// Benchmark "./test_runs/structural2_key-2-3-4-5--s-120240927_164306/ITC99/b15_encrypted" written by ABC on Fri Sep 27 18:32:53 2024

module b15_encrypted  ( clock, 
    DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
    DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
    DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
    DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
    DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
    DATAI_0_, NA_N, BS16_N, READY_N, HOLD, keyinput0, keyinput1, keyinput2,
    BE_N_REG_3_, BE_N_REG_2_, BE_N_REG_1_, BE_N_REG_0_, ADDRESS_REG_29_,
    ADDRESS_REG_28_, ADDRESS_REG_27_, ADDRESS_REG_26_, ADDRESS_REG_25_,
    ADDRESS_REG_24_, ADDRESS_REG_23_, ADDRESS_REG_22_, ADDRESS_REG_21_,
    ADDRESS_REG_20_, ADDRESS_REG_19_, ADDRESS_REG_18_, ADDRESS_REG_17_,
    ADDRESS_REG_16_, ADDRESS_REG_15_, ADDRESS_REG_14_, ADDRESS_REG_13_,
    ADDRESS_REG_12_, ADDRESS_REG_11_, ADDRESS_REG_10_, ADDRESS_REG_9_,
    ADDRESS_REG_8_, ADDRESS_REG_7_, ADDRESS_REG_6_, ADDRESS_REG_5_,
    ADDRESS_REG_4_, ADDRESS_REG_3_, ADDRESS_REG_2_, ADDRESS_REG_1_,
    ADDRESS_REG_0_, W_R_N_REG, D_C_N_REG, M_IO_N_REG, ADS_N_REG,
    DATAO_REG_31_, DATAO_REG_30_, DATAO_REG_29_, DATAO_REG_28_,
    DATAO_REG_27_, DATAO_REG_26_, DATAO_REG_25_, DATAO_REG_24_,
    DATAO_REG_23_, DATAO_REG_22_, DATAO_REG_21_, DATAO_REG_20_,
    DATAO_REG_19_, DATAO_REG_18_, DATAO_REG_17_, DATAO_REG_16_,
    DATAO_REG_15_, DATAO_REG_14_, DATAO_REG_13_, DATAO_REG_12_,
    DATAO_REG_11_, DATAO_REG_10_, DATAO_REG_9_, DATAO_REG_8_, DATAO_REG_7_,
    DATAO_REG_6_, DATAO_REG_5_, DATAO_REG_4_, DATAO_REG_3_, DATAO_REG_2_,
    DATAO_REG_1_, DATAO_REG_0_  );
  input  clock;
  input  DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_,
    DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_,
    DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_,
    DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_,
    DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_,
    DATAI_1_, DATAI_0_, NA_N, BS16_N, READY_N, HOLD, keyinput0, keyinput1,
    keyinput2;
  output BE_N_REG_3_, BE_N_REG_2_, BE_N_REG_1_, BE_N_REG_0_, ADDRESS_REG_29_,
    ADDRESS_REG_28_, ADDRESS_REG_27_, ADDRESS_REG_26_, ADDRESS_REG_25_,
    ADDRESS_REG_24_, ADDRESS_REG_23_, ADDRESS_REG_22_, ADDRESS_REG_21_,
    ADDRESS_REG_20_, ADDRESS_REG_19_, ADDRESS_REG_18_, ADDRESS_REG_17_,
    ADDRESS_REG_16_, ADDRESS_REG_15_, ADDRESS_REG_14_, ADDRESS_REG_13_,
    ADDRESS_REG_12_, ADDRESS_REG_11_, ADDRESS_REG_10_, ADDRESS_REG_9_,
    ADDRESS_REG_8_, ADDRESS_REG_7_, ADDRESS_REG_6_, ADDRESS_REG_5_,
    ADDRESS_REG_4_, ADDRESS_REG_3_, ADDRESS_REG_2_, ADDRESS_REG_1_,
    ADDRESS_REG_0_, W_R_N_REG, D_C_N_REG, M_IO_N_REG, ADS_N_REG,
    DATAO_REG_31_, DATAO_REG_30_, DATAO_REG_29_, DATAO_REG_28_,
    DATAO_REG_27_, DATAO_REG_26_, DATAO_REG_25_, DATAO_REG_24_,
    DATAO_REG_23_, DATAO_REG_22_, DATAO_REG_21_, DATAO_REG_20_,
    DATAO_REG_19_, DATAO_REG_18_, DATAO_REG_17_, DATAO_REG_16_,
    DATAO_REG_15_, DATAO_REG_14_, DATAO_REG_13_, DATAO_REG_12_,
    DATAO_REG_11_, DATAO_REG_10_, DATAO_REG_9_, DATAO_REG_8_, DATAO_REG_7_,
    DATAO_REG_6_, DATAO_REG_5_, DATAO_REG_4_, DATAO_REG_3_, DATAO_REG_2_,
    DATAO_REG_1_, DATAO_REG_0_;
  reg BE_N_REG_3_, BE_N_REG_2_, BE_N_REG_1_, BE_N_REG_0_, ADDRESS_REG_29_,
    ADDRESS_REG_28_, ADDRESS_REG_27_, ADDRESS_REG_26_, ADDRESS_REG_25_,
    ADDRESS_REG_24_, ADDRESS_REG_23_, ADDRESS_REG_22_, ADDRESS_REG_21_,
    ADDRESS_REG_20_, ADDRESS_REG_19_, ADDRESS_REG_18_, ADDRESS_REG_17_,
    ADDRESS_REG_16_, ADDRESS_REG_15_, ADDRESS_REG_14_, ADDRESS_REG_13_,
    ADDRESS_REG_12_, ADDRESS_REG_11_, ADDRESS_REG_10_, ADDRESS_REG_9_,
    ADDRESS_REG_8_, ADDRESS_REG_7_, ADDRESS_REG_6_, ADDRESS_REG_5_,
    ADDRESS_REG_4_, ADDRESS_REG_3_, ADDRESS_REG_2_, ADDRESS_REG_1_,
    ADDRESS_REG_0_, STATE_REG_2_, STATE_REG_1_, STATE_REG_0_,
    DATAWIDTH_REG_0_, DATAWIDTH_REG_1_, DATAWIDTH_REG_2_, DATAWIDTH_REG_3_,
    DATAWIDTH_REG_4_, DATAWIDTH_REG_5_, DATAWIDTH_REG_6_, DATAWIDTH_REG_7_,
    DATAWIDTH_REG_8_, DATAWIDTH_REG_9_, DATAWIDTH_REG_10_,
    DATAWIDTH_REG_11_, DATAWIDTH_REG_12_, DATAWIDTH_REG_13_,
    DATAWIDTH_REG_14_, DATAWIDTH_REG_15_, DATAWIDTH_REG_16_,
    DATAWIDTH_REG_17_, DATAWIDTH_REG_18_, DATAWIDTH_REG_19_,
    DATAWIDTH_REG_20_, DATAWIDTH_REG_21_, DATAWIDTH_REG_22_,
    DATAWIDTH_REG_23_, DATAWIDTH_REG_24_, DATAWIDTH_REG_25_,
    DATAWIDTH_REG_26_, DATAWIDTH_REG_27_, DATAWIDTH_REG_28_,
    DATAWIDTH_REG_29_, DATAWIDTH_REG_30_, DATAWIDTH_REG_31_, STATE2_REG_3_,
    STATE2_REG_2_, STATE2_REG_1_, STATE2_REG_0_, INSTQUEUE_REG_15__7_,
    INSTQUEUE_REG_15__6_, INSTQUEUE_REG_15__5_, INSTQUEUE_REG_15__4_,
    INSTQUEUE_REG_15__3_, INSTQUEUE_REG_15__2_, INSTQUEUE_REG_15__1_,
    INSTQUEUE_REG_15__0_, INSTQUEUE_REG_14__7_, INSTQUEUE_REG_14__6_,
    INSTQUEUE_REG_14__5_, INSTQUEUE_REG_14__4_, INSTQUEUE_REG_14__3_,
    INSTQUEUE_REG_14__2_, INSTQUEUE_REG_14__1_, INSTQUEUE_REG_14__0_,
    INSTQUEUE_REG_13__7_, INSTQUEUE_REG_13__6_, INSTQUEUE_REG_13__5_,
    INSTQUEUE_REG_13__4_, INSTQUEUE_REG_13__3_, INSTQUEUE_REG_13__2_,
    INSTQUEUE_REG_13__1_, INSTQUEUE_REG_13__0_, INSTQUEUE_REG_12__7_,
    INSTQUEUE_REG_12__6_, INSTQUEUE_REG_12__5_, INSTQUEUE_REG_12__4_,
    INSTQUEUE_REG_12__3_, INSTQUEUE_REG_12__2_, INSTQUEUE_REG_12__1_,
    INSTQUEUE_REG_12__0_, INSTQUEUE_REG_11__7_, INSTQUEUE_REG_11__6_,
    INSTQUEUE_REG_11__5_, INSTQUEUE_REG_11__4_, INSTQUEUE_REG_11__3_,
    INSTQUEUE_REG_11__2_, INSTQUEUE_REG_11__1_, INSTQUEUE_REG_11__0_,
    INSTQUEUE_REG_10__7_, INSTQUEUE_REG_10__6_, INSTQUEUE_REG_10__5_,
    INSTQUEUE_REG_10__4_, INSTQUEUE_REG_10__3_, INSTQUEUE_REG_10__2_,
    INSTQUEUE_REG_10__1_, INSTQUEUE_REG_10__0_, INSTQUEUE_REG_9__7_,
    INSTQUEUE_REG_9__6_, INSTQUEUE_REG_9__5_, INSTQUEUE_REG_9__4_,
    INSTQUEUE_REG_9__3_, INSTQUEUE_REG_9__2_, INSTQUEUE_REG_9__1_,
    INSTQUEUE_REG_9__0_, INSTQUEUE_REG_8__7_, INSTQUEUE_REG_8__6_,
    INSTQUEUE_REG_8__5_, INSTQUEUE_REG_8__4_, INSTQUEUE_REG_8__3_,
    INSTQUEUE_REG_8__2_, INSTQUEUE_REG_8__1_, INSTQUEUE_REG_8__0_,
    INSTQUEUE_REG_7__7_, INSTQUEUE_REG_7__6_, INSTQUEUE_REG_7__5_,
    INSTQUEUE_REG_7__4_, INSTQUEUE_REG_7__3_, INSTQUEUE_REG_7__2_,
    INSTQUEUE_REG_7__1_, INSTQUEUE_REG_7__0_, INSTQUEUE_REG_6__7_,
    INSTQUEUE_REG_6__6_, INSTQUEUE_REG_6__5_, INSTQUEUE_REG_6__4_,
    INSTQUEUE_REG_6__3_, INSTQUEUE_REG_6__2_, INSTQUEUE_REG_6__1_,
    INSTQUEUE_REG_6__0_, INSTQUEUE_REG_5__7_, INSTQUEUE_REG_5__6_,
    INSTQUEUE_REG_5__5_, INSTQUEUE_REG_5__4_, INSTQUEUE_REG_5__3_,
    INSTQUEUE_REG_5__2_, INSTQUEUE_REG_5__1_, INSTQUEUE_REG_5__0_,
    INSTQUEUE_REG_4__7_, INSTQUEUE_REG_4__6_, INSTQUEUE_REG_4__5_,
    INSTQUEUE_REG_4__4_, INSTQUEUE_REG_4__3_, INSTQUEUE_REG_4__2_,
    INSTQUEUE_REG_4__1_, INSTQUEUE_REG_4__0_, INSTQUEUE_REG_3__7_,
    INSTQUEUE_REG_3__6_, INSTQUEUE_REG_3__5_, INSTQUEUE_REG_3__4_,
    INSTQUEUE_REG_3__3_, INSTQUEUE_REG_3__2_, INSTQUEUE_REG_3__1_,
    INSTQUEUE_REG_3__0_, INSTQUEUE_REG_2__7_, INSTQUEUE_REG_2__6_,
    INSTQUEUE_REG_2__5_, INSTQUEUE_REG_2__4_, INSTQUEUE_REG_2__3_,
    INSTQUEUE_REG_2__2_, INSTQUEUE_REG_2__1_, INSTQUEUE_REG_2__0_,
    INSTQUEUE_REG_1__7_, INSTQUEUE_REG_1__6_, INSTQUEUE_REG_1__5_,
    INSTQUEUE_REG_1__4_, INSTQUEUE_REG_1__3_, INSTQUEUE_REG_1__2_,
    INSTQUEUE_REG_1__1_, INSTQUEUE_REG_1__0_, INSTQUEUE_REG_0__7_,
    INSTQUEUE_REG_0__6_, INSTQUEUE_REG_0__5_, INSTQUEUE_REG_0__4_,
    INSTQUEUE_REG_0__3_, INSTQUEUE_REG_0__2_, INSTQUEUE_REG_0__1_,
    INSTQUEUE_REG_0__0_, INSTQUEUERD_ADDR_REG_4_, INSTQUEUERD_ADDR_REG_3_,
    INSTQUEUERD_ADDR_REG_2_, INSTQUEUERD_ADDR_REG_1_,
    INSTQUEUERD_ADDR_REG_0_, INSTQUEUEWR_ADDR_REG_4_,
    INSTQUEUEWR_ADDR_REG_3_, INSTQUEUEWR_ADDR_REG_2_,
    INSTQUEUEWR_ADDR_REG_1_, INSTQUEUEWR_ADDR_REG_0_,
    INSTADDRPOINTER_REG_0_, INSTADDRPOINTER_REG_1_, INSTADDRPOINTER_REG_2_,
    INSTADDRPOINTER_REG_3_, INSTADDRPOINTER_REG_4_, INSTADDRPOINTER_REG_5_,
    INSTADDRPOINTER_REG_6_, INSTADDRPOINTER_REG_7_, INSTADDRPOINTER_REG_8_,
    INSTADDRPOINTER_REG_9_, INSTADDRPOINTER_REG_10_,
    INSTADDRPOINTER_REG_11_, INSTADDRPOINTER_REG_12_,
    INSTADDRPOINTER_REG_13_, INSTADDRPOINTER_REG_14_,
    INSTADDRPOINTER_REG_15_, INSTADDRPOINTER_REG_16_,
    INSTADDRPOINTER_REG_17_, INSTADDRPOINTER_REG_18_,
    INSTADDRPOINTER_REG_19_, INSTADDRPOINTER_REG_20_,
    INSTADDRPOINTER_REG_21_, INSTADDRPOINTER_REG_22_,
    INSTADDRPOINTER_REG_23_, INSTADDRPOINTER_REG_24_,
    INSTADDRPOINTER_REG_25_, INSTADDRPOINTER_REG_26_,
    INSTADDRPOINTER_REG_27_, INSTADDRPOINTER_REG_28_,
    INSTADDRPOINTER_REG_29_, INSTADDRPOINTER_REG_30_,
    INSTADDRPOINTER_REG_31_, PHYADDRPOINTER_REG_0_, PHYADDRPOINTER_REG_1_,
    PHYADDRPOINTER_REG_2_, PHYADDRPOINTER_REG_3_, PHYADDRPOINTER_REG_4_,
    PHYADDRPOINTER_REG_5_, PHYADDRPOINTER_REG_6_, PHYADDRPOINTER_REG_7_,
    PHYADDRPOINTER_REG_8_, PHYADDRPOINTER_REG_9_, PHYADDRPOINTER_REG_10_,
    PHYADDRPOINTER_REG_11_, PHYADDRPOINTER_REG_12_, PHYADDRPOINTER_REG_13_,
    PHYADDRPOINTER_REG_14_, PHYADDRPOINTER_REG_15_, PHYADDRPOINTER_REG_16_,
    PHYADDRPOINTER_REG_17_, PHYADDRPOINTER_REG_18_, PHYADDRPOINTER_REG_19_,
    PHYADDRPOINTER_REG_20_, PHYADDRPOINTER_REG_21_, PHYADDRPOINTER_REG_22_,
    PHYADDRPOINTER_REG_23_, PHYADDRPOINTER_REG_24_, PHYADDRPOINTER_REG_25_,
    PHYADDRPOINTER_REG_26_, PHYADDRPOINTER_REG_27_, PHYADDRPOINTER_REG_28_,
    PHYADDRPOINTER_REG_29_, PHYADDRPOINTER_REG_30_, PHYADDRPOINTER_REG_31_,
    LWORD_REG_15_, LWORD_REG_14_, LWORD_REG_13_, LWORD_REG_12_,
    LWORD_REG_11_, LWORD_REG_10_, LWORD_REG_9_, LWORD_REG_8_, LWORD_REG_7_,
    LWORD_REG_6_, LWORD_REG_5_, LWORD_REG_4_, LWORD_REG_3_, LWORD_REG_2_,
    LWORD_REG_1_, LWORD_REG_0_, UWORD_REG_14_, UWORD_REG_13_,
    UWORD_REG_12_, UWORD_REG_11_, UWORD_REG_10_, UWORD_REG_9_,
    UWORD_REG_8_, UWORD_REG_7_, UWORD_REG_6_, UWORD_REG_5_, UWORD_REG_4_,
    UWORD_REG_3_, UWORD_REG_2_, UWORD_REG_1_, UWORD_REG_0_, DATAO_REG_0_,
    DATAO_REG_1_, DATAO_REG_2_, DATAO_REG_3_, DATAO_REG_4_, DATAO_REG_5_,
    DATAO_REG_6_, DATAO_REG_7_, DATAO_REG_8_, DATAO_REG_9_, DATAO_REG_10_,
    DATAO_REG_11_, DATAO_REG_12_, DATAO_REG_13_, DATAO_REG_14_,
    DATAO_REG_15_, DATAO_REG_16_, DATAO_REG_17_, DATAO_REG_18_,
    DATAO_REG_19_, DATAO_REG_20_, DATAO_REG_21_, DATAO_REG_22_,
    DATAO_REG_23_, DATAO_REG_24_, DATAO_REG_25_, DATAO_REG_26_,
    DATAO_REG_27_, DATAO_REG_28_, DATAO_REG_29_, DATAO_REG_30_,
    DATAO_REG_31_, EAX_REG_0_, EAX_REG_1_, EAX_REG_2_, EAX_REG_3_,
    EAX_REG_4_, EAX_REG_5_, EAX_REG_6_, EAX_REG_7_, EAX_REG_8_, EAX_REG_9_,
    EAX_REG_10_, EAX_REG_11_, EAX_REG_12_, EAX_REG_13_, EAX_REG_14_,
    EAX_REG_15_, EAX_REG_16_, EAX_REG_17_, EAX_REG_18_, EAX_REG_19_,
    EAX_REG_20_, EAX_REG_21_, EAX_REG_22_, EAX_REG_23_, EAX_REG_24_,
    EAX_REG_25_, EAX_REG_26_, EAX_REG_27_, EAX_REG_28_, EAX_REG_29_,
    EAX_REG_30_, EAX_REG_31_, EBX_REG_0_, EBX_REG_1_, EBX_REG_2_,
    EBX_REG_3_, EBX_REG_4_, EBX_REG_5_, EBX_REG_6_, EBX_REG_7_, EBX_REG_8_,
    EBX_REG_9_, EBX_REG_10_, EBX_REG_11_, EBX_REG_12_, EBX_REG_13_,
    EBX_REG_14_, EBX_REG_15_, EBX_REG_16_, EBX_REG_17_, EBX_REG_18_,
    EBX_REG_19_, EBX_REG_20_, EBX_REG_21_, EBX_REG_22_, EBX_REG_23_,
    EBX_REG_24_, EBX_REG_25_, EBX_REG_26_, EBX_REG_27_, EBX_REG_28_,
    EBX_REG_29_, EBX_REG_30_, EBX_REG_31_, REIP_REG_0_, REIP_REG_1_,
    REIP_REG_2_, REIP_REG_3_, REIP_REG_4_, REIP_REG_5_, REIP_REG_6_,
    REIP_REG_7_, REIP_REG_8_, REIP_REG_9_, REIP_REG_10_, REIP_REG_11_,
    REIP_REG_12_, REIP_REG_13_, REIP_REG_14_, REIP_REG_15_, REIP_REG_16_,
    REIP_REG_17_, REIP_REG_18_, REIP_REG_19_, REIP_REG_20_, REIP_REG_21_,
    REIP_REG_22_, REIP_REG_23_, REIP_REG_24_, REIP_REG_25_, REIP_REG_26_,
    REIP_REG_27_, REIP_REG_28_, REIP_REG_29_, REIP_REG_30_, REIP_REG_31_,
    BYTEENABLE_REG_3_, BYTEENABLE_REG_2_, BYTEENABLE_REG_1_,
    BYTEENABLE_REG_0_, W_R_N_REG, FLUSH_REG, MORE_REG, STATEBS16_REG,
    REQUESTPENDING_REG, D_C_N_REG, M_IO_N_REG, CODEFETCH_REG, ADS_N_REG,
    READREQUEST_REG, MEMORYFETCH_REG, Q_0, Q_1;
  wire new_ADD_515_U182, new_ADD_515_U181, new_ADD_515_U180, new_U2352,
    new_U2353, new_U2354, new_U2355, new_U2356, new_U2357, new_U2358,
    new_U2359, new_U2360, new_U2361, new_U2362, new_U2363, new_U2364,
    new_U2365, new_U2366, new_U2367, new_U2368, new_U2369, new_U2370,
    new_U2371, new_U2372, new_U2373, new_U2374, new_U2375, new_U2376,
    new_U2377, new_U2378, new_U2379, new_U2380, new_U2381, new_U2382,
    new_U2383, new_U2384, new_U2385, new_U2386, new_U2387, new_U2388,
    new_U2389, new_U2390, new_U2391, new_U2392, new_U2393, new_U2394,
    new_U2395, new_U2396, new_U2397, new_U2398, new_U2399, new_U2400,
    new_U2401, new_U2402, new_U2403, new_U2404, new_U2405, new_U2406,
    new_U2407, new_U2408, new_U2409, new_U2410, new_U2411, new_U2412,
    new_U2413, new_U2414, new_U2415, new_U2416, new_U2417, new_U2418,
    new_U2419, new_U2420, new_U2421, new_U2422, new_U2423, new_U2424,
    new_U2425, new_U2426, new_U2427, new_U2428, new_U2429, new_U2430,
    new_U2431, new_U2432, new_U2433, new_U2434, new_U2435, new_U2436,
    new_U2437, new_U2438, new_U2439, new_U2440, new_U2441, new_U2442,
    new_U2443, new_U2444, new_U2445, new_U2446, new_U2447, new_U2448,
    new_U2449, new_U2450, new_U2451, new_U2452, new_U2453, new_U2454,
    new_U2455, new_U2456, new_U2457, new_U2458, new_U2459, new_U2460,
    new_U2461, new_U2462, new_U2463, new_U2464, new_U2465, new_U2466,
    new_U2467, new_U2468, new_U2469, new_U2470, new_U2471, new_U2472,
    new_U2473, new_U2474, new_U2475, new_U2476, new_U2477, new_U2478,
    new_U2479, new_U2480, new_U2481, new_U2482, new_U2483, new_U2484,
    new_U2485, new_U2486, new_U2487, new_U2488, new_U2489, new_U2490,
    new_U2491, new_U2492, new_U2493, new_U2494, new_U2495, new_U2496,
    new_U2497, new_U2498, new_U2499, new_U2500, new_U2501, new_U2502,
    new_U2503, new_U2504, new_U2505, new_U2506, new_U2507, new_U2508,
    new_U2509, new_U2510, new_U2511, new_U2512, new_U2513, new_U2514,
    new_U2515, new_U2516, new_U2517, new_U2518, new_U2519, new_U2520,
    new_U2521, new_U2522, new_U2523, new_U2524, new_U2525, new_U2526,
    new_U2527, new_U2528, new_U2529, new_U2530, new_U2531, new_U2532,
    new_U2533, new_U2534, new_U2535, new_U2536, new_U2537, new_U2538,
    new_U2539, new_U2540, new_U2541, new_U2542, new_U2543, new_U2544,
    new_U2545, new_U2546, new_U2547, new_U2548, new_U2549, new_U2550,
    new_U2551, new_U2552, new_U2553, new_U2554, new_U2555, new_U2556,
    new_U2557, new_U2558, new_U2559, new_U2560, new_U2561, new_U2562,
    new_U2563, new_U2564, new_U2565, new_U2566, new_U2567, new_U2568,
    new_U2569, new_U2570, new_U2571, new_U2572, new_U2573, new_U2574,
    new_U2575, new_U2576, new_U2577, new_U2578, new_U2579, new_U2580,
    new_U2581, new_U2582, new_U2583, new_U2584, new_U2585, new_U2586,
    new_U2587, new_U2588, new_U2589, new_U2590, new_U2591, new_U2592,
    new_U2593, new_U2594, new_U2595, new_U2596, new_U2597, new_U2598,
    new_U2599, new_U2600, new_U2601, new_U2602, new_U2603, new_U2604,
    new_U2605, new_U2606, new_U2607, new_U2608, new_U2609, new_U2610,
    new_U2611, new_U2612, new_U2613, new_U2614, new_U2615, new_U2616,
    new_U2617, new_U2618, new_ADD_515_U179, new_U2620, new_U2621,
    new_U2622, new_U2623, new_U2624, new_U2625, new_U2626, new_U2627,
    new_U2628, new_U2629, new_U2630, new_U2631, new_U2632, new_U2633,
    new_U2634, new_U2635, new_U2636, new_U2637, new_U2638, new_U2639,
    new_U2640, new_U2641, new_U2642, new_U2643, new_U2644, new_U2645,
    new_U2646, new_U2647, new_U2648, new_U2649, new_U2650, new_U2651,
    new_U2652, new_U2653, new_U2654, new_U2655, new_U2656, new_U2657,
    new_U2658, new_U2659, new_U2660, new_U2661, new_U2662, new_U2663,
    new_U2664, new_U2665, new_U2666, new_U2667, new_U2668, new_U2669,
    new_U2670, new_U2671, new_U2672, new_U2673, new_U2674, new_U2675,
    new_U2676, new_U2677, new_U2678, new_U2679, new_U2680, new_U2681,
    new_U2682, new_U2683, new_U2684, new_U2685, new_U2686, new_U2687,
    new_U2688, new_U2689, new_U2690, new_U2691, new_U2692, new_U2693,
    new_U2694, new_U2695, new_U2696, new_U2697, new_U2698, new_U2699,
    new_U2700, new_U2701, new_U2702, new_U2703, new_U2704, new_U2705,
    new_U2706, new_U2707, new_U2708, new_U2709, new_U2710, new_U2711,
    new_U2712, new_U2713, new_U2714, new_U2715, new_U2716, new_U2717,
    new_U2718, new_U2719, new_U2720, new_U2721, new_U2722, new_U2723,
    new_U2724, new_U2725, new_U2726, new_U2727, new_U2728, new_U2729,
    new_U2730, new_U2731, new_U2732, new_U2733, new_U2734, new_U2735,
    new_U2736, new_U2737, new_U2738, new_U2739, new_U2740, new_U2741,
    new_U2742, new_U2743, new_U2744, new_U2745, new_U2746, new_U2747,
    new_U2748, new_U2749, new_U2750, new_U2751, new_U2752, new_U2753,
    new_U2754, new_U2755, new_U2756, new_U2757, new_U2758, new_U2759,
    new_U2760, new_U2761, new_U2762, new_U2763, new_U2764, new_U2765,
    new_U2766, new_U2767, new_U2768, new_U2769, new_U2770, new_U2771,
    new_U2772, new_U2773, new_U2774, new_U2775, new_U2776, new_U2777,
    new_U2778, new_U2779, new_U2780, new_U2781, new_U2782, new_U2783,
    new_U2784, new_U2785, new_U2786, new_U2787, new_U3214, new_U3215,
    new_U3216, new_U3217, new_U3218, new_U3219, new_U3220, new_U3221,
    new_U3222, new_U3223, new_U3224, new_U3225, new_U3226, new_U3227,
    new_U3228, new_U3229, new_U3230, new_U3231, new_U3232, new_U3233,
    new_U3234, new_U3235, new_U3236, new_U3237, new_U3238, new_U3239,
    new_U3240, new_U3241, new_U3242, new_U3243, new_U3244, new_U3245,
    new_U3246, new_U3247, new_U3248, new_U3249, new_U3250, new_U3251,
    new_U3252, new_U3253, new_U3254, new_U3255, new_U3256, new_U3257,
    new_U3258, new_U3259, new_U3260, new_U3261, new_U3262, new_U3263,
    new_U3264, new_U3265, new_U3266, new_U3267, new_U3268, new_U3269,
    new_U3270, new_U3271, new_U3272, new_U3273, new_U3274, new_U3275,
    new_U3276, new_U3277, new_U3278, new_U3279, new_U3280, new_U3281,
    new_U3282, new_U3283, new_U3284, new_U3285, new_U3286, new_U3287,
    new_U3288, new_U3289, new_U3290, new_U3291, new_U3292, new_U3293,
    new_U3294, new_U3295, new_U3296, new_U3297, new_U3298, new_U3299,
    new_U3300, new_U3301, new_U3302, new_U3303, new_U3304, new_U3305,
    new_U3306, new_U3307, new_U3308, new_U3309, new_U3310, new_U3311,
    new_U3312, new_U3313, new_U3314, new_U3315, new_U3316, new_U3317,
    new_U3318, new_U3319, new_U3320, new_U3321, new_U3322, new_U3323,
    new_U3324, new_U3325, new_U3326, new_U3327, new_U3328, new_U3329,
    new_U3330, new_U3331, new_U3332, new_U3333, new_U3334, new_U3335,
    new_U3336, new_U3337, new_U3338, new_U3339, new_U3340, new_U3341,
    new_U3342, new_U3343, new_U3344, new_U3345, new_U3346, new_U3347,
    new_U3348, new_U3349, new_U3350, new_U3351, new_U3352, new_U3353,
    new_U3354, new_U3355, new_U3356, new_U3357, new_U3358, new_U3359,
    new_U3360, new_U3361, new_U3362, new_U3363, new_U3364, new_U3365,
    new_U3366, new_U3367, new_U3368, new_U3369, new_U3370, new_U3371,
    new_U3372, new_U3373, new_U3374, new_U3375, new_U3376, new_U3377,
    new_U3378, new_U3379, new_U3380, new_U3381, new_U3382, new_U3383,
    new_U3384, new_U3385, new_U3386, new_U3387, new_U3388, new_U3389,
    new_U3390, new_U3391, new_U3392, new_U3393, new_U3394, new_U3395,
    new_U3396, new_U3397, new_U3398, new_U3399, new_U3400, new_U3401,
    new_U3402, new_U3403, new_U3404, new_U3405, new_U3406, new_U3407,
    new_U3408, new_U3409, new_U3410, new_U3411, new_U3412, new_U3413,
    new_U3414, new_U3415, new_U3416, new_U3417, new_U3418, new_U3419,
    new_U3420, new_U3421, new_U3422, new_U3423, new_U3424, new_U3425,
    new_U3426, new_U3427, new_U3428, new_U3429, new_U3430, new_U3431,
    new_U3432, new_U3433, new_U3434, new_U3435, new_U3436, new_U3437,
    new_U3438, new_U3439, new_U3440, new_U3441, new_U3442, new_U3443,
    new_U3444, new_U3445, new_U3449, new_U3450, new_U3454, new_U3457,
    new_U3458, new_U3466, new_U3467, new_U3475, new_U3476, new_U3477,
    new_U3478, new_U3479, new_U3480, new_U3481, new_U3482, new_U3483,
    new_U3484, new_U3485, new_U3486, new_U3487, new_U3488, new_U3489,
    new_U3490, new_U3491, new_U3492, new_U3493, new_U3494, new_U3495,
    new_U3496, new_U3497, new_U3498, new_U3499, new_U3500, new_U3501,
    new_U3502, new_U3503, new_U3504, new_U3505, new_U3506, new_U3507,
    new_U3508, new_U3509, new_U3510, new_U3511, new_U3512, new_U3513,
    new_U3514, new_U3515, new_U3516, new_U3517, new_U3518, new_U3519,
    new_U3520, new_U3521, new_U3522, new_U3523, new_U3524, new_U3525,
    new_U3526, new_U3527, new_U3528, new_U3529, new_U3530, new_U3531,
    new_U3532, new_U3533, new_U3534, new_U3535, new_U3536, new_U3537,
    new_U3538, new_U3539, new_U3540, new_U3541, new_U3542, new_U3543,
    new_U3544, new_U3545, new_U3546, new_U3547, new_U3548, new_U3549,
    new_U3550, new_U3551, new_U3552, new_U3553, new_U3554, new_U3555,
    new_U3556, new_U3557, new_U3558, new_U3559, new_U3560, new_U3561,
    new_U3562, new_U3563, new_U3564, new_U3565, new_U3566, new_U3567,
    new_U3568, new_U3569, new_U3570, new_U3571, new_U3572, new_U3573,
    new_U3574, new_U3575, new_U3576, new_U3577, new_U3578, new_U3579,
    new_U3580, new_U3581, new_U3582, new_U3583, new_U3584, new_U3585,
    new_U3586, new_U3587, new_U3588, new_U3589, new_U3590, new_U3591,
    new_U3592, new_U3593, new_U3594, new_U3595, new_U3596, new_U3597,
    new_U3598, new_U3599, new_U3600, new_U3601, new_U3602, new_U3603,
    new_U3604, new_U3605, new_U3606, new_U3607, new_U3608, new_U3609,
    new_U3610, new_U3611, new_U3612, new_U3613, new_U3614, new_U3615,
    new_U3616, new_U3617, new_U3618, new_U3619, new_U3620, new_U3621,
    new_U3622, new_U3623, new_U3624, new_U3625, new_U3626, new_U3627,
    new_U3628, new_U3629, new_U3630, new_U3631, new_U3632, new_U3633,
    new_U3634, new_U3635, new_U3636, new_U3637, new_U3638, new_U3639,
    new_U3640, new_U3641, new_U3642, new_U3643, new_U3644, new_U3645,
    new_U3646, new_U3647, new_U3648, new_U3649, new_U3650, new_U3651,
    new_U3652, new_U3653, new_U3654, new_U3655, new_U3656, new_U3657,
    new_U3658, new_U3659, new_U3660, new_U3661, new_U3662, new_U3663,
    new_U3664, new_U3665, new_U3666, new_U3667, new_U3668, new_U3669,
    new_U3670, new_U3671, new_U3672, new_U3673, new_U3674, new_U3675,
    new_U3676, new_U3677, new_U3678, new_U3679, new_U3680, new_U3681,
    new_U3682, new_U3683, new_U3684, new_U3685, new_U3686, new_U3687,
    new_U3688, new_U3689, new_U3690, new_U3691, new_U3692, new_U3693,
    new_U3694, new_U3695, new_U3696, new_U3697, new_U3698, new_U3699,
    new_U3700, new_U3701, new_U3702, new_U3703, new_U3704, new_U3705,
    new_U3706, new_U3707, new_U3708, new_U3709, new_U3710, new_U3711,
    new_U3712, new_U3713, new_U3714, new_U3715, new_U3716, new_U3717,
    new_U3718, new_U3719, new_U3720, new_U3721, new_U3722, new_U3723,
    new_U3724, new_U3725, new_U3726, new_U3727, new_U3728, new_U3729,
    new_U3730, new_U3731, new_U3732, new_U3733, new_U3734, new_U3735,
    new_U3736, new_U3737, new_U3738, new_U3739, new_U3740, new_U3741,
    new_U3742, new_U3743, new_U3744, new_U3745, new_U3746, new_U3747,
    new_U3748, new_U3749, new_U3750, new_U3751, new_U3752, new_U3753,
    new_U3754, new_U3755, new_U3756, new_U3757, new_U3758, new_U3759,
    new_U3760, new_U3761, new_U3762, new_U3763, new_U3764, new_U3765,
    new_U3766, new_U3767, new_U3768, new_U3769, new_U3770, new_U3771,
    new_U3772, new_U3773, new_U3774, new_U3775, new_U3776, new_U3777,
    new_U3778, new_U3779, new_U3780, new_U3781, new_U3782, new_U3783,
    new_U3784, new_U3785, new_U3786, new_U3787, new_U3788, new_U3789,
    new_U3790, new_U3791, new_U3792, new_U3793, new_U3794, new_U3795,
    new_U3796, new_U3797, new_U3798, new_U3799, new_U3800, new_U3801,
    new_U3802, new_U3803, new_U3804, new_U3805, new_U3806, new_U3807,
    new_U3808, new_U3809, new_U3810, new_U3811, new_U3812, new_U3813,
    new_U3814, new_U3815, new_U3816, new_U3817, new_U3818, new_U3819,
    new_U3820, new_U3821, new_U3822, new_U3823, new_U3824, new_U3825,
    new_U3826, new_U3827, new_U3828, new_U3829, new_U3830, new_U3831,
    new_U3832, new_U3833, new_U3834, new_U3835, new_U3836, new_U3837,
    new_U3838, new_U3839, new_U3840, new_U3841, new_U3842, new_U3843,
    new_U3844, new_U3845, new_U3846, new_U3847, new_U3848, new_U3849,
    new_U3850, new_U3851, new_U3852, new_U3853, new_U3854, new_U3855,
    new_U3856, new_U3857, new_U3858, new_U3859, new_U3860, new_U3861,
    new_U3862, new_U3863, new_U3864, new_U3865, new_U3866, new_U3867,
    new_U3868, new_U3869, new_U3870, new_U3871, new_U3872, new_U3873,
    new_U3874, new_U3875, new_U3876, new_U3877, new_U3878, new_U3879,
    new_U3880, new_U3881, new_U3882, new_U3883, new_U3884, new_U3885,
    new_U3886, new_U3887, new_U3888, new_U3889, new_U3890, new_U3891,
    new_U3892, new_U3893, new_U3894, new_U3895, new_U3896, new_U3897,
    new_U3898, new_U3899, new_U3900, new_U3901, new_U3902, new_U3903,
    new_U3904, new_U3905, new_U3906, new_U3907, new_U3908, new_U3909,
    new_U3910, new_U3911, new_U3912, new_U3913, new_U3914, new_U3915,
    new_U3916, new_U3917, new_U3918, new_U3919, new_U3920, new_U3921,
    new_U3922, new_U3923, new_U3924, new_U3925, new_U3926, new_U3927,
    new_U3928, new_U3929, new_U3930, new_U3931, new_U3932, new_U3933,
    new_U3934, new_U3935, new_U3936, new_U3937, new_U3938, new_U3939,
    new_U3940, new_U3941, new_U3942, new_U3943, new_U3944, new_U3945,
    new_U3946, new_U3947, new_U3948, new_U3949, new_U3950, new_U3951,
    new_U3952, new_U3953, new_U3954, new_U3955, new_U3956, new_U3957,
    new_U3958, new_U3959, new_U3960, new_U3961, new_U3962, new_U3963,
    new_U3964, new_U3965, new_U3966, new_U3967, new_U3968, new_U3969,
    new_U3970, new_U3971, new_U3972, new_U3973, new_U3974, new_U3975,
    new_U3976, new_U3977, new_U3978, new_U3979, new_U3980, new_U3981,
    new_U3982, new_U3983, new_U3984, new_U3985, new_U3986, new_U3987,
    new_U3988, new_U3989, new_U3990, new_U3991, new_U3992, new_U3993,
    new_U3994, new_U3995, new_U3996, new_U3997, new_U3998, new_U3999,
    new_U4000, new_U4001, new_U4002, new_U4003, new_U4004, new_U4005,
    new_U4006, new_U4007, new_U4008, new_U4009, new_U4010, new_U4011,
    new_U4012, new_U4013, new_U4014, new_U4015, new_U4016, new_U4017,
    new_U4018, new_U4019, new_U4020, new_U4021, new_U4022, new_U4023,
    new_U4024, new_U4025, new_U4026, new_U4027, new_U4028, new_U4029,
    new_U4030, new_U4031, new_U4032, new_U4033, new_U4034, new_U4035,
    new_U4036, new_U4037, new_U4038, new_U4039, new_U4040, new_U4041,
    new_U4042, new_U4043, new_U4044, new_U4045, new_U4046, new_U4047,
    new_U4048, new_U4049, new_U4050, new_U4051, new_U4052, new_U4053,
    new_U4054, new_U4055, new_U4056, new_U4057, new_U4058, new_U4059,
    new_U4060, new_U4061, new_U4062, new_U4063, new_U4064, new_U4065,
    new_U4066, new_U4067, new_U4068, new_U4069, new_U4070, new_U4071,
    new_U4072, new_U4073, new_U4074, new_U4075, new_U4076, new_U4077,
    new_U4078, new_U4079, new_U4080, new_U4081, new_U4082, new_U4083,
    new_U4084, new_U4085, new_U4086, new_U4087, new_U4088, new_U4089,
    new_U4090, new_U4091, new_U4092, new_U4093, new_U4094, new_U4095,
    new_U4096, new_U4097, new_U4098, new_U4099, new_U4100, new_U4101,
    new_U4102, new_U4103, new_U4104, new_U4105, new_U4106, new_U4107,
    new_U4108, new_U4109, new_U4110, new_U4111, new_U4112, new_U4113,
    new_U4114, new_U4115, new_U4116, new_U4117, new_U4118, new_U4119,
    new_U4120, new_U4121, new_U4122, new_U4123, new_U4124, new_U4125,
    new_U4126, new_U4127, new_U4128, new_U4129, new_U4130, new_U4131,
    new_U4132, new_U4133, new_U4134, new_U4135, new_U4136, new_U4137,
    new_U4138, new_U4139, new_U4140, new_U4141, new_U4142, new_U4143,
    new_U4144, new_U4145, new_U4146, new_U4147, new_U4148, new_U4149,
    new_U4150, new_U4151, new_U4152, new_U4153, new_U4154, new_U4155,
    new_U4156, new_U4157, new_U4158, new_U4159, new_U4160, new_U4161,
    new_U4162, new_U4163, new_U4164, new_U4165, new_U4166, new_U4167,
    new_U4168, new_U4169, new_U4170, new_U4171, new_U4172, new_U4173,
    new_U4174, new_U4175, new_U4176, new_U4177, new_U4178, new_U4179,
    new_U4180, new_U4181, new_U4182, new_U4183, new_U4184, new_U4185,
    new_U4186, new_U4187, new_U4188, new_U4189, new_U4190, new_U4191,
    new_U4192, new_U4193, new_U4194, new_U4195, new_U4196, new_U4197,
    new_U4198, new_U4199, new_U4200, new_U4201, new_U4202, new_U4203,
    new_U4204, new_U4205, new_U4206, new_U4207, new_U4208, new_U4209,
    new_U4210, new_U4211, new_U4212, new_U4213, new_U4214, new_U4215,
    new_U4216, new_U4217, new_U4218, new_U4219, new_U4220, new_U4221,
    new_U4222, new_U4223, new_U4224, new_U4225, new_U4226, new_U4227,
    new_U4228, new_U4229, new_U4230, new_U4231, new_U4232, new_U4233,
    new_U4234, new_U4235, new_U4236, new_U4237, new_U4238, new_U4239,
    new_U4240, new_U4241, new_U4242, new_U4243, new_U4244, new_U4245,
    new_U4246, new_U4247, new_U4248, new_U4249, new_U4250, new_U4251,
    new_U4252, new_U4253, new_U4254, new_U4255, new_U4256, new_U4257,
    new_U4258, new_U4259, new_U4260, new_U4261, new_U4262, new_U4263,
    new_U4264, new_U4265, new_U4266, new_U4267, new_U4268, new_U4269,
    new_U4270, new_U4271, new_U4272, new_U4273, new_U4274, new_U4275,
    new_U4276, new_U4277, new_U4278, new_U4279, new_U4280, new_U4281,
    new_U4282, new_U4283, new_U4284, new_U4285, new_U4286, new_U4287,
    new_U4288, new_U4289, new_U4290, new_U4291, new_U4292, new_U4293,
    new_U4294, new_U4295, new_U4296, new_U4297, new_U4298, new_U4299,
    new_U4300, new_U4301, new_U4302, new_U4303, new_U4304, new_U4305,
    new_U4306, new_U4307, new_U4308, new_U4309, new_U4310, new_U4311,
    new_U4312, new_U4313, new_U4314, new_U4315, new_U4316, new_U4317,
    new_U4318, new_U4319, new_U4320, new_U4321, new_U4322, new_U4323,
    new_U4324, new_U4325, new_U4326, new_U4327, new_U4328, new_U4329,
    new_U4330, new_U4331, new_U4332, new_U4333, new_U4334, new_U4335,
    new_U4336, new_U4337, new_U4338, new_U4339, new_U4340, new_U4341,
    new_U4342, new_U4343, new_U4344, new_U4345, new_U4346, new_U4347,
    new_U4348, new_U4349, new_U4350, new_U4351, new_U4352, new_U4353,
    new_U4354, new_U4355, new_U4356, new_U4357, new_U4358, new_U4359,
    new_U4360, new_U4361, new_U4362, new_U4363, new_U4364, new_U4365,
    new_U4366, new_U4367, new_U4368, new_U4369, new_U4370, new_U4371,
    new_U4372, new_U4373, new_U4374, new_U4375, new_U4376, new_U4377,
    new_U4378, new_U4379, new_U4380, new_U4381, new_U4382, new_U4383,
    new_U4384, new_U4385, new_U4386, new_U4387, new_U4388, new_U4389,
    new_U4390, new_U4391, new_U4392, new_U4393, new_U4394, new_U4395,
    new_U4396, new_U4397, new_U4398, new_U4399, new_U4400, new_U4401,
    new_U4402, new_U4403, new_U4404, new_U4405, new_U4406, new_U4407,
    new_U4408, new_U4409, new_U4410, new_U4411, new_U4412, new_U4413,
    new_U4414, new_U4415, new_U4416, new_U4417, new_U4418, new_U4419,
    new_U4420, new_U4421, new_U4422, new_U4423, new_U4424, new_U4425,
    new_U4426, new_U4427, new_U4428, new_U4429, new_U4430, new_U4431,
    new_U4432, new_U4433, new_U4434, new_U4435, new_U4436, new_U4437,
    new_U4438, new_U4439, new_U4440, new_U4441, new_U4442, new_U4443,
    new_U4444, new_U4445, new_U4446, new_U4447, new_U4448, new_U4449,
    new_U4450, new_U4451, new_U4452, new_U4453, new_U4454, new_U4455,
    new_U4456, new_U4457, new_U4458, new_U4459, new_U4460, new_U4461,
    new_U4462, new_U4463, new_U4464, new_U4465, new_U4466, new_U4467,
    new_U4468, new_U4469, new_U4470, new_U4471, new_U4472, new_U4473,
    new_U4474, new_U4475, new_U4476, new_U4477, new_U4478, new_U4479,
    new_U4480, new_U4481, new_U4482, new_U4483, new_U4484, new_U4485,
    new_U4486, new_U4487, new_U4488, new_U4489, new_U4490, new_U4491,
    new_U4492, new_U4493, new_U4494, new_U4495, new_U4496, new_U4497,
    new_U4498, new_U4499, new_U4500, new_U4501, new_U4502, new_U4503,
    new_U4504, new_U4505, new_U4506, new_U4507, new_U4508, new_U4509,
    new_U4510, new_U4511, new_U4512, new_U4513, new_U4514, new_U4515,
    new_U4516, new_U4517, new_U4518, new_U4519, new_U4520, new_U4521,
    new_U4522, new_U4523, new_U4524, new_U4525, new_U4526, new_U4527,
    new_U4528, new_U4529, new_U4530, new_U4531, new_U4532, new_U4533,
    new_U4534, new_U4535, new_U4536, new_U4537, new_U4538, new_U4539,
    new_U4540, new_U4541, new_U4542, new_U4543, new_U4544, new_U4545,
    new_U4546, new_U4547, new_U4548, new_U4549, new_U4550, new_U4551,
    new_U4552, new_U4553, new_U4554, new_U4555, new_U4556, new_U4557,
    new_U4558, new_U4559, new_U4560, new_U4561, new_U4562, new_U4563,
    new_U4564, new_U4565, new_U4566, new_U4567, new_U4568, new_U4569,
    new_U4570, new_U4571, new_U4572, new_U4573, new_U4574, new_U4575,
    new_U4576, new_U4577, new_U4578, new_U4579, new_U4580, new_U4581,
    new_U4582, new_U4583, new_U4584, new_U4585, new_U4586, new_U4587,
    new_U4588, new_U4589, new_U4590, new_U4591, new_U4592, new_U4593,
    new_U4594, new_U4595, new_U4596, new_U4597, new_U4598, new_U4599,
    new_U4600, new_U4601, new_U4602, new_U4603, new_U4604, new_U4605,
    new_U4606, new_U4607, new_U4608, new_U4609, new_U4610, new_U4611,
    new_U4612, new_U4613, new_U4614, new_U4615, new_U4616, new_U4617,
    new_U4618, new_U4619, new_U4620, new_U4621, new_U4622, new_U4623,
    new_U4624, new_U4625, new_U4626, new_U4627, new_U4628, new_U4629,
    new_U4630, new_U4631, new_U4632, new_U4633, new_U4634, new_U4635,
    new_U4636, new_U4637, new_U4638, new_U4639, new_U4640, new_U4641,
    new_U4642, new_U4643, new_U4644, new_U4645, new_U4646, new_U4647,
    new_U4648, new_U4649, new_U4650, new_U4651, new_U4652, new_U4653,
    new_U4654, new_U4655, new_U4656, new_U4657, new_U4658, new_U4659,
    new_U4660, new_U4661, new_U4662, new_U4663, new_U4664, new_U4665,
    new_U4666, new_U4667, new_U4668, new_U4669, new_U4670, new_U4671,
    new_U4672, new_U4673, new_U4674, new_U4675, new_U4676, new_U4677,
    new_U4678, new_U4679, new_U4680, new_U4681, new_U4682, new_U4683,
    new_U4684, new_U4685, new_U4686, new_U4687, new_U4688, new_U4689,
    new_U4690, new_U4691, new_U4692, new_U4693, new_U4694, new_U4695,
    new_U4696, new_U4697, new_U4698, new_U4699, new_U4700, new_U4701,
    new_U4702, new_U4703, new_U4704, new_U4705, new_U4706, new_U4707,
    new_U4708, new_U4709, new_U4710, new_U4711, new_U4712, new_U4713,
    new_U4714, new_U4715, new_U4716, new_U4717, new_U4718, new_U4719,
    new_U4720, new_U4721, new_U4722, new_U4723, new_U4724, new_U4725,
    new_U4726, new_U4727, new_U4728, new_U4729, new_U4730, new_U4731,
    new_U4732, new_U4733, new_U4734, new_U4735, new_U4736, new_U4737,
    new_U4738, new_U4739, new_U4740, new_U4741, new_U4742, new_U4743,
    new_U4744, new_U4745, new_U4746, new_U4747, new_U4748, new_U4749,
    new_U4750, new_U4751, new_U4752, new_U4753, new_U4754, new_U4755,
    new_U4756, new_U4757, new_U4758, new_U4759, new_U4760, new_U4761,
    new_U4762, new_U4763, new_U4764, new_U4765, new_U4766, new_U4767,
    new_U4768, new_U4769, new_U4770, new_U4771, new_U4772, new_U4773,
    new_U4774, new_U4775, new_U4776, new_U4777, new_U4778, new_U4779,
    new_U4780, new_U4781, new_U4782, new_U4783, new_U4784, new_U4785,
    new_U4786, new_U4787, new_U4788, new_U4789, new_U4790, new_U4791,
    new_U4792, new_U4793, new_U4794, new_U4795, new_U4796, new_U4797,
    new_U4798, new_U4799, new_U4800, new_U4801, new_U4802, new_U4803,
    new_U4804, new_U4805, new_U4806, new_U4807, new_U4808, new_U4809,
    new_U4810, new_U4811, new_U4812, new_U4813, new_U4814, new_U4815,
    new_U4816, new_U4817, new_U4818, new_U4819, new_U4820, new_U4821,
    new_U4822, new_U4823, new_U4824, new_U4825, new_U4826, new_U4827,
    new_U4828, new_U4829, new_U4830, new_U4831, new_U4832, new_U4833,
    new_U4834, new_U4835, new_U4836, new_U4837, new_U4838, new_U4839,
    new_U4840, new_U4841, new_U4842, new_U4843, new_U4844, new_U4845,
    new_U4846, new_U4847, new_U4848, new_U4849, new_U4850, new_U4851,
    new_U4852, new_U4853, new_U4854, new_U4855, new_U4856, new_U4857,
    new_U4858, new_U4859, new_U4860, new_U4861, new_U4862, new_U4863,
    new_U4864, new_U4865, new_U4866, new_U4867, new_U4868, new_U4869,
    new_U4870, new_U4871, new_U4872, new_U4873, new_U4874, new_U4875,
    new_U4876, new_U4877, new_U4878, new_U4879, new_U4880, new_U4881,
    new_U4882, new_U4883, new_U4884, new_U4885, new_U4886, new_U4887,
    new_U4888, new_U4889, new_U4890, new_U4891, new_U4892, new_U4893,
    new_U4894, new_U4895, new_U4896, new_U4897, new_U4898, new_U4899,
    new_U4900, new_U4901, new_U4902, new_U4903, new_U4904, new_U4905,
    new_U4906, new_U4907, new_U4908, new_U4909, new_U4910, new_U4911,
    new_U4912, new_U4913, new_U4914, new_U4915, new_U4916, new_U4917,
    new_U4918, new_U4919, new_U4920, new_U4921, new_U4922, new_U4923,
    new_U4924, new_U4925, new_U4926, new_U4927, new_U4928, new_U4929,
    new_U4930, new_U4931, new_U4932, new_U4933, new_U4934, new_U4935,
    new_U4936, new_U4937, new_U4938, new_U4939, new_U4940, new_U4941,
    new_U4942, new_U4943, new_U4944, new_U4945, new_U4946, new_U4947,
    new_U4948, new_U4949, new_U4950, new_U4951, new_U4952, new_U4953,
    new_U4954, new_U4955, new_U4956, new_U4957, new_U4958, new_U4959,
    new_U4960, new_U4961, new_U4962, new_U4963, new_U4964, new_U4965,
    new_U4966, new_U4967, new_U4968, new_U4969, new_U4970, new_U4971,
    new_U4972, new_U4973, new_U4974, new_U4975, new_U4976, new_U4977,
    new_U4978, new_U4979, new_U4980, new_U4981, new_U4982, new_U4983,
    new_U4984, new_U4985, new_U4986, new_U4987, new_U4988, new_U4989,
    new_U4990, new_U4991, new_U4992, new_U4993, new_U4994, new_U4995,
    new_U4996, new_U4997, new_U4998, new_U4999, new_U5000, new_U5001,
    new_U5002, new_U5003, new_U5004, new_U5005, new_U5006, new_U5007,
    new_U5008, new_U5009, new_U5010, new_U5011, new_U5012, new_U5013,
    new_U5014, new_U5015, new_U5016, new_U5017, new_U5018, new_U5019,
    new_U5020, new_U5021, new_U5022, new_U5023, new_U5024, new_U5025,
    new_U5026, new_U5027, new_U5028, new_U5029, new_U5030, new_U5031,
    new_U5032, new_U5033, new_U5034, new_U5035, new_U5036, new_U5037,
    new_U5038, new_U5039, new_U5040, new_U5041, new_U5042, new_U5043,
    new_U5044, new_U5045, new_U5046, new_U5047, new_U5048, new_U5049,
    new_U5050, new_U5051, new_U5052, new_U5053, new_U5054, new_U5055,
    new_U5056, new_U5057, new_U5058, new_U5059, new_U5060, new_U5061,
    new_U5062, new_U5063, new_U5064, new_U5065, new_U5066, new_U5067,
    new_U5068, new_U5069, new_U5070, new_U5071, new_U5072, new_U5073,
    new_U5074, new_U5075, new_U5076, new_U5077, new_U5078, new_U5079,
    new_U5080, new_U5081, new_U5082, new_U5083, new_U5084, new_U5085,
    new_U5086, new_U5087, new_U5088, new_U5089, new_U5090, new_U5091,
    new_U5092, new_U5093, new_U5094, new_U5095, new_U5096, new_U5097,
    new_U5098, new_U5099, new_U5100, new_U5101, new_U5102, new_U5103,
    new_U5104, new_U5105, new_U5106, new_U5107, new_U5108, new_U5109,
    new_U5110, new_U5111, new_U5112, new_U5113, new_U5114, new_U5115,
    new_U5116, new_U5117, new_U5118, new_U5119, new_U5120, new_U5121,
    new_U5122, new_U5123, new_U5124, new_U5125, new_U5126, new_U5127,
    new_U5128, new_U5129, new_U5130, new_U5131, new_U5132, new_U5133,
    new_U5134, new_U5135, new_U5136, new_U5137, new_U5138, new_U5139,
    new_U5140, new_U5141, new_U5142, new_U5143, new_U5144, new_U5145,
    new_U5146, new_U5147, new_U5148, new_U5149, new_U5150, new_U5151,
    new_U5152, new_U5153, new_U5154, new_U5155, new_U5156, new_U5157,
    new_U5158, new_U5159, new_U5160, new_U5161, new_U5162, new_U5163,
    new_U5164, new_U5165, new_U5166, new_U5167, new_U5168, new_U5169,
    new_U5170, new_U5171, new_U5172, new_U5173, new_U5174, new_U5175,
    new_U5176, new_U5177, new_U5178, new_U5179, new_U5180, new_U5181,
    new_U5182, new_U5183, new_U5184, new_U5185, new_U5186, new_U5187,
    new_U5188, new_U5189, new_U5190, new_U5191, new_U5192, new_U5193,
    new_U5194, new_U5195, new_U5196, new_U5197, new_U5198, new_U5199,
    new_U5200, new_U5201, new_U5202, new_U5203, new_U5204, new_U5205,
    new_U5206, new_U5207, new_U5208, new_U5209, new_U5210, new_U5211,
    new_U5212, new_U5213, new_U5214, new_U5215, new_U5216, new_U5217,
    new_U5218, new_U5219, new_U5220, new_U5221, new_U5222, new_U5223,
    new_U5224, new_U5225, new_U5226, new_U5227, new_U5228, new_U5229,
    new_U5230, new_U5231, new_U5232, new_U5233, new_U5234, new_U5235,
    new_U5236, new_U5237, new_U5238, new_U5239, new_U5240, new_U5241,
    new_U5242, new_U5243, new_U5244, new_U5245, new_U5246, new_U5247,
    new_U5248, new_U5249, new_U5250, new_U5251, new_U5252, new_U5253,
    new_U5254, new_U5255, new_U5256, new_U5257, new_U5258, new_U5259,
    new_U5260, new_U5261, new_U5262, new_U5263, new_U5264, new_U5265,
    new_U5266, new_U5267, new_U5268, new_U5269, new_U5270, new_U5271,
    new_U5272, new_U5273, new_U5274, new_U5275, new_U5276, new_U5277,
    new_U5278, new_U5279, new_U5280, new_U5281, new_U5282, new_U5283,
    new_U5284, new_U5285, new_U5286, new_U5287, new_U5288, new_U5289,
    new_U5290, new_U5291, new_U5292, new_U5293, new_U5294, new_U5295,
    new_U5296, new_U5297, new_U5298, new_U5299, new_U5300, new_U5301,
    new_U5302, new_U5303, new_U5304, new_U5305, new_U5306, new_U5307,
    new_U5308, new_U5309, new_U5310, new_U5311, new_U5312, new_U5313,
    new_U5314, new_U5315, new_U5316, new_U5317, new_U5318, new_U5319,
    new_U5320, new_U5321, new_U5322, new_U5323, new_U5324, new_U5325,
    new_U5326, new_U5327, new_U5328, new_U5329, new_U5330, new_U5331,
    new_U5332, new_U5333, new_U5334, new_U5335, new_U5336, new_U5337,
    new_U5338, new_U5339, new_U5340, new_U5341, new_U5342, new_U5343,
    new_U5344, new_U5345, new_U5346, new_U5347, new_U5348, new_U5349,
    new_U5350, new_U5351, new_U5352, new_U5353, new_U5354, new_U5355,
    new_U5356, new_U5357, new_U5358, new_U5359, new_U5360, new_U5361,
    new_U5362, new_U5363, new_U5364, new_U5365, new_U5366, new_U5367,
    new_U5368, new_U5369, new_U5370, new_U5371, new_U5372, new_U5373,
    new_U5374, new_U5375, new_U5376, new_U5377, new_U5378, new_U5379,
    new_U5380, new_U5381, new_U5382, new_U5383, new_U5384, new_U5385,
    new_U5386, new_U5387, new_U5388, new_U5389, new_U5390, new_U5391,
    new_U5392, new_U5393, new_U5394, new_U5395, new_U5396, new_U5397,
    new_U5398, new_U5399, new_U5400, new_U5401, new_U5402, new_U5403,
    new_U5404, new_U5405, new_U5406, new_U5407, new_U5408, new_U5409,
    new_U5410, new_U5411, new_U5412, new_U5413, new_U5414, new_U5415,
    new_U5416, new_U5417, new_U5418, new_U5419, new_U5420, new_U5421,
    new_U5422, new_U5423, new_U5424, new_U5425, new_U5426, new_U5427,
    new_U5428, new_U5429, new_U5430, new_U5431, new_U5432, new_U5433,
    new_U5434, new_U5435, new_U5436, new_U5437, new_U5438, new_U5439,
    new_U5440, new_U5441, new_U5442, new_U5443, new_U5444, new_U5445,
    new_U5446, new_U5447, new_U5448, new_U5449, new_U5450, new_U5451,
    new_U5452, new_U5453, new_U5454, new_U5455, new_U5456, new_U5457,
    new_U5458, new_U5459, new_U5460, new_U5461, new_U5462, new_U5463,
    new_U5464, new_U5465, new_U5466, new_U5467, new_U5468, new_U5469,
    new_U5470, new_U5471, new_U5472, new_U5473, new_U5474, new_U5475,
    new_U5476, new_U5477, new_U5478, new_U5479, new_U5480, new_U5481,
    new_U5482, new_U5483, new_U5484, new_U5485, new_U5486, new_U5487,
    new_U5488, new_U5489, new_U5490, new_U5491, new_U5492, new_U5493,
    new_U5494, new_U5495, new_U5496, new_U5497, new_U5498, new_U5499,
    new_U5500, new_U5501, new_U5502, new_U5503, new_U5504, new_U5505,
    new_U5506, new_U5507, new_U5508, new_U5509, new_U5510, new_U5511,
    new_U5512, new_U5513, new_U5514, new_U5515, new_U5516, new_U5517,
    new_U5518, new_U5519, new_U5520, new_U5521, new_U5522, new_U5523,
    new_U5524, new_U5525, new_U5526, new_U5527, new_U5528, new_U5529,
    new_U5530, new_U5531, new_U5532, new_U5533, new_U5534, new_U5535,
    new_U5536, new_U5537, new_U5538, new_U5539, new_U5540, new_U5541,
    new_U5542, new_U5543, new_U5544, new_U5545, new_U5546, new_U5547,
    new_U5548, new_U5549, new_U5550, new_U5551, new_U5552, new_U5553,
    new_U5554, new_U5555, new_U5556, new_U5557, new_U5558, new_U5559,
    new_U5560, new_U5561, new_U5562, new_U5563, new_U5564, new_U5565,
    new_U5566, new_U5567, new_U5568, new_U5569, new_U5570, new_U5571,
    new_U5572, new_U5573, new_U5574, new_U5575, new_U5576, new_U5577,
    new_U5578, new_U5579, new_U5580, new_U5581, new_U5582, new_U5583,
    new_U5584, new_U5585, new_U5586, new_U5587, new_U5588, new_U5589,
    new_U5590, new_U5591, new_U5592, new_U5593, new_U5594, new_U5595,
    new_U5596, new_U5597, new_U5598, new_U5599, new_U5600, new_U5601,
    new_U5602, new_U5603, new_U5604, new_U5605, new_U5606, new_U5607,
    new_U5608, new_U5609, new_U5610, new_U5611, new_U5612, new_U5613,
    new_U5614, new_U5615, new_U5616, new_U5617, new_U5618, new_U5619,
    new_U5620, new_U5621, new_U5622, new_U5623, new_U5624, new_U5625,
    new_U5626, new_U5627, new_U5628, new_U5629, new_U5630, new_U5631,
    new_U5632, new_U5633, new_U5634, new_U5635, new_U5636, new_U5637,
    new_U5638, new_U5639, new_U5640, new_U5641, new_U5642, new_U5643,
    new_U5644, new_U5645, new_U5646, new_U5647, new_U5648, new_U5649,
    new_U5650, new_U5651, new_U5652, new_U5653, new_U5654, new_U5655,
    new_U5656, new_U5657, new_U5658, new_U5659, new_U5660, new_U5661,
    new_U5662, new_U5663, new_U5664, new_U5665, new_U5666, new_U5667,
    new_U5668, new_U5669, new_U5670, new_U5671, new_U5672, new_U5673,
    new_U5674, new_U5675, new_U5676, new_U5677, new_U5678, new_U5679,
    new_U5680, new_U5681, new_U5682, new_U5683, new_U5684, new_U5685,
    new_U5686, new_U5687, new_U5688, new_U5689, new_U5690, new_U5691,
    new_U5692, new_U5693, new_U5694, new_U5695, new_U5696, new_U5697,
    new_U5698, new_U5699, new_U5700, new_U5701, new_U5702, new_U5703,
    new_U5704, new_U5705, new_U5706, new_U5707, new_U5708, new_U5709,
    new_U5710, new_U5711, new_U5712, new_U5713, new_U5714, new_U5715,
    new_U5716, new_U5717, new_U5718, new_U5719, new_U5720, new_U5721,
    new_U5722, new_U5723, new_U5724, new_U5725, new_U5726, new_U5727,
    new_U5728, new_U5729, new_U5730, new_U5731, new_U5732, new_U5733,
    new_U5734, new_U5735, new_U5736, new_U5737, new_U5738, new_U5739,
    new_U5740, new_U5741, new_U5742, new_U5743, new_U5744, new_U5745,
    new_U5746, new_U5747, new_U5748, new_U5749, new_U5750, new_U5751,
    new_U5752, new_U5753, new_U5754, new_U5755, new_U5756, new_U5757,
    new_U5758, new_U5759, new_U5760, new_U5761, new_U5762, new_U5763,
    new_U5764, new_U5765, new_U5766, new_U5767, new_U5768, new_U5769,
    new_U5770, new_U5771, new_U5772, new_U5773, new_U5774, new_U5775,
    new_U5776, new_U5777, new_U5778, new_U5779, new_U5780, new_U5781,
    new_U5782, new_U5783, new_U5784, new_U5785, new_U5786, new_U5787,
    new_U5788, new_U5789, new_U5790, new_U5791, new_U5792, new_U5793,
    new_U5794, new_U5795, new_U5796, new_U5797, new_U5798, new_U5799,
    new_U5800, new_U5801, new_U5802, new_U5803, new_U5804, new_U5805,
    new_U5806, new_U5807, new_U5808, new_U5809, new_U5810, new_U5811,
    new_U5812, new_U5813, new_U5814, new_U5815, new_U5816, new_U5817,
    new_U5818, new_U5819, new_U5820, new_U5821, new_U5822, new_U5823,
    new_U5824, new_U5825, new_U5826, new_U5827, new_U5828, new_U5829,
    new_U5830, new_U5831, new_U5832, new_U5833, new_U5834, new_U5835,
    new_U5836, new_U5837, new_U5838, new_U5839, new_U5840, new_U5841,
    new_U5842, new_U5843, new_U5844, new_U5845, new_U5846, new_U5847,
    new_U5848, new_U5849, new_U5850, new_U5851, new_U5852, new_U5853,
    new_U5854, new_U5855, new_U5856, new_U5857, new_U5858, new_U5859,
    new_U5860, new_U5861, new_U5862, new_U5863, new_U5864, new_U5865,
    new_U5866, new_U5867, new_U5868, new_U5869, new_U5870, new_U5871,
    new_U5872, new_U5873, new_U5874, new_U5875, new_U5876, new_U5877,
    new_U5878, new_U5879, new_U5880, new_U5881, new_U5882, new_U5883,
    new_U5884, new_U5885, new_U5886, new_U5887, new_U5888, new_U5889,
    new_U5890, new_U5891, new_U5892, new_U5893, new_U5894, new_U5895,
    new_U5896, new_U5897, new_U5898, new_U5899, new_U5900, new_U5901,
    new_U5902, new_U5903, new_U5904, new_U5905, new_U5906, new_U5907,
    new_U5908, new_U5909, new_U5910, new_U5911, new_U5912, new_U5913,
    new_U5914, new_U5915, new_U5916, new_U5917, new_U5918, new_U5919,
    new_U5920, new_U5921, new_U5922, new_U5923, new_U5924, new_U5925,
    new_U5926, new_U5927, new_U5928, new_U5929, new_U5930, new_U5931,
    new_U5932, new_U5933, new_U5934, new_U5935, new_U5936, new_U5937,
    new_U5938, new_U5939, new_U5940, new_U5941, new_U5942, new_U5943,
    new_U5944, new_U5945, new_U5946, new_U5947, new_U5948, new_U5949,
    new_U5950, new_U5951, new_U5952, new_U5953, new_U5954, new_U5955,
    new_U5956, new_U5957, new_U5958, new_U5959, new_U5960, new_U5961,
    new_U5962, new_U5963, new_U5964, new_U5965, new_U5966, new_U5967,
    new_U5968, new_U5969, new_U5970, new_U5971, new_U5972, new_U5973,
    new_U5974, new_U5975, new_U5976, new_U5977, new_U5978, new_U5979,
    new_U5980, new_U5981, new_U5982, new_U5983, new_U5984, new_U5985,
    new_U5986, new_U5987, new_U5988, new_U5989, new_U5990, new_U5991,
    new_U5992, new_U5993, new_U5994, new_U5995, new_U5996, new_U5997,
    new_U5998, new_U5999, new_U6000, new_U6001, new_U6002, new_U6003,
    new_U6004, new_U6005, new_U6006, new_U6007, new_U6008, new_U6009,
    new_U6010, new_U6011, new_U6012, new_U6013, new_U6014, new_U6015,
    new_U6016, new_U6017, new_U6018, new_U6019, new_U6020, new_U6021,
    new_U6022, new_U6023, new_U6024, new_U6025, new_U6026, new_U6027,
    new_U6028, new_U6029, new_U6030, new_U6031, new_U6032, new_U6033,
    new_U6034, new_U6035, new_U6036, new_U6037, new_U6038, new_U6039,
    new_U6040, new_U6041, new_U6042, new_U6043, new_U6044, new_U6045,
    new_U6046, new_U6047, new_U6048, new_U6049, new_U6050, new_U6051,
    new_U6052, new_U6053, new_U6054, new_U6055, new_U6056, new_U6057,
    new_U6058, new_U6059, new_U6060, new_U6061, new_U6062, new_U6063,
    new_U6064, new_U6065, new_U6066, new_U6067, new_U6068, new_U6069,
    new_U6070, new_U6071, new_U6072, new_U6073, new_U6074, new_U6075,
    new_U6076, new_U6077, new_U6078, new_U6079, new_U6080, new_U6081,
    new_U6082, new_U6083, new_U6084, new_U6085, new_U6086, new_U6087,
    new_U6088, new_U6089, new_U6090, new_U6091, new_U6092, new_U6093,
    new_U6094, new_U6095, new_U6096, new_U6097, new_U6098, new_U6099,
    new_U6100, new_U6101, new_U6102, new_U6103, new_U6104, new_U6105,
    new_U6106, new_U6107, new_U6108, new_U6109, new_U6110, new_U6111,
    new_U6112, new_U6113, new_U6114, new_U6115, new_U6116, new_U6117,
    new_U6118, new_U6119, new_U6120, new_U6121, new_U6122, new_U6123,
    new_U6124, new_U6125, new_U6126, new_U6127, new_U6128, new_U6129,
    new_U6130, new_U6131, new_U6132, new_U6133, new_U6134, new_U6135,
    new_U6136, new_U6137, new_U6138, new_U6139, new_U6140, new_U6141,
    new_U6142, new_U6143, new_U6144, new_U6145, new_U6146, new_U6147,
    new_U6148, new_U6149, new_U6150, new_U6151, new_U6152, new_U6153,
    new_U6154, new_U6155, new_U6156, new_U6157, new_U6158, new_U6159,
    new_U6160, new_U6161, new_U6162, new_U6163, new_U6164, new_U6165,
    new_U6166, new_U6167, new_U6168, new_U6169, new_U6170, new_U6171,
    new_U6172, new_U6173, new_U6174, new_U6175, new_U6176, new_U6177,
    new_U6178, new_U6179, new_U6180, new_U6181, new_U6182, new_U6183,
    new_U6184, new_U6185, new_U6186, new_U6187, new_U6188, new_U6189,
    new_U6190, new_U6191, new_U6192, new_U6193, new_U6194, new_U6195,
    new_U6196, new_U6197, new_U6198, new_U6199, new_U6200, new_U6201,
    new_U6202, new_U6203, new_U6204, new_U6205, new_U6206, new_U6207,
    new_U6208, new_U6209, new_U6210, new_U6211, new_U6212, new_U6213,
    new_U6214, new_U6215, new_U6216, new_U6217, new_U6218, new_U6219,
    new_U6220, new_U6221, new_U6222, new_U6223, new_U6224, new_U6225,
    new_U6226, new_U6227, new_U6228, new_U6229, new_U6230, new_U6231,
    new_U6232, new_U6233, new_U6234, new_U6235, new_U6236, new_U6237,
    new_U6238, new_U6239, new_U6240, new_U6241, new_U6242, new_U6243,
    new_U6244, new_U6245, new_U6246, new_U6247, new_U6248, new_U6249,
    new_U6250, new_U6251, new_U6252, new_U6253, new_U6254, new_U6255,
    new_U6256, new_U6257, new_U6258, new_U6259, new_U6260, new_U6261,
    new_U6262, new_U6263, new_U6264, new_U6265, new_U6266, new_U6267,
    new_U6268, new_U6269, new_U6270, new_U6271, new_U6272, new_U6273,
    new_U6274, new_U6275, new_U6276, new_U6277, new_U6278, new_U6279,
    new_U6280, new_U6281, new_U6282, new_U6283, new_U6284, new_U6285,
    new_U6286, new_U6287, new_U6288, new_U6289, new_U6290, new_U6291,
    new_U6292, new_U6293, new_U6294, new_U6295, new_U6296, new_U6297,
    new_U6298, new_U6299, new_U6300, new_U6301, new_U6302, new_U6303,
    new_U6304, new_U6305, new_U6306, new_U6307, new_U6308, new_U6309,
    new_U6310, new_U6311, new_U6312, new_U6313, new_U6314, new_U6315,
    new_U6316, new_U6317, new_U6318, new_U6319, new_U6320, new_U6321,
    new_U6322, new_U6323, new_U6324, new_U6325, new_U6326, new_U6327,
    new_U6328, new_U6329, new_U6330, new_U6331, new_U6332, new_U6333,
    new_U6334, new_U6335, new_U6336, new_U6337, new_U6338, new_U6339,
    new_U6340, new_U6341, new_U6342, new_U6343, new_U6344, new_U6345,
    new_U6346, new_U6347, new_U6348, new_U6349, new_U6350, new_U6351,
    new_U6352, new_U6353, new_U6354, new_U6355, new_U6356, new_U6357,
    new_U6358, new_U6359, new_U6360, new_U6361, new_U6362, new_U6363,
    new_U6364, new_U6365, new_U6366, new_U6367, new_U6368, new_U6369,
    new_U6370, new_U6371, new_U6372, new_U6373, new_U6374, new_U6375,
    new_U6376, new_U6377, new_U6378, new_U6379, new_U6380, new_U6381,
    new_U6382, new_U6383, new_U6384, new_U6385, new_U6386, new_U6387,
    new_U6388, new_U6389, new_U6390, new_U6391, new_U6392, new_U6393,
    new_U6394, new_U6395, new_U6396, new_U6397, new_U6398, new_U6399,
    new_U6400, new_U6401, new_U6402, new_U6403, new_U6404, new_U6405,
    new_U6406, new_U6407, new_U6408, new_U6409, new_U6410, new_U6411,
    new_U6412, new_U6413, new_U6414, new_U6415, new_U6416, new_U6417,
    new_U6418, new_U6419, new_U6420, new_U6421, new_U6422, new_U6423,
    new_U6424, new_U6425, new_U6426, new_U6427, new_U6428, new_U6429,
    new_U6430, new_U6431, new_U6432, new_U6433, new_U6434, new_U6435,
    new_U6436, new_U6437, new_U6438, new_U6439, new_U6440, new_U6441,
    new_U6442, new_U6443, new_U6444, new_U6445, new_U6446, new_U6447,
    new_U6448, new_U6449, new_U6450, new_U6451, new_U6452, new_U6453,
    new_U6454, new_U6455, new_U6456, new_U6457, new_U6458, new_U6459,
    new_U6460, new_U6461, new_U6462, new_U6463, new_U6464, new_U6465,
    new_U6466, new_U6467, new_U6468, new_U6469, new_U6470, new_U6471,
    new_U6472, new_U6473, new_U6474, new_U6475, new_U6476, new_U6477,
    new_U6478, new_U6479, new_U6480, new_U6481, new_U6482, new_U6483,
    new_U6484, new_U6485, new_U6486, new_U6487, new_U6488, new_U6489,
    new_U6490, new_U6491, new_U6492, new_U6493, new_U6494, new_U6495,
    new_U6496, new_U6497, new_U6498, new_U6499, new_U6500, new_U6501,
    new_U6502, new_U6503, new_U6504, new_U6505, new_U6506, new_U6507,
    new_U6508, new_U6509, new_U6510, new_U6511, new_U6512, new_U6513,
    new_U6514, new_U6515, new_U6516, new_U6517, new_U6518, new_U6519,
    new_U6520, new_U6521, new_U6522, new_U6523, new_U6524, new_U6525,
    new_U6526, new_U6527, new_U6528, new_U6529, new_U6530, new_U6531,
    new_U6532, new_U6533, new_U6534, new_U6535, new_U6536, new_U6537,
    new_U6538, new_U6539, new_U6540, new_U6541, new_U6542, new_U6543,
    new_U6544, new_U6545, new_U6546, new_U6547, new_U6548, new_U6549,
    new_U6550, new_U6551, new_U6552, new_U6553, new_U6554, new_U6555,
    new_U6556, new_U6557, new_U6558, new_U6559, new_U6560, new_U6561,
    new_U6562, new_U6563, new_U6564, new_U6565, new_U6566, new_U6567,
    new_U6568, new_U6569, new_U6570, new_U6571, new_U6572, new_U6573,
    new_U6574, new_U6575, new_U6576, new_U6577, new_U6578, new_U6579,
    new_U6580, new_U6581, new_U6582, new_U6583, new_U6584, new_U6585,
    new_U6586, new_U6587, new_U6588, new_U6589, new_U6590, new_U6591,
    new_U6592, new_U6593, new_U6594, new_U6595, new_U6596, new_U6597,
    new_U6598, new_U6599, new_U6600, new_U6601, new_U6602, new_U6603,
    new_U6604, new_U6605, new_U6606, new_U6607, new_U6608, new_U6609,
    new_U6610, new_U6611, new_U6612, new_U6613, new_U6614, new_U6615,
    new_U6616, new_U6617, new_U6618, new_U6619, new_U6620, new_U6621,
    new_U6622, new_U6623, new_U6624, new_U6625, new_U6626, new_U6627,
    new_U6628, new_U6629, new_U6630, new_U6631, new_U6632, new_U6633,
    new_U6634, new_U6635, new_U6636, new_U6637, new_U6638, new_U6639,
    new_U6640, new_U6641, new_U6642, new_U6643, new_U6644, new_U6645,
    new_U6646, new_U6647, new_U6648, new_U6649, new_U6650, new_U6651,
    new_U6652, new_U6653, new_U6654, new_U6655, new_U6656, new_U6657,
    new_U6658, new_U6659, new_U6660, new_U6661, new_U6662, new_U6663,
    new_U6664, new_U6665, new_U6666, new_U6667, new_U6668, new_U6669,
    new_U6670, new_U6671, new_U6672, new_U6673, new_U6674, new_U6675,
    new_U6676, new_U6677, new_U6678, new_U6679, new_U6680, new_U6681,
    new_U6682, new_U6683, new_U6684, new_U6685, new_U6686, new_U6687,
    new_U6688, new_U6689, new_U6690, new_U6691, new_U6692, new_U6693,
    new_U6694, new_U6695, new_U6696, new_U6697, new_U6698, new_U6699,
    new_U6700, new_U6701, new_U6702, new_U6703, new_U6704, new_U6705,
    new_U6706, new_U6707, new_U6708, new_U6709, new_U6710, new_U6711,
    new_U6712, new_U6713, new_U6714, new_U6715, new_U6716, new_U6717,
    new_U6718, new_U6719, new_U6720, new_U6721, new_U6722, new_U6723,
    new_U6724, new_U6725, new_U6726, new_U6727, new_U6728, new_U6729,
    new_U6730, new_U6731, new_U6732, new_U6733, new_U6734, new_U6735,
    new_U6736, new_U6737, new_U6738, new_U6739, new_U6740, new_U6741,
    new_U6742, new_U6743, new_U6744, new_U6745, new_U6746, new_U6747,
    new_U6748, new_U6749, new_U6750, new_U6751, new_U6752, new_U6753,
    new_U6754, new_U6755, new_U6756, new_U6757, new_U6758, new_U6759,
    new_U6760, new_U6761, new_U6762, new_U6763, new_U6764, new_U6765,
    new_U6766, new_U6767, new_U6768, new_U6769, new_U6770, new_U6771,
    new_U6772, new_U6773, new_U6774, new_U6775, new_U6776, new_U6777,
    new_U6778, new_U6779, new_U6780, new_U6781, new_U6782, new_U6783,
    new_U6784, new_U6785, new_U6786, new_U6787, new_U6788, new_U6789,
    new_U6790, new_U6791, new_U6792, new_U6793, new_U6794, new_U6795,
    new_U6796, new_U6797, new_U6798, new_U6799, new_U6800, new_U6801,
    new_U6802, new_U6803, new_U6804, new_U6805, new_U6806, new_U6807,
    new_U6808, new_U6809, new_U6810, new_U6811, new_U6812, new_U6813,
    new_U6814, new_U6815, new_U6816, new_U6817, new_U6818, new_U6819,
    new_U6820, new_U6821, new_U6822, new_U6823, new_U6824, new_U6825,
    new_U6826, new_U6827, new_U6828, new_U6829, new_U6830, new_U6831,
    new_U6832, new_U6833, new_U6834, new_U6835, new_U6836, new_U6837,
    new_U6838, new_U6839, new_U6840, new_U6841, new_U6842, new_U6843,
    new_U6844, new_U6845, new_U6846, new_U6847, new_U6848, new_U6849,
    new_U6850, new_U6851, new_U6852, new_U6853, new_U6854, new_U6855,
    new_U6856, new_U6857, new_U6858, new_U6859, new_U6860, new_U6861,
    new_U6862, new_U6863, new_U6864, new_U6865, new_U6866, new_U6867,
    new_U6868, new_U6869, new_U6870, new_U6871, new_U6872, new_U6873,
    new_U6874, new_U6875, new_U6876, new_U6877, new_U6878, new_U6879,
    new_U6880, new_U6881, new_U6882, new_U6883, new_U6884, new_U6885,
    new_U6886, new_U6887, new_U6888, new_U6889, new_U6890, new_U6891,
    new_U6892, new_U6893, new_U6894, new_U6895, new_U6896, new_U6897,
    new_U6898, new_U6899, new_U6900, new_U6901, new_U6902, new_U6903,
    new_U6904, new_U6905, new_U6906, new_U6907, new_U6908, new_U6909,
    new_U6910, new_U6911, new_U6912, new_U6913, new_U6914, new_U6915,
    new_U6916, new_U6917, new_U6918, new_U6919, new_U6920, new_U6921,
    new_U6922, new_U6923, new_U6924, new_U6925, new_U6926, new_U6927,
    new_U6928, new_U6929, new_U6930, new_U6931, new_U6932, new_U6933,
    new_U6934, new_U6935, new_U6936, new_U6937, new_U6938, new_U6939,
    new_U6940, new_U6941, new_U6942, new_U6943, new_U6944, new_U6945,
    new_U6946, new_U6947, new_U6948, new_U6949, new_U6950, new_U6951,
    new_U6952, new_U6953, new_U6954, new_U6955, new_U6956, new_U6957,
    new_U6958, new_U6959, new_U6960, new_U6961, new_U6962, new_U6963,
    new_U6964, new_U6965, new_U6966, new_U6967, new_U6968, new_U6969,
    new_U6970, new_U6971, new_U6972, new_U6973, new_U6974, new_U6975,
    new_U6976, new_U6977, new_U6978, new_U6979, new_U6980, new_U6981,
    new_U6982, new_U6983, new_U6984, new_U6985, new_U6986, new_U6987,
    new_U6988, new_U6989, new_U6990, new_U6991, new_U6992, new_U6993,
    new_U6994, new_U6995, new_U6996, new_U6997, new_U6998, new_U6999,
    new_U7000, new_U7001, new_U7002, new_U7003, new_U7004, new_U7005,
    new_U7006, new_U7007, new_U7008, new_U7009, new_U7010, new_U7011,
    new_U7012, new_U7013, new_U7014, new_U7015, new_U7016, new_U7017,
    new_U7018, new_U7019, new_U7020, new_U7021, new_U7022, new_U7023,
    new_U7024, new_U7025, new_U7026, new_U7027, new_U7028, new_U7029,
    new_U7030, new_U7031, new_U7032, new_U7033, new_U7034, new_U7035,
    new_U7036, new_U7037, new_U7038, new_U7039, new_U7040, new_U7041,
    new_U7042, new_U7043, new_U7044, new_U7045, new_U7046, new_U7047,
    new_U7048, new_U7049, new_U7050, new_U7051, new_U7052, new_U7053,
    new_U7054, new_U7055, new_U7056, new_U7057, new_U7058, new_U7059,
    new_U7060, new_U7061, new_U7062, new_U7063, new_U7064, new_U7065,
    new_U7066, new_U7067, new_U7068, new_U7069, new_U7070, new_U7071,
    new_U7072, new_U7073, new_U7074, new_U7075, new_U7076, new_U7077,
    new_U7078, new_U7079, new_U7080, new_U7081, new_U7082, new_U7083,
    new_U7084, new_U7085, new_U7086, new_U7087, new_U7088, new_U7089,
    new_U7090, new_U7091, new_U7092, new_U7093, new_U7094, new_U7095,
    new_U7096, new_U7097, new_U7098, new_U7099, new_U7100, new_U7101,
    new_U7102, new_U7103, new_U7104, new_U7105, new_U7106, new_U7107,
    new_U7108, new_U7109, new_U7110, new_U7111, new_U7112, new_U7113,
    new_U7114, new_U7115, new_U7116, new_U7117, new_U7118, new_U7119,
    new_U7120, new_U7121, new_U7122, new_U7123, new_U7124, new_U7125,
    new_U7126, new_U7127, new_U7128, new_U7129, new_U7130, new_U7131,
    new_U7132, new_U7133, new_U7134, new_U7135, new_U7136, new_U7137,
    new_U7138, new_U7139, new_U7140, new_U7141, new_U7142, new_U7143,
    new_U7144, new_U7145, new_U7146, new_U7147, new_U7148, new_U7149,
    new_U7150, new_U7151, new_U7152, new_U7153, new_U7154, new_U7155,
    new_U7156, new_U7157, new_U7158, new_U7159, new_U7160, new_U7161,
    new_U7162, new_U7163, new_U7164, new_U7165, new_U7166, new_U7167,
    new_U7168, new_U7169, new_U7170, new_U7171, new_U7172, new_U7173,
    new_U7174, new_U7175, new_U7176, new_U7177, new_U7178, new_U7179,
    new_U7180, new_U7181, new_U7182, new_U7183, new_U7184, new_U7185,
    new_U7186, new_U7187, new_U7188, new_U7189, new_U7190, new_U7191,
    new_U7192, new_U7193, new_U7194, new_U7195, new_U7196, new_U7197,
    new_U7198, new_U7199, new_U7200, new_U7201, new_U7202, new_U7203,
    new_U7204, new_U7205, new_U7206, new_U7207, new_U7208, new_U7209,
    new_U7210, new_U7211, new_U7212, new_U7213, new_U7214, new_U7215,
    new_U7216, new_U7217, new_U7218, new_U7219, new_U7220, new_U7221,
    new_U7222, new_U7223, new_U7224, new_U7225, new_U7226, new_U7227,
    new_U7228, new_U7229, new_U7230, new_U7231, new_U7232, new_U7233,
    new_U7234, new_U7235, new_U7236, new_U7237, new_U7238, new_U7239,
    new_U7240, new_U7241, new_U7242, new_U7243, new_U7244, new_U7245,
    new_U7246, new_U7247, new_U7248, new_U7249, new_U7250, new_U7251,
    new_U7252, new_U7253, new_U7254, new_U7255, new_U7256, new_U7257,
    new_U7258, new_U7259, new_U7260, new_U7261, new_U7262, new_U7263,
    new_U7264, new_U7265, new_U7266, new_U7267, new_U7268, new_U7269,
    new_U7270, new_U7271, new_U7272, new_U7273, new_U7274, new_U7275,
    new_U7276, new_U7277, new_U7278, new_U7279, new_U7280, new_U7281,
    new_U7282, new_U7283, new_U7284, new_U7285, new_U7286, new_U7287,
    new_U7288, new_U7289, new_U7290, new_U7291, new_U7292, new_U7293,
    new_U7294, new_U7295, new_U7296, new_U7297, new_U7298, new_U7299,
    new_U7300, new_U7301, new_U7302, new_U7303, new_U7304, new_U7305,
    new_U7306, new_U7307, new_U7308, new_U7309, new_U7310, new_U7311,
    new_U7312, new_U7313, new_U7314, new_U7315, new_U7316, new_U7317,
    new_U7318, new_U7319, new_U7320, new_U7321, new_U7322, new_U7323,
    new_U7324, new_U7325, new_U7326, new_U7327, new_U7328, new_U7329,
    new_U7330, new_U7331, new_U7332, new_U7333, new_U7334, new_U7335,
    new_U7336, new_U7337, new_U7338, new_U7339, new_U7340, new_U7341,
    new_U7342, new_U7343, new_U7344, new_U7345, new_U7346, new_U7347,
    new_U7348, new_U7349, new_U7350, new_U7351, new_U7352, new_U7353,
    new_U7354, new_U7355, new_U7356, new_U7357, new_U7358, new_U7359,
    new_U7360, new_U7361, new_U7362, new_U7363, new_U7364, new_U7365,
    new_U7366, new_U7367, new_U7368, new_U7369, new_U7370, new_U7371,
    new_U7372, new_U7373, new_U7374, new_U7375, new_U7376, new_U7377,
    new_U7378, new_U7379, new_U7380, new_U7381, new_U7382, new_U7383,
    new_U7384, new_U7385, new_U7386, new_U7387, new_U7388, new_U7389,
    new_U7390, new_U7391, new_U7392, new_U7393, new_U7394, new_U7395,
    new_U7396, new_U7397, new_U7398, new_U7399, new_U7400, new_U7401,
    new_U7402, new_U7403, new_U7404, new_U7405, new_U7406, new_U7407,
    new_U7408, new_U7409, new_U7410, new_U7411, new_U7412, new_U7413,
    new_U7414, new_U7415, new_U7416, new_U7417, new_U7418, new_U7419,
    new_U7420, new_U7421, new_U7422, new_U7423, new_U7424, new_U7425,
    new_U7426, new_U7427, new_U7428, new_U7429, new_U7430, new_U7431,
    new_U7432, new_U7433, new_U7434, new_U7435, new_U7436, new_U7437,
    new_U7438, new_U7439, new_U7440, new_U7441, new_U7442, new_U7443,
    new_U7444, new_U7445, new_U7446, new_U7447, new_U7448, new_U7449,
    new_U7450, new_U7451, new_U7452, new_U7453, new_U7454, new_U7455,
    new_U7456, new_U7457, new_U7458, new_U7459, new_U7460, new_U7461,
    new_U7462, new_U7463, new_U7464, new_U7465, new_U7466, new_U7467,
    new_U7468, new_U7469, new_U7470, new_U7471, new_U7472, new_U7473,
    new_U7474, new_U7475, new_U7476, new_U7477, new_U7478, new_U7479,
    new_U7480, new_U7481, new_U7482, new_U7483, new_U7484, new_U7485,
    new_U7486, new_U7487, new_U7488, new_U7489, new_U7490, new_U7491,
    new_U7492, new_U7493, new_U7494, new_U7495, new_U7496, new_U7497,
    new_U7498, new_U7499, new_U7500, new_U7501, new_U7502, new_U7503,
    new_U7504, new_U7505, new_U7506, new_U7507, new_U7508, new_U7509,
    new_U7510, new_U7511, new_U7512, new_U7513, new_U7514, new_U7515,
    new_U7516, new_U7517, new_U7518, new_U7519, new_U7520, new_U7521,
    new_U7522, new_U7523, new_U7524, new_U7525, new_U7526, new_U7527,
    new_U7528, new_U7529, new_U7530, new_U7531, new_U7532, new_U7533,
    new_U7534, new_U7535, new_U7536, new_U7537, new_U7538, new_U7539,
    new_U7540, new_U7541, new_U7542, new_U7543, new_U7544, new_U7545,
    new_U7546, new_U7547, new_U7548, new_U7549, new_U7550, new_U7551,
    new_U7552, new_U7553, new_U7554, new_U7555, new_U7556, new_U7557,
    new_U7558, new_U7559, new_U7560, new_U7561, new_U7562, new_U7563,
    new_U7564, new_U7565, new_U7566, new_U7567, new_U7568, new_U7569,
    new_U7570, new_U7571, new_U7572, new_U7573, new_U7574, new_U7575,
    new_U7576, new_U7577, new_U7578, new_U7579, new_U7580, new_U7581,
    new_U7582, new_U7583, new_U7584, new_U7585, new_U7586, new_U7587,
    new_U7588, new_U7589, new_U7590, new_U7591, new_U7592, new_U7593,
    new_U7594, new_U7595, new_U7596, new_U7597, new_U7598, new_U7599,
    new_U7600, new_U7601, new_U7602, new_U7603, new_U7604, new_U7605,
    new_U7606, new_U7607, new_U7608, new_U7609, new_U7610, new_U7611,
    new_U7612, new_U7613, new_U7614, new_U7615, new_U7616, new_U7617,
    new_U7618, new_U7619, new_U7620, new_U7621, new_U7622, new_U7623,
    new_U7624, new_U7625, new_U7626, new_U7627, new_U7628, new_U7629,
    new_U7630, new_U7631, new_U7632, new_U7633, new_U7634, new_U7635,
    new_U7636, new_U7637, new_U7638, new_U7639, new_U7640, new_U7641,
    new_U7642, new_U7643, new_U7644, new_U7645, new_U7646, new_U7647,
    new_U7648, new_U7649, new_U7650, new_U7651, new_U7652, new_U7653,
    new_U7654, new_U7655, new_U7656, new_U7657, new_U7658, new_U7659,
    new_U7660, new_U7661, new_U7662, new_U7663, new_U7664, new_U7665,
    new_U7666, new_U7667, new_U7668, new_U7669, new_U7670, new_U7671,
    new_U7672, new_U7673, new_U7674, new_U7675, new_U7676, new_U7677,
    new_U7678, new_U7679, new_U7680, new_U7681, new_U7682, new_U7683,
    new_U7684, new_U7685, new_U7686, new_U7687, new_U7688, new_U7689,
    new_U7690, new_U7691, new_U7692, new_U7693, new_U7694, new_U7695,
    new_U7696, new_U7697, new_U7698, new_U7699, new_U7700, new_U7701,
    new_U7702, new_U7703, new_U7704, new_U7705, new_U7706, new_U7707,
    new_U7708, new_U7709, new_U7710, new_U7711, new_U7712, new_U7713,
    new_U7714, new_U7715, new_U7716, new_U7717, new_U7718, new_U7719,
    new_U7720, new_U7721, new_U7722, new_U7723, new_U7724, new_U7725,
    new_U7726, new_U7727, new_U7728, new_U7729, new_U7730, new_U7731,
    new_U7732, new_U7733, new_U7734, new_U7735, new_U7736, new_U7737,
    new_U7738, new_U7739, new_U7740, new_U7741, new_U7742, new_U7743,
    new_U7744, new_U7745, new_U7746, new_U7747, new_U7748, new_U7749,
    new_U7750, new_U7751, new_U7752, new_U7753, new_U7754, new_U7755,
    new_U7756, new_U7757, new_U7758, new_U7759, new_U7760, new_U7761,
    new_U7762, new_U7763, new_U7764, new_U7765, new_U7766, new_U7767,
    new_U7768, new_U7769, new_U7770, new_U7771, new_U7772, new_U7773,
    new_U7774, new_U7775, new_U7776, new_U7777, new_U7778, new_U7779,
    new_U7780, new_U7781, new_U7782, new_ADD_515_U178, new_ADD_515_U177,
    new_ADD_515_U176, new_ADD_515_U175, new_ADD_515_U174, new_ADD_515_U173,
    new_ADD_515_U172, new_ADD_515_U171, new_ADD_515_U170, new_ADD_515_U169,
    new_ADD_515_U168, new_ADD_515_U167, new_ADD_515_U166, new_ADD_515_U165,
    new_ADD_515_U164, new_ADD_515_U163, new_ADD_515_U162, new_ADD_515_U161,
    new_ADD_515_U160, new_ADD_515_U159, new_ADD_515_U158, new_ADD_515_U157,
    new_ADD_515_U156, new_ADD_515_U155, new_ADD_515_U154, new_ADD_515_U153,
    new_ADD_515_U152, new_R2027_U5, new_R2027_U6, new_R2027_U7,
    new_R2027_U8, new_R2027_U9, new_R2027_U10, new_R2027_U11,
    new_R2027_U12, new_R2027_U13, new_R2027_U14, new_R2027_U15,
    new_R2027_U16, new_R2027_U17, new_R2027_U18, new_R2027_U19,
    new_R2027_U20, new_R2027_U21, new_R2027_U22, new_R2027_U23,
    new_R2027_U24, new_R2027_U25, new_R2027_U26, new_R2027_U27,
    new_R2027_U28, new_R2027_U29, new_R2027_U30, new_R2027_U31,
    new_R2027_U32, new_R2027_U33, new_R2027_U34, new_R2027_U35,
    new_R2027_U36, new_R2027_U37, new_R2027_U38, new_R2027_U39,
    new_R2027_U40, new_R2027_U41, new_R2027_U42, new_R2027_U43,
    new_R2027_U44, new_R2027_U45, new_R2027_U46, new_R2027_U47,
    new_R2027_U48, new_R2027_U49, new_R2027_U50, new_R2027_U51,
    new_R2027_U52, new_R2027_U53, new_R2027_U54, new_R2027_U55,
    new_R2027_U56, new_R2027_U57, new_R2027_U58, new_R2027_U59,
    new_R2027_U60, new_R2027_U61, new_R2027_U62, new_R2027_U63,
    new_R2027_U64, new_R2027_U65, new_R2027_U66, new_R2027_U67,
    new_R2027_U68, new_R2027_U69, new_R2027_U70, new_R2027_U71,
    new_R2027_U72, new_R2027_U73, new_R2027_U74, new_R2027_U75,
    new_R2027_U76, new_R2027_U77, new_R2027_U78, new_R2027_U79,
    new_R2027_U80, new_R2027_U81, new_R2027_U82, new_R2027_U83,
    new_R2027_U84, new_R2027_U85, new_R2027_U86, new_R2027_U87,
    new_R2027_U88, new_R2027_U89, new_R2027_U90, new_R2027_U91,
    new_R2027_U92, new_R2027_U93, new_R2027_U94, new_R2027_U95,
    new_R2027_U96, new_R2027_U97, new_R2027_U98, new_R2027_U99,
    new_R2027_U100, new_R2027_U101, new_R2027_U102, new_R2027_U103,
    new_R2027_U104, new_R2027_U105, new_R2027_U106, new_R2027_U107,
    new_R2027_U108, new_R2027_U109, new_R2027_U110, new_R2027_U111,
    new_R2027_U112, new_R2027_U113, new_R2027_U114, new_R2027_U115,
    new_R2027_U116, new_R2027_U117, new_R2027_U118, new_R2027_U119,
    new_R2027_U120, new_R2027_U121, new_R2027_U122, new_R2027_U123,
    new_R2027_U124, new_R2027_U125, new_R2027_U126, new_R2027_U127,
    new_R2027_U128, new_R2027_U129, new_R2027_U130, new_R2027_U131,
    new_R2027_U132, new_R2027_U133, new_R2027_U134, new_R2027_U135,
    new_R2027_U136, new_R2027_U137, new_R2027_U138, new_R2027_U139,
    new_R2027_U140, new_R2027_U141, new_R2027_U142, new_R2027_U143,
    new_R2027_U144, new_R2027_U145, new_R2027_U146, new_R2027_U147,
    new_R2027_U148, new_R2027_U149, new_R2027_U150, new_R2027_U151,
    new_R2027_U152, new_R2027_U153, new_R2027_U154, new_R2027_U155,
    new_R2027_U156, new_R2027_U157, new_R2027_U158, new_R2027_U159,
    new_R2027_U160, new_R2027_U161, new_R2027_U162, new_R2027_U163,
    new_R2027_U164, new_R2027_U165, new_R2027_U166, new_R2027_U167,
    new_R2027_U168, new_R2027_U169, new_R2027_U170, new_R2027_U171,
    new_R2027_U172, new_R2027_U173, new_R2027_U174, new_R2027_U175,
    new_R2027_U176, new_R2027_U177, new_R2027_U178, new_R2027_U179,
    new_R2027_U180, new_R2027_U181, new_R2027_U182, new_R2027_U183,
    new_R2027_U184, new_R2027_U185, new_R2027_U186, new_R2027_U187,
    new_R2027_U188, new_R2027_U189, new_R2027_U190, new_R2027_U191,
    new_R2027_U192, new_R2027_U193, new_R2027_U194, new_R2027_U195,
    new_R2027_U196, new_R2027_U197, new_R2027_U198, new_R2027_U199,
    new_R2027_U200, new_R2027_U201, new_R2027_U202, new_R2278_U5,
    new_R2278_U6, new_R2278_U7, new_R2278_U8, new_R2278_U9, new_R2278_U10,
    new_R2278_U11, new_R2278_U12, new_R2278_U13, new_R2278_U14,
    new_R2278_U15, new_R2278_U16, new_R2278_U17, new_R2278_U18,
    new_R2278_U19, new_R2278_U20, new_R2278_U21, new_R2278_U22,
    new_R2278_U23, new_R2278_U24, new_R2278_U25, new_R2278_U26,
    new_R2278_U27, new_R2278_U28, new_R2278_U29, new_R2278_U30,
    new_R2278_U31, new_R2278_U32, new_R2278_U33, new_R2278_U34,
    new_R2278_U35, new_R2278_U36, new_R2278_U37, new_R2278_U38,
    new_R2278_U39, new_R2278_U40, new_R2278_U41, new_R2278_U42,
    new_R2278_U43, new_R2278_U44, new_R2278_U45, new_R2278_U46,
    new_R2278_U47, new_R2278_U48, new_R2278_U49, new_R2278_U50,
    new_R2278_U51, new_R2278_U52, new_R2278_U53, new_R2278_U54,
    new_R2278_U55, new_R2278_U56, new_R2278_U57, new_R2278_U58,
    new_R2278_U59, new_R2278_U60, new_R2278_U61, new_R2278_U62,
    new_R2278_U63, new_R2278_U64, new_R2278_U65, new_R2278_U66,
    new_R2278_U67, new_R2278_U68, new_R2278_U69, new_R2278_U70,
    new_R2278_U71, new_R2278_U72, new_R2278_U73, new_R2278_U74,
    new_R2278_U75, new_R2278_U76, new_R2278_U77, new_R2278_U78,
    new_R2278_U79, new_R2278_U80, new_R2278_U81, new_R2278_U82,
    new_R2278_U83, new_R2278_U84, new_R2278_U85, new_R2278_U86,
    new_R2278_U87, new_R2278_U88, new_R2278_U89, new_R2278_U90,
    new_R2278_U91, new_R2278_U92, new_R2278_U93, new_R2278_U94,
    new_R2278_U95, new_R2278_U96, new_R2278_U97, new_R2278_U98,
    new_R2278_U99, new_R2278_U100, new_R2278_U101, new_R2278_U102,
    new_R2278_U103, new_R2278_U104, new_R2278_U105, new_R2278_U106,
    new_R2278_U107, new_R2278_U108, new_R2278_U109, new_R2278_U110,
    new_R2278_U111, new_R2278_U112, new_R2278_U113, new_R2278_U114,
    new_R2278_U115, new_R2278_U116, new_R2278_U117, new_R2278_U118,
    new_R2278_U119, new_R2278_U120, new_R2278_U121, new_R2278_U122,
    new_R2278_U123, new_R2278_U124, new_R2278_U125, new_R2278_U126,
    new_R2278_U127, new_R2278_U128, new_R2278_U129, new_R2278_U130,
    new_R2278_U131, new_R2278_U132, new_R2278_U133, new_R2278_U134,
    new_R2278_U135, new_R2278_U136, new_R2278_U137, new_R2278_U138,
    new_R2278_U139, new_R2278_U140, new_R2278_U141, new_R2278_U142,
    new_R2278_U143, new_R2278_U144, new_R2278_U145, new_R2278_U146,
    new_R2278_U147, new_R2278_U148, new_R2278_U149, new_R2278_U150,
    new_R2278_U151, new_R2278_U152, new_R2278_U153, new_R2278_U154,
    new_R2278_U155, new_R2278_U156, new_R2278_U157, new_R2278_U158,
    new_R2278_U159, new_R2278_U160, new_R2278_U161, new_R2278_U162,
    new_R2278_U163, new_R2278_U164, new_R2278_U165, new_R2278_U166,
    new_R2278_U167, new_R2278_U168, new_R2278_U169, new_R2278_U170,
    new_R2278_U171, new_R2278_U172, new_R2278_U173, new_R2278_U174,
    new_R2278_U175, new_R2278_U176, new_R2278_U177, new_R2278_U178,
    new_R2278_U179, new_R2278_U180, new_R2278_U181, new_R2278_U182,
    new_R2278_U183, new_R2278_U184, new_R2278_U185, new_R2278_U186,
    new_R2278_U187, new_R2278_U188, new_R2278_U189, new_R2278_U190,
    new_R2278_U191, new_R2278_U192, new_R2278_U193, new_R2278_U194,
    new_R2278_U195, new_R2278_U196, new_R2278_U197, new_R2278_U198,
    new_R2278_U199, new_R2278_U200, new_R2278_U201, new_R2278_U202,
    new_R2278_U203, new_R2278_U204, new_R2278_U205, new_R2278_U206,
    new_R2278_U207, new_R2278_U208, new_R2278_U209, new_R2278_U210,
    new_R2278_U211, new_R2278_U212, new_R2278_U213, new_R2278_U214,
    new_R2278_U215, new_R2278_U216, new_R2278_U217, new_R2278_U218,
    new_R2278_U219, new_R2278_U220, new_R2278_U221, new_R2278_U222,
    new_R2278_U223, new_R2278_U224, new_R2278_U225, new_R2278_U226,
    new_R2278_U227, new_R2278_U228, new_R2278_U229, new_R2278_U230,
    new_R2278_U231, new_R2278_U232, new_R2278_U233, new_R2278_U234,
    new_R2278_U235, new_R2278_U236, new_R2278_U237, new_R2278_U238,
    new_R2278_U239, new_R2278_U240, new_R2278_U241, new_R2278_U242,
    new_R2278_U243, new_R2278_U244, new_R2278_U245, new_R2278_U246,
    new_R2278_U247, new_R2278_U248, new_R2278_U249, new_R2278_U250,
    new_R2278_U251, new_R2278_U252, new_R2278_U253, new_R2278_U254,
    new_R2278_U255, new_R2278_U256, new_R2278_U257, new_R2278_U258,
    new_R2278_U259, new_R2278_U260, new_R2278_U261, new_R2278_U262,
    new_R2278_U263, new_R2278_U264, new_R2278_U265, new_R2278_U266,
    new_R2278_U267, new_R2278_U268, new_R2278_U269, new_R2278_U270,
    new_R2278_U271, new_R2278_U272, new_R2278_U273, new_R2278_U274,
    new_R2278_U275, new_R2278_U276, new_R2278_U277, new_R2278_U278,
    new_R2278_U279, new_R2278_U280, new_R2278_U281, new_R2278_U282,
    new_R2278_U283, new_R2278_U284, new_R2278_U285, new_R2278_U286,
    new_R2278_U287, new_R2278_U288, new_R2278_U289, new_R2278_U290,
    new_R2278_U291, new_R2278_U292, new_R2278_U293, new_R2278_U294,
    new_R2278_U295, new_R2278_U296, new_R2278_U297, new_R2278_U298,
    new_R2278_U299, new_R2278_U300, new_R2278_U301, new_R2278_U302,
    new_R2278_U303, new_R2278_U304, new_R2278_U305, new_R2278_U306,
    new_R2278_U307, new_R2278_U308, new_R2278_U309, new_R2278_U310,
    new_R2278_U311, new_R2278_U312, new_R2278_U313, new_R2278_U314,
    new_R2278_U315, new_R2278_U316, new_R2278_U317, new_R2278_U318,
    new_R2278_U319, new_R2278_U320, new_R2278_U321, new_R2278_U322,
    new_R2278_U323, new_R2278_U324, new_R2278_U325, new_R2278_U326,
    new_R2278_U327, new_R2278_U328, new_R2278_U329, new_R2278_U330,
    new_R2278_U331, new_R2278_U332, new_R2278_U333, new_R2278_U334,
    new_R2278_U335, new_R2278_U336, new_R2278_U337, new_R2278_U338,
    new_R2278_U339, new_R2278_U340, new_R2278_U341, new_R2278_U342,
    new_R2278_U343, new_R2278_U344, new_R2278_U345, new_R2278_U346,
    new_R2278_U347, new_R2278_U348, new_R2278_U349, new_R2278_U350,
    new_R2278_U351, new_R2278_U352, new_R2278_U353, new_R2278_U354,
    new_R2278_U355, new_R2278_U356, new_R2278_U357, new_R2278_U358,
    new_R2278_U359, new_R2278_U360, new_R2278_U361, new_R2278_U362,
    new_R2278_U363, new_R2278_U364, new_R2278_U365, new_R2278_U366,
    new_R2278_U367, new_R2278_U368, new_R2278_U369, new_R2278_U370,
    new_R2278_U371, new_R2278_U372, new_R2278_U373, new_R2278_U374,
    new_R2278_U375, new_R2278_U376, new_R2278_U377, new_R2278_U378,
    new_R2278_U379, new_R2278_U380, new_R2278_U381, new_R2278_U382,
    new_R2278_U383, new_R2278_U384, new_R2278_U385, new_R2278_U386,
    new_R2278_U387, new_R2278_U388, new_R2278_U389, new_R2278_U390,
    new_R2278_U391, new_R2278_U392, new_R2278_U393, new_R2278_U394,
    new_R2278_U395, new_R2278_U396, new_R2278_U397, new_R2278_U398,
    new_R2278_U399, new_R2278_U400, new_R2278_U401, new_R2278_U402,
    new_R2278_U403, new_R2278_U404, new_R2278_U405, new_R2278_U406,
    new_R2278_U407, new_R2278_U408, new_R2278_U409, new_R2278_U410,
    new_R2278_U411, new_R2278_U412, new_R2278_U413, new_R2278_U414,
    new_R2278_U415, new_R2278_U416, new_R2278_U417, new_R2278_U418,
    new_R2278_U419, new_R2278_U420, new_R2278_U421, new_R2278_U422,
    new_R2358_U5, new_R2358_U6, new_R2358_U7, new_R2358_U8, new_R2358_U9,
    new_R2358_U10, new_R2358_U11, new_R2358_U12, new_R2358_U13,
    new_R2358_U14, new_R2358_U15, new_R2358_U16, new_R2358_U17,
    new_R2358_U18, new_R2358_U19, new_R2358_U20, new_R2358_U21,
    new_R2358_U22, new_R2358_U23, new_R2358_U24, new_R2358_U25,
    new_R2358_U26, new_R2358_U27, new_R2358_U28, new_R2358_U29,
    new_R2358_U30, new_R2358_U31, new_R2358_U32, new_R2358_U33,
    new_R2358_U34, new_R2358_U35, new_R2358_U36, new_R2358_U37,
    new_R2358_U38, new_R2358_U39, new_R2358_U40, new_R2358_U41,
    new_R2358_U42, new_R2358_U43, new_R2358_U44, new_R2358_U45,
    new_R2358_U46, new_R2358_U47, new_R2358_U48, new_R2358_U49,
    new_R2358_U50, new_R2358_U51, new_R2358_U52, new_R2358_U53,
    new_R2358_U54, new_R2358_U55, new_R2358_U56, new_R2358_U57,
    new_R2358_U58, new_R2358_U59, new_R2358_U60, new_R2358_U61,
    new_R2358_U62, new_R2358_U63, new_R2358_U64, new_R2358_U65,
    new_R2358_U66, new_R2358_U67, new_R2358_U68, new_R2358_U69,
    new_R2358_U70, new_R2358_U71, new_R2358_U72, new_R2358_U73,
    new_R2358_U74, new_R2358_U75, new_R2358_U76, new_R2358_U77,
    new_R2358_U78, new_R2358_U79, new_R2358_U80, new_R2358_U81,
    new_R2358_U82, new_R2358_U83, new_R2358_U84, new_R2358_U85,
    new_R2358_U86, new_R2358_U87, new_R2358_U88, new_R2358_U89,
    new_R2358_U90, new_R2358_U91, new_R2358_U92, new_R2358_U93,
    new_R2358_U94, new_R2358_U95, new_R2358_U96, new_R2358_U97,
    new_R2358_U98, new_R2358_U99, new_R2358_U100, new_R2358_U101,
    new_R2358_U102, new_R2358_U103, new_R2358_U104, new_R2358_U105,
    new_R2358_U106, new_R2358_U107, new_R2358_U108, new_R2358_U109,
    new_R2358_U110, new_R2358_U111, new_R2358_U112, new_R2358_U113,
    new_R2358_U114, new_R2358_U115, new_R2358_U116, new_R2358_U117,
    new_R2358_U118, new_R2358_U119, new_R2358_U120, new_R2358_U121,
    new_R2358_U122, new_R2358_U123, new_R2358_U124, new_R2358_U125,
    new_R2358_U126, new_R2358_U127, new_R2358_U128, new_R2358_U129,
    new_R2358_U130, new_R2358_U131, new_R2358_U132, new_R2358_U133,
    new_R2358_U134, new_R2358_U135, new_R2358_U136, new_R2358_U137,
    new_R2358_U138, new_R2358_U139, new_R2358_U140, new_R2358_U141,
    new_R2358_U142, new_R2358_U143, new_R2358_U144, new_R2358_U145,
    new_R2358_U146, new_R2358_U147, new_R2358_U148, new_R2358_U149,
    new_R2358_U150, new_R2358_U151, new_R2358_U152, new_R2358_U153,
    new_R2358_U154, new_R2358_U155, new_R2358_U156, new_R2358_U157,
    new_R2358_U158, new_R2358_U159, new_R2358_U160, new_R2358_U161,
    new_R2358_U162, new_R2358_U163, new_R2358_U164, new_R2358_U165,
    new_R2358_U166, new_R2358_U167, new_R2358_U168, new_R2358_U169,
    new_R2358_U170, new_R2358_U171, new_R2358_U172, new_R2358_U173,
    new_R2358_U174, new_R2358_U175, new_R2358_U176, new_R2358_U177,
    new_R2358_U178, new_R2358_U179, new_R2358_U180, new_R2358_U181,
    new_R2358_U182, new_R2358_U183, new_R2358_U184, new_R2358_U185,
    new_R2358_U186, new_R2358_U187, new_R2358_U188, new_R2358_U189,
    new_R2358_U190, new_R2358_U191, new_R2358_U192, new_R2358_U193,
    new_R2358_U194, new_R2358_U195, new_R2358_U196, new_R2358_U197,
    new_R2358_U198, new_R2358_U199, new_R2358_U200, new_R2358_U201,
    new_R2358_U202, new_R2358_U203, new_R2358_U204, new_R2358_U205,
    new_R2358_U206, new_R2358_U207, new_R2358_U208, new_R2358_U209,
    new_R2358_U210, new_R2358_U211, new_R2358_U212, new_R2358_U213,
    new_R2358_U214, new_R2358_U215, new_R2358_U216, new_R2358_U217,
    new_R2358_U218, new_R2358_U219, new_R2358_U220, new_R2358_U221,
    new_R2358_U222, new_R2358_U223, new_R2358_U224, new_R2358_U225,
    new_R2358_U226, new_R2358_U227, new_R2358_U228, new_R2358_U229,
    new_R2358_U230, new_R2358_U231, new_R2358_U232, new_R2358_U233,
    new_R2358_U234, new_R2358_U235, new_R2358_U236, new_R2358_U237,
    new_R2358_U238, new_R2358_U239, new_R2358_U240, new_R2358_U241,
    new_R2358_U242, new_R2358_U243, new_R2358_U244, new_R2358_U245,
    new_R2358_U246, new_R2358_U247, new_R2358_U248, new_R2358_U249,
    new_R2358_U250, new_R2358_U251, new_R2358_U252, new_R2358_U253,
    new_R2358_U254, new_R2358_U255, new_R2358_U256, new_R2358_U257,
    new_R2358_U258, new_R2358_U259, new_R2358_U260, new_R2358_U261,
    new_R2358_U262, new_R2358_U263, new_R2358_U264, new_R2358_U265,
    new_R2358_U266, new_R2358_U267, new_R2358_U268, new_R2358_U269,
    new_R2358_U270, new_R2358_U271, new_R2358_U272, new_R2358_U273,
    new_R2358_U274, new_R2358_U275, new_R2358_U276, new_R2358_U277,
    new_R2358_U278, new_R2358_U279, new_R2358_U280, new_R2358_U281,
    new_R2358_U282, new_R2358_U283, new_R2358_U284, new_R2358_U285,
    new_R2358_U286, new_R2358_U287, new_R2358_U288, new_R2358_U289,
    new_R2358_U290, new_R2358_U291, new_R2358_U292, new_R2358_U293,
    new_R2358_U294, new_R2358_U295, new_R2358_U296, new_R2358_U297,
    new_R2358_U298, new_R2358_U299, new_R2358_U300, new_R2358_U301,
    new_R2358_U302, new_R2358_U303, new_R2358_U304, new_R2358_U305,
    new_R2358_U306, new_R2358_U307, new_R2358_U308, new_R2358_U309,
    new_R2358_U310, new_R2358_U311, new_R2358_U312, new_R2358_U313,
    new_R2358_U314, new_R2358_U315, new_R2358_U316, new_R2358_U317,
    new_R2358_U318, new_R2358_U319, new_R2358_U320, new_R2358_U321,
    new_R2358_U322, new_R2358_U323, new_R2358_U324, new_R2358_U325,
    new_R2358_U326, new_R2358_U327, new_R2358_U328, new_R2358_U329,
    new_R2358_U330, new_R2358_U331, new_R2358_U332, new_R2358_U333,
    new_R2358_U334, new_R2358_U335, new_R2358_U336, new_R2358_U337,
    new_R2358_U338, new_R2358_U339, new_R2358_U340, new_R2358_U341,
    new_R2358_U342, new_R2358_U343, new_R2358_U344, new_R2358_U345,
    new_R2358_U346, new_R2358_U347, new_R2358_U348, new_R2358_U349,
    new_R2358_U350, new_R2358_U351, new_R2358_U352, new_R2358_U353,
    new_R2358_U354, new_R2358_U355, new_R2358_U356, new_R2358_U357,
    new_R2358_U358, new_R2358_U359, new_R2358_U360, new_R2358_U361,
    new_R2358_U362, new_R2358_U363, new_R2358_U364, new_R2358_U365,
    new_R2358_U366, new_R2358_U367, new_R2358_U368, new_R2358_U369,
    new_R2358_U370, new_R2358_U371, new_R2358_U372, new_R2358_U373,
    new_R2358_U374, new_R2358_U375, new_R2358_U376, new_R2358_U377,
    new_R2358_U378, new_R2358_U379, new_R2358_U380, new_R2358_U381,
    new_R2358_U382, new_R2358_U383, new_R2358_U384, new_R2358_U385,
    new_R2358_U386, new_R2358_U387, new_R2358_U388, new_R2358_U389,
    new_R2358_U390, new_R2358_U391, new_R2358_U392, new_R2358_U393,
    new_R2358_U394, new_R2358_U395, new_R2358_U396, new_R2358_U397,
    new_R2358_U398, new_R2358_U399, new_R2358_U400, new_R2358_U401,
    new_R2358_U402, new_R2358_U403, new_R2358_U404, new_R2358_U405,
    new_R2358_U406, new_R2358_U407, new_R2358_U408, new_R2358_U409,
    new_R2358_U410, new_R2358_U411, new_R2358_U412, new_R2358_U413,
    new_R2358_U414, new_R2358_U415, new_R2358_U416, new_R2358_U417,
    new_R2358_U418, new_R2358_U419, new_R2358_U420, new_R2358_U421,
    new_R2358_U422, new_R2358_U423, new_R2358_U424, new_R2358_U425,
    new_R2358_U426, new_R2358_U427, new_R2358_U428, new_R2358_U429,
    new_R2358_U430, new_R2358_U431, new_R2358_U432, new_R2358_U433,
    new_R2358_U434, new_R2358_U435, new_R2358_U436, new_R2358_U437,
    new_R2358_U438, new_R2358_U439, new_R2358_U440, new_R2358_U441,
    new_R2358_U442, new_R2358_U443, new_R2358_U444, new_R2358_U445,
    new_R2358_U446, new_R2358_U447, new_R2358_U448, new_R2358_U449,
    new_R2358_U450, new_R2358_U451, new_R2358_U452, new_R2358_U453,
    new_R2358_U454, new_R2358_U455, new_R2358_U456, new_R2358_U457,
    new_R2358_U458, new_R2358_U459, new_R2358_U460, new_R2358_U461,
    new_R2358_U462, new_R2358_U463, new_R2358_U464, new_R2358_U465,
    new_R2358_U466, new_R2358_U467, new_R2358_U468, new_R2358_U469,
    new_R2358_U470, new_R2358_U471, new_R2358_U472, new_R2358_U473,
    new_R2358_U474, new_R2358_U475, new_R2358_U476, new_R2358_U477,
    new_R2358_U478, new_R2358_U479, new_R2358_U480, new_R2358_U481,
    new_R2358_U482, new_R2358_U483, new_R2358_U484, new_R2358_U485,
    new_R2358_U486, new_R2358_U487, new_R2358_U488, new_R2358_U489,
    new_R2358_U490, new_R2358_U491, new_R2358_U492, new_R2358_U493,
    new_R2358_U494, new_R2358_U495, new_R2358_U496, new_R2358_U497,
    new_R2358_U498, new_R2358_U499, new_R2358_U500, new_R2358_U501,
    new_R2358_U502, new_R2358_U503, new_R2358_U504, new_R2358_U505,
    new_R2358_U506, new_R2358_U507, new_R2358_U508, new_R2358_U509,
    new_R2358_U510, new_R2358_U511, new_R2358_U512, new_R2358_U513,
    new_R2358_U514, new_R2358_U515, new_R2358_U516, new_R2358_U517,
    new_R2358_U518, new_R2358_U519, new_R2358_U520, new_R2358_U521,
    new_R2358_U522, new_R2358_U523, new_R2358_U524, new_R2358_U525,
    new_R2358_U526, new_R2358_U527, new_R2358_U528, new_R2358_U529,
    new_R2358_U530, new_R2358_U531, new_R2358_U532, new_R2358_U533,
    new_R2358_U534, new_R2358_U535, new_R2358_U536, new_R2358_U537,
    new_R2358_U538, new_R2358_U539, new_R2358_U540, new_R2358_U541,
    new_R2358_U542, new_R2358_U543, new_R2358_U544, new_R2358_U545,
    new_R2358_U546, new_R2358_U547, new_R2358_U548, new_R2358_U549,
    new_R2358_U550, new_R2358_U551, new_R2358_U552, new_R2358_U553,
    new_R2358_U554, new_R2358_U555, new_R2358_U556, new_R2358_U557,
    new_R2358_U558, new_R2358_U559, new_R2358_U560, new_R2358_U561,
    new_R2358_U562, new_R2358_U563, new_R2358_U564, new_R2358_U565,
    new_R2358_U566, new_R2358_U567, new_R2358_U568, new_R2358_U569,
    new_R2358_U570, new_R2358_U571, new_R2358_U572, new_R2358_U573,
    new_R2358_U574, new_R2358_U575, new_R2358_U576, new_R2358_U577,
    new_R2358_U578, new_R2358_U579, new_R2358_U580, new_R2358_U581,
    new_R2358_U582, new_R2358_U583, new_R2358_U584, new_R2358_U585,
    new_R2358_U586, new_R2358_U587, new_R2358_U588, new_R2358_U589,
    new_R2358_U590, new_R2358_U591, new_R2358_U592, new_R2358_U593,
    new_R2358_U594, new_R2358_U595, new_R2358_U596, new_R2358_U597,
    new_R2358_U598, new_R2358_U599, new_R2358_U600, new_R2358_U601,
    new_R2358_U602, new_R2358_U603, new_R2358_U604, new_R2358_U605,
    new_R2358_U606, new_R2358_U607, new_R2358_U608, new_R2358_U609,
    new_R2358_U610, new_R2358_U611, new_R2358_U612, new_R2358_U613,
    new_R2358_U614, new_R2358_U615, new_R2358_U616, new_R2358_U617,
    new_R2358_U618, new_R2358_U619, new_R2358_U620, new_R2358_U621,
    new_R2358_U622, new_R2358_U623, new_R2358_U624, new_R2358_U625,
    new_R2358_U626, new_R2358_U627, new_R2358_U628, new_R2358_U629,
    new_R2358_U630, new_R2358_U631, new_R2358_U632, new_R2358_U633,
    new_R2358_U634, new_R2358_U635, new_R2358_U636, new_R2358_U637,
    new_R2358_U638, new_R2358_U639, new_R2358_U640, new_R2358_U641,
    new_R2358_U642, new_R2358_U643, new_R2358_U644, new_R2358_U645,
    new_R2358_U646, new_R2358_U647, new_R2358_U648, new_R2358_U649,
    new_R2358_U650, new_R2358_U651, new_R2358_U652, new_R2358_U653,
    new_R2358_U654, new_R2337_U5, new_R2337_U6, new_R2337_U7, new_R2337_U8,
    new_R2337_U9, new_R2337_U10, new_R2337_U11, new_R2337_U12,
    new_R2337_U13, new_R2337_U14, new_R2337_U15, new_R2337_U16,
    new_R2337_U17, new_R2337_U18, new_R2337_U19, new_R2337_U20,
    new_R2337_U21, new_R2337_U22, new_R2337_U23, new_R2337_U24,
    new_R2337_U25, new_R2337_U26, new_R2337_U27, new_R2337_U28,
    new_R2337_U29, new_R2337_U30, new_R2337_U31, new_R2337_U32,
    new_R2337_U33, new_R2337_U34, new_R2337_U35, new_R2337_U36,
    new_R2337_U37, new_R2337_U38, new_R2337_U39, new_R2337_U40,
    new_R2337_U41, new_R2337_U42, new_R2337_U43, new_R2337_U44,
    new_R2337_U45, new_R2337_U46, new_R2337_U47, new_R2337_U48,
    new_R2337_U49, new_R2337_U50, new_R2337_U51, new_R2337_U52,
    new_R2337_U53, new_R2337_U54, new_R2337_U55, new_R2337_U56,
    new_R2337_U57, new_R2337_U58, new_R2337_U59, new_R2337_U60,
    new_R2337_U61, new_R2337_U62, new_R2337_U63, new_R2337_U64,
    new_R2337_U65, new_R2337_U66, new_R2337_U67, new_R2337_U68,
    new_R2337_U69, new_R2337_U70, new_R2337_U71, new_R2337_U72,
    new_R2337_U73, new_R2337_U74, new_R2337_U75, new_R2337_U76,
    new_R2337_U77, new_R2337_U78, new_R2337_U79, new_R2337_U80,
    new_R2337_U81, new_R2337_U82, new_R2337_U83, new_R2337_U84,
    new_R2337_U85, new_R2337_U86, new_R2337_U87, new_R2337_U88,
    new_R2337_U89, new_R2337_U90, new_R2337_U91, new_R2337_U92,
    new_R2337_U93, new_R2337_U94, new_R2337_U95, new_R2337_U96,
    new_R2337_U97, new_R2337_U98, new_R2337_U99, new_R2337_U100,
    new_R2337_U101, new_R2337_U102, new_R2337_U103, new_R2337_U104,
    new_R2337_U105, new_R2337_U106, new_R2337_U107, new_R2337_U108,
    new_R2337_U109, new_R2337_U110, new_R2337_U111, new_R2337_U112,
    new_R2337_U113, new_R2337_U114, new_R2337_U115, new_R2337_U116,
    new_R2337_U117, new_R2337_U118, new_R2337_U119, new_R2337_U120,
    new_R2337_U121, new_R2337_U122, new_R2337_U123, new_R2337_U124,
    new_R2337_U125, new_R2337_U126, new_R2337_U127, new_R2337_U128,
    new_R2337_U129, new_R2337_U130, new_R2337_U131, new_R2337_U132,
    new_R2337_U133, new_R2337_U134, new_R2337_U135, new_R2337_U136,
    new_R2337_U137, new_R2337_U138, new_R2337_U139, new_R2337_U140,
    new_R2337_U141, new_R2337_U142, new_R2337_U143, new_R2337_U144,
    new_R2337_U145, new_R2337_U146, new_R2337_U147, new_R2337_U148,
    new_R2337_U149, new_R2337_U150, new_R2337_U151, new_R2337_U152,
    new_R2337_U153, new_R2337_U154, new_R2337_U155, new_R2337_U156,
    new_R2337_U157, new_R2337_U158, new_R2337_U159, new_R2337_U160,
    new_R2337_U161, new_R2337_U162, new_R2337_U163, new_R2337_U164,
    new_R2337_U165, new_R2337_U166, new_R2337_U167, new_R2337_U168,
    new_R2337_U169, new_R2337_U170, new_R2337_U171, new_R2337_U172,
    new_R2337_U173, new_R2337_U174, new_R2337_U175, new_R2337_U176,
    new_R2337_U177, new_R2337_U178, new_R2337_U179, new_R2337_U180,
    new_R2337_U181, new_R2337_U182, new_R2337_U183, new_R2337_U184,
    new_R2337_U185, new_R2337_U186, new_R2337_U187, new_R2337_U188,
    new_R2337_U189, new_R2337_U190, new_R2337_U191, new_R2337_U192,
    new_R2337_U193, new_R2182_U5, new_R2182_U6, new_R2182_U7, new_R2182_U8,
    new_R2182_U9, new_R2182_U10, new_R2182_U11, new_R2182_U12,
    new_R2182_U13, new_R2182_U14, new_R2182_U15, new_R2182_U16,
    new_R2182_U17, new_R2182_U18, new_R2182_U19, new_R2182_U20,
    new_R2182_U21, new_R2182_U22, new_R2182_U23, new_R2182_U24,
    new_R2182_U25, new_R2182_U26, new_R2182_U27, new_R2182_U28,
    new_R2182_U29, new_R2182_U30, new_R2182_U31, new_R2182_U32,
    new_R2182_U33, new_R2182_U34, new_R2182_U35, new_R2182_U36,
    new_R2182_U37, new_R2182_U38, new_R2182_U39, new_R2182_U40,
    new_R2182_U41, new_R2182_U42, new_R2182_U43, new_R2182_U44,
    new_R2182_U45, new_R2182_U46, new_R2182_U47, new_R2182_U48,
    new_R2182_U49, new_R2182_U50, new_R2182_U51, new_R2182_U52,
    new_R2182_U53, new_R2182_U54, new_R2182_U55, new_R2182_U56,
    new_R2182_U57, new_R2182_U58, new_R2182_U59, new_R2182_U60,
    new_R2182_U61, new_R2182_U62, new_R2182_U63, new_R2182_U64,
    new_R2182_U65, new_R2182_U66, new_R2182_U67, new_R2182_U68,
    new_R2182_U69, new_R2182_U70, new_R2182_U71, new_R2182_U72,
    new_R2182_U73, new_R2182_U74, new_R2182_U75, new_R2182_U76,
    new_R2182_U77, new_R2182_U78, new_R2182_U79, new_R2182_U80,
    new_R2182_U81, new_R2182_U82, new_R2182_U83, new_R2182_U84,
    new_R2182_U85, new_R2182_U86, new_R2144_U5, new_R2144_U6, new_R2144_U7,
    new_R2144_U8, new_R2144_U9, new_R2144_U10, new_R2144_U11,
    new_R2144_U12, new_R2144_U13, new_R2144_U14, new_R2144_U15,
    new_R2144_U16, new_R2144_U17, new_R2144_U18, new_R2144_U19,
    new_R2144_U20, new_R2144_U21, new_R2144_U22, new_R2144_U23,
    new_R2144_U24, new_R2144_U25, new_R2144_U26, new_R2144_U27,
    new_R2144_U28, new_R2144_U29, new_R2144_U30, new_R2144_U31,
    new_R2144_U32, new_R2144_U33, new_R2144_U34, new_R2144_U35,
    new_R2144_U36, new_R2144_U37, new_R2144_U38, new_R2144_U39,
    new_R2144_U40, new_R2144_U41, new_R2144_U42, new_R2144_U43,
    new_R2144_U44, new_R2144_U45, new_R2144_U46, new_R2144_U47,
    new_R2144_U48, new_R2144_U49, new_R2144_U50, new_R2144_U51,
    new_R2144_U52, new_R2144_U53, new_R2144_U54, new_R2144_U55,
    new_R2144_U56, new_R2144_U57, new_R2144_U58, new_R2144_U59,
    new_R2144_U60, new_R2144_U61, new_R2144_U62, new_R2144_U63,
    new_R2144_U64, new_R2144_U65, new_R2144_U66, new_R2144_U67,
    new_R2144_U68, new_R2144_U69, new_R2144_U70, new_R2144_U71,
    new_R2144_U72, new_R2144_U73, new_R2144_U74, new_R2144_U75,
    new_R2144_U76, new_R2144_U77, new_R2144_U78, new_R2144_U79,
    new_R2144_U80, new_R2144_U81, new_R2144_U82, new_R2144_U83,
    new_R2144_U84, new_R2144_U85, new_R2144_U86, new_R2144_U87,
    new_R2144_U88, new_R2144_U89, new_R2144_U90, new_R2144_U91,
    new_R2144_U92, new_R2144_U93, new_R2144_U94, new_R2144_U95,
    new_R2144_U96, new_R2144_U97, new_R2144_U98, new_R2144_U99,
    new_R2144_U100, new_R2144_U101, new_R2144_U102, new_R2144_U103,
    new_R2144_U104, new_R2144_U105, new_R2144_U106, new_R2144_U107,
    new_R2144_U108, new_R2144_U109, new_R2144_U110, new_R2144_U111,
    new_R2144_U112, new_R2144_U113, new_R2144_U114, new_R2144_U115,
    new_R2144_U116, new_R2144_U117, new_R2144_U118, new_R2144_U119,
    new_R2144_U120, new_R2144_U121, new_R2144_U122, new_R2144_U123,
    new_R2144_U124, new_R2144_U125, new_R2144_U126, new_R2144_U127,
    new_R2144_U128, new_R2144_U129, new_R2144_U130, new_R2144_U131,
    new_R2144_U132, new_R2144_U133, new_R2144_U134, new_R2144_U135,
    new_R2144_U136, new_R2144_U137, new_R2144_U138, new_R2144_U139,
    new_R2144_U140, new_R2144_U141, new_R2144_U142, new_R2144_U143,
    new_R2144_U144, new_R2144_U145, new_R2144_U146, new_R2144_U147,
    new_R2144_U148, new_R2144_U149, new_R2144_U150, new_R2144_U151,
    new_R2144_U152, new_R2144_U153, new_R2144_U154, new_R2144_U155,
    new_R2144_U156, new_R2144_U157, new_R2144_U158, new_R2144_U159,
    new_R2144_U160, new_R2144_U161, new_R2144_U162, new_R2144_U163,
    new_R2144_U164, new_R2144_U165, new_R2144_U166, new_R2144_U167,
    new_R2144_U168, new_R2144_U169, new_R2144_U170, new_R2144_U171,
    new_R2144_U172, new_R2144_U173, new_R2144_U174, new_R2144_U175,
    new_R2144_U176, new_R2144_U177, new_R2144_U178, new_R2144_U179,
    new_R2144_U180, new_R2144_U181, new_R2144_U182, new_R2144_U183,
    new_R2144_U184, new_R2144_U185, new_R2144_U186, new_R2144_U187,
    new_R2144_U188, new_R2144_U189, new_R2144_U190, new_R2144_U191,
    new_R2144_U192, new_R2144_U193, new_R2144_U194, new_R2144_U195,
    new_R2144_U196, new_R2144_U197, new_R2144_U198, new_R2144_U199,
    new_R2144_U200, new_R2144_U201, new_R2144_U202, new_R2144_U203,
    new_R2144_U204, new_R2144_U205, new_R2144_U206, new_R2144_U207,
    new_R2144_U208, new_R2144_U209, new_R2144_U210, new_R2144_U211,
    new_R2144_U212, new_R2144_U213, new_R2144_U214, new_R2144_U215,
    new_R2144_U216, new_R2144_U217, new_R2144_U218, new_R2144_U219,
    new_R2144_U220, new_R2144_U221, new_R2144_U222, new_R2144_U223,
    new_R2144_U224, new_R2144_U225, new_R2144_U226, new_R2144_U227,
    new_R2144_U228, new_R2144_U229, new_R2144_U230, new_R2144_U231,
    new_R2144_U232, new_R2144_U233, new_R2144_U234, new_R2144_U235,
    new_R2144_U236, new_R2144_U237, new_R2144_U238, new_R2144_U239,
    new_R2144_U240, new_R2144_U241, new_R2144_U242, new_R2144_U243,
    new_R2144_U244, new_R2144_U245, new_R2144_U246, new_R2144_U247,
    new_R2144_U248, new_R2144_U249, new_R2144_U250, new_R2144_U251,
    new_R2144_U252, new_R2144_U253, new_R2144_U254, new_R2144_U255,
    new_R2144_U256, new_R2144_U257, new_R2144_U258, new_R2144_U259,
    new_R2144_U260, new_LT_589_U6, new_LT_589_U7, new_LT_589_U8,
    new_R584_U6, new_R584_U7, new_R584_U8, new_R584_U9, new_R2099_U4,
    new_R2099_U5, new_R2099_U6, new_R2099_U7, new_R2099_U8, new_R2099_U9,
    new_R2099_U10, new_R2099_U11, new_R2099_U12, new_R2099_U13,
    new_R2099_U14, new_R2099_U15, new_R2099_U16, new_R2099_U17,
    new_R2099_U18, new_R2099_U19, new_R2099_U20, new_R2099_U21,
    new_R2099_U22, new_R2099_U23, new_R2099_U24, new_R2099_U25,
    new_R2099_U26, new_R2099_U27, new_R2099_U28, new_R2099_U29,
    new_R2099_U30, new_R2099_U31, new_R2099_U32, new_R2099_U33,
    new_R2099_U34, new_R2099_U35, new_R2099_U36, new_R2099_U37,
    new_R2099_U38, new_R2099_U39, new_R2099_U40, new_R2099_U41,
    new_R2099_U42, new_R2099_U43, new_R2099_U44, new_R2099_U45,
    new_R2099_U46, new_R2099_U47, new_R2099_U48, new_R2099_U49,
    new_R2099_U50, new_R2099_U51, new_R2099_U52, new_R2099_U53,
    new_R2099_U54, new_R2099_U55, new_R2099_U56, new_R2099_U57,
    new_R2099_U58, new_R2099_U59, new_R2099_U60, new_R2099_U61,
    new_R2099_U62, new_R2099_U63, new_R2099_U64, new_R2099_U65,
    new_R2099_U66, new_R2099_U67, new_R2099_U68, new_R2099_U69,
    new_R2099_U70, new_R2099_U71, new_R2099_U72, new_R2099_U73,
    new_R2099_U74, new_R2099_U75, new_R2099_U76, new_R2099_U77,
    new_R2099_U78, new_R2099_U79, new_R2099_U80, new_R2099_U81,
    new_R2099_U82, new_R2099_U83, new_R2099_U84, new_R2099_U85,
    new_R2099_U86, new_R2099_U87, new_R2099_U88, new_R2099_U89,
    new_R2099_U90, new_R2099_U91, new_R2099_U92, new_R2099_U93,
    new_R2099_U94, new_R2099_U95, new_R2099_U96, new_R2099_U97,
    new_R2099_U98, new_R2099_U99, new_R2099_U100, new_R2099_U101,
    new_R2099_U102, new_R2099_U103, new_R2099_U104, new_R2099_U105,
    new_R2099_U106, new_R2099_U107, new_R2099_U108, new_R2099_U109,
    new_R2099_U110, new_R2099_U111, new_R2099_U112, new_R2099_U113,
    new_R2099_U114, new_R2099_U115, new_R2099_U116, new_R2099_U117,
    new_R2099_U118, new_R2099_U119, new_R2099_U120, new_R2099_U121,
    new_R2099_U122, new_R2099_U123, new_R2099_U124, new_R2099_U125,
    new_R2099_U126, new_R2099_U127, new_R2099_U128, new_R2099_U129,
    new_R2099_U130, new_R2099_U131, new_R2099_U132, new_R2099_U133,
    new_R2099_U134, new_R2099_U135, new_R2099_U136, new_R2099_U137,
    new_R2099_U138, new_R2099_U139, new_R2099_U140, new_R2099_U141,
    new_R2099_U142, new_R2099_U143, new_R2099_U144, new_R2099_U145,
    new_R2099_U146, new_R2099_U147, new_R2099_U148, new_R2099_U149,
    new_R2099_U150, new_R2099_U151, new_R2099_U152, new_R2099_U153,
    new_R2099_U154, new_R2099_U155, new_R2099_U156, new_R2099_U157,
    new_R2099_U158, new_R2099_U159, new_R2099_U160, new_R2099_U161,
    new_R2099_U162, new_R2099_U163, new_R2099_U164, new_R2099_U165,
    new_R2099_U166, new_R2099_U167, new_R2099_U168, new_R2099_U169,
    new_R2099_U170, new_R2099_U171, new_R2099_U172, new_R2099_U173,
    new_R2099_U174, new_R2099_U175, new_R2099_U176, new_R2099_U177,
    new_R2099_U178, new_R2099_U179, new_R2099_U180, new_R2099_U181,
    new_R2099_U182, new_R2099_U183, new_R2099_U184, new_R2099_U185,
    new_R2099_U186, new_R2099_U187, new_R2099_U188, new_R2099_U189,
    new_R2099_U190, new_R2099_U191, new_R2099_U192, new_R2099_U193,
    new_R2099_U194, new_R2099_U195, new_R2099_U196, new_R2099_U197,
    new_R2099_U198, new_R2099_U199, new_R2099_U200, new_R2099_U201,
    new_R2099_U202, new_R2099_U203, new_R2099_U204, new_R2099_U205,
    new_R2099_U206, new_R2099_U207, new_R2099_U208, new_R2099_U209,
    new_R2099_U210, new_R2099_U211, new_R2099_U212, new_R2099_U213,
    new_R2099_U214, new_R2099_U215, new_R2099_U216, new_R2099_U217,
    new_R2099_U218, new_R2099_U219, new_R2099_U220, new_R2099_U221,
    new_R2099_U222, new_R2099_U223, new_R2099_U224, new_R2099_U225,
    new_R2099_U226, new_R2099_U227, new_R2099_U228, new_R2099_U229,
    new_R2099_U230, new_R2099_U231, new_R2099_U232, new_R2099_U233,
    new_R2099_U234, new_R2099_U235, new_R2099_U236, new_R2099_U237,
    new_R2099_U238, new_R2099_U239, new_R2099_U240, new_R2099_U241,
    new_R2099_U242, new_R2099_U243, new_R2099_U244, new_R2099_U245,
    new_R2099_U246, new_R2099_U247, new_R2099_U248, new_R2099_U249,
    new_R2099_U250, new_R2099_U251, new_R2099_U252, new_R2099_U253,
    new_R2099_U254, new_R2099_U255, new_R2099_U256, new_R2099_U257,
    new_R2099_U258, new_R2099_U259, new_R2099_U260, new_R2099_U261,
    new_R2099_U262, new_R2099_U263, new_R2099_U264, new_R2099_U265,
    new_R2099_U266, new_R2099_U267, new_R2099_U268, new_R2099_U269,
    new_R2099_U270, new_R2099_U271, new_R2099_U272, new_R2099_U273,
    new_R2099_U274, new_R2099_U275, new_R2099_U276, new_R2099_U277,
    new_R2099_U278, new_R2099_U279, new_R2099_U280, new_R2099_U281,
    new_R2099_U282, new_R2099_U283, new_R2099_U284, new_R2099_U285,
    new_R2099_U286, new_R2099_U287, new_R2099_U288, new_R2099_U289,
    new_R2099_U290, new_R2099_U291, new_R2099_U292, new_R2099_U293,
    new_R2099_U294, new_R2099_U295, new_R2099_U296, new_R2099_U297,
    new_R2099_U298, new_R2099_U299, new_R2099_U300, new_R2099_U301,
    new_R2099_U302, new_R2099_U303, new_R2099_U304, new_R2099_U305,
    new_R2099_U306, new_R2099_U307, new_R2099_U308, new_R2099_U309,
    new_R2099_U310, new_R2099_U311, new_R2099_U312, new_R2099_U313,
    new_R2099_U314, new_R2099_U315, new_R2099_U316, new_R2099_U317,
    new_R2099_U318, new_R2099_U319, new_R2099_U320, new_R2099_U321,
    new_R2099_U322, new_R2099_U323, new_R2099_U324, new_R2099_U325,
    new_R2099_U326, new_R2099_U327, new_R2099_U328, new_R2099_U329,
    new_R2099_U330, new_R2099_U331, new_R2099_U332, new_R2099_U333,
    new_R2099_U334, new_R2099_U335, new_R2099_U336, new_R2099_U337,
    new_R2099_U338, new_R2099_U339, new_R2099_U340, new_R2099_U341,
    new_R2099_U342, new_R2099_U343, new_R2099_U344, new_R2099_U345,
    new_R2099_U346, new_R2099_U347, new_R2099_U348, new_R2099_U349,
    new_R2167_U6, new_R2167_U7, new_R2167_U8, new_R2167_U9, new_R2167_U10,
    new_R2167_U11, new_R2167_U12, new_R2167_U13, new_R2167_U14,
    new_R2167_U15, new_R2167_U16, new_R2167_U17, new_R2167_U18,
    new_R2167_U19, new_R2167_U20, new_R2167_U21, new_R2167_U22,
    new_R2167_U23, new_R2167_U24, new_R2167_U25, new_R2167_U26,
    new_R2167_U27, new_R2167_U28, new_R2167_U29, new_R2167_U30,
    new_R2167_U31, new_R2167_U32, new_R2167_U33, new_R2167_U34,
    new_R2167_U35, new_R2167_U36, new_R2167_U37, new_R2167_U38,
    new_R2167_U39, new_R2167_U40, new_R2167_U41, new_R2167_U42,
    new_R2167_U43, new_R2167_U44, new_R2167_U45, new_R2167_U46,
    new_R2167_U47, new_R2167_U48, new_R2167_U49, new_R2167_U50,
    new_SUB_357_U6, new_SUB_357_U7, new_SUB_357_U8, new_SUB_357_U9,
    new_SUB_357_U10, new_SUB_357_U11, new_SUB_357_U12, new_SUB_357_U13,
    new_LT_563_1260_U6, new_LT_563_1260_U7, new_LT_563_1260_U8,
    new_LT_563_1260_U9, new_SUB_580_U6, new_SUB_580_U7, new_SUB_580_U8,
    new_SUB_580_U9, new_SUB_580_U10, new_R2096_U4, new_R2096_U5,
    new_R2096_U6, new_R2096_U7, new_R2096_U8, new_R2096_U9, new_R2096_U10,
    new_R2096_U11, new_R2096_U12, new_R2096_U13, new_R2096_U14,
    new_R2096_U15, new_R2096_U16, new_R2096_U17, new_R2096_U18,
    new_R2096_U19, new_R2096_U20, new_R2096_U21, new_R2096_U22,
    new_R2096_U23, new_R2096_U24, new_R2096_U25, new_R2096_U26,
    new_R2096_U27, new_R2096_U28, new_R2096_U29, new_R2096_U30,
    new_R2096_U31, new_R2096_U32, new_R2096_U33, new_R2096_U34,
    new_R2096_U35, new_R2096_U36, new_R2096_U37, new_R2096_U38,
    new_R2096_U39, new_R2096_U40, new_R2096_U41, new_R2096_U42,
    new_R2096_U43, new_R2096_U44, new_R2096_U45, new_R2096_U46,
    new_R2096_U47, new_R2096_U48, new_R2096_U49, new_R2096_U50,
    new_R2096_U51, new_R2096_U52, new_R2096_U53, new_R2096_U54,
    new_R2096_U55, new_R2096_U56, new_R2096_U57, new_R2096_U58,
    new_R2096_U59, new_R2096_U60, new_R2096_U61, new_R2096_U62,
    new_R2096_U63, new_R2096_U64, new_R2096_U65, new_R2096_U66,
    new_R2096_U67, new_R2096_U68, new_R2096_U69, new_R2096_U70,
    new_R2096_U71, new_R2096_U72, new_R2096_U73, new_R2096_U74,
    new_R2096_U75, new_R2096_U76, new_R2096_U77, new_R2096_U78,
    new_R2096_U79, new_R2096_U80, new_R2096_U81, new_R2096_U82,
    new_R2096_U83, new_R2096_U84, new_R2096_U85, new_R2096_U86,
    new_R2096_U87, new_R2096_U88, new_R2096_U89, new_R2096_U90,
    new_R2096_U91, new_R2096_U92, new_R2096_U93, new_R2096_U94,
    new_R2096_U95, new_R2096_U96, new_R2096_U97, new_R2096_U98,
    new_R2096_U99, new_R2096_U100, new_R2096_U101, new_R2096_U102,
    new_R2096_U103, new_R2096_U104, new_R2096_U105, new_R2096_U106,
    new_R2096_U107, new_R2096_U108, new_R2096_U109, new_R2096_U110,
    new_R2096_U111, new_R2096_U112, new_R2096_U113, new_R2096_U114,
    new_R2096_U115, new_R2096_U116, new_R2096_U117, new_R2096_U118,
    new_R2096_U119, new_R2096_U120, new_R2096_U121, new_R2096_U122,
    new_R2096_U123, new_R2096_U124, new_R2096_U125, new_R2096_U126,
    new_R2096_U127, new_R2096_U128, new_R2096_U129, new_R2096_U130,
    new_R2096_U131, new_R2096_U132, new_R2096_U133, new_R2096_U134,
    new_R2096_U135, new_R2096_U136, new_R2096_U137, new_R2096_U138,
    new_R2096_U139, new_R2096_U140, new_R2096_U141, new_R2096_U142,
    new_R2096_U143, new_R2096_U144, new_R2096_U145, new_R2096_U146,
    new_R2096_U147, new_R2096_U148, new_R2096_U149, new_R2096_U150,
    new_R2096_U151, new_R2096_U152, new_R2096_U153, new_R2096_U154,
    new_R2096_U155, new_R2096_U156, new_R2096_U157, new_R2096_U158,
    new_R2096_U159, new_R2096_U160, new_R2096_U161, new_R2096_U162,
    new_R2096_U163, new_R2096_U164, new_R2096_U165, new_R2096_U166,
    new_R2096_U167, new_R2096_U168, new_R2096_U169, new_R2096_U170,
    new_R2096_U171, new_R2096_U172, new_R2096_U173, new_R2096_U174,
    new_R2096_U175, new_R2096_U176, new_R2096_U177, new_R2096_U178,
    new_R2096_U179, new_R2096_U180, new_R2096_U181, new_R2096_U182,
    new_LT_563_U6, new_LT_563_U7, new_LT_563_U8, new_LT_563_U9,
    new_LT_563_U10, new_LT_563_U11, new_LT_563_U12, new_LT_563_U13,
    new_LT_563_U14, new_LT_563_U15, new_LT_563_U16, new_LT_563_U17,
    new_LT_563_U18, new_LT_563_U19, new_LT_563_U20, new_LT_563_U21,
    new_LT_563_U22, new_LT_563_U23, new_LT_563_U24, new_LT_563_U25,
    new_LT_563_U26, new_LT_563_U27, new_LT_563_U28, new_R2238_U6,
    new_R2238_U7, new_R2238_U8, new_R2238_U9, new_R2238_U10, new_R2238_U11,
    new_R2238_U12, new_R2238_U13, new_R2238_U14, new_R2238_U15,
    new_R2238_U16, new_R2238_U17, new_R2238_U18, new_R2238_U19,
    new_R2238_U20, new_R2238_U21, new_R2238_U22, new_R2238_U23,
    new_R2238_U24, new_R2238_U25, new_R2238_U26, new_R2238_U27,
    new_R2238_U28, new_R2238_U29, new_R2238_U30, new_R2238_U31,
    new_R2238_U32, new_R2238_U33, new_R2238_U34, new_R2238_U35,
    new_R2238_U36, new_R2238_U37, new_R2238_U38, new_R2238_U39,
    new_R2238_U40, new_R2238_U41, new_R2238_U42, new_R2238_U43,
    new_R2238_U44, new_R2238_U45, new_R2238_U46, new_R2238_U47,
    new_R2238_U48, new_R2238_U49, new_R2238_U50, new_R2238_U51,
    new_R2238_U52, new_R2238_U53, new_R2238_U54, new_R2238_U55,
    new_R2238_U56, new_R2238_U57, new_R2238_U58, new_R2238_U59,
    new_R2238_U60, new_R2238_U61, new_R2238_U62, new_R2238_U63,
    new_R2238_U64, new_R2238_U65, new_R2238_U66, new_SUB_450_U6,
    new_SUB_450_U7, new_SUB_450_U8, new_SUB_450_U9, new_SUB_450_U10,
    new_SUB_450_U11, new_SUB_450_U12, new_SUB_450_U13, new_SUB_450_U14,
    new_SUB_450_U15, new_SUB_450_U16, new_SUB_450_U17, new_SUB_450_U18,
    new_SUB_450_U19, new_SUB_450_U20, new_SUB_450_U21, new_SUB_450_U22,
    new_SUB_450_U23, new_SUB_450_U24, new_SUB_450_U25, new_SUB_450_U26,
    new_SUB_450_U27, new_SUB_450_U28, new_SUB_450_U29, new_SUB_450_U30,
    new_SUB_450_U31, new_SUB_450_U32, new_SUB_450_U33, new_SUB_450_U34,
    new_SUB_450_U35, new_SUB_450_U36, new_SUB_450_U37, new_SUB_450_U38,
    new_SUB_450_U39, new_SUB_450_U40, new_SUB_450_U41, new_SUB_450_U42,
    new_SUB_450_U43, new_SUB_450_U44, new_SUB_450_U45, new_SUB_450_U46,
    new_SUB_450_U47, new_SUB_450_U48, new_SUB_450_U49, new_SUB_450_U50,
    new_SUB_450_U51, new_SUB_450_U52, new_SUB_450_U53, new_SUB_450_U54,
    new_SUB_450_U55, new_SUB_450_U56, new_SUB_450_U57, new_SUB_450_U58,
    new_SUB_450_U59, new_SUB_450_U60, new_SUB_450_U61, new_SUB_450_U62,
    new_SUB_450_U63, new_SUB_450_U64, new_SUB_450_U65, new_SUB_450_U66,
    new_ADD_371_U4, new_ADD_371_U5, new_ADD_371_U6, new_ADD_371_U7,
    new_ADD_371_U8, new_ADD_371_U9, new_ADD_371_U10, new_ADD_371_U11,
    new_ADD_371_U12, new_ADD_371_U13, new_ADD_371_U14, new_ADD_371_U15,
    new_ADD_371_U16, new_ADD_371_U17, new_ADD_371_U18, new_ADD_371_U19,
    new_ADD_371_U20, new_ADD_371_U21, new_ADD_371_U22, new_ADD_371_U23,
    new_ADD_371_U24, new_ADD_371_U25, new_ADD_371_U26, new_ADD_371_U27,
    new_ADD_371_U28, new_ADD_371_U29, new_ADD_371_U30, new_ADD_371_U31,
    new_ADD_371_U32, new_ADD_371_U33, new_ADD_371_U34, new_ADD_371_U35,
    new_ADD_371_U36, new_ADD_371_U37, new_ADD_371_U38, new_ADD_371_U39,
    new_ADD_371_U40, new_ADD_371_U41, new_ADD_371_U42, new_ADD_371_U43,
    new_ADD_371_U44, new_ADD_405_U4, new_ADD_405_U5, new_ADD_405_U6,
    new_ADD_405_U7, new_ADD_405_U8, new_ADD_405_U9, new_ADD_405_U10,
    new_ADD_405_U11, new_ADD_405_U12, new_ADD_405_U13, new_ADD_405_U14,
    new_ADD_405_U15, new_ADD_405_U16, new_ADD_405_U17, new_ADD_405_U18,
    new_ADD_405_U19, new_ADD_405_U20, new_ADD_405_U21, new_ADD_405_U22,
    new_ADD_405_U23, new_ADD_405_U24, new_ADD_405_U25, new_ADD_405_U26,
    new_ADD_405_U27, new_ADD_405_U28, new_ADD_405_U29, new_ADD_405_U30,
    new_ADD_405_U31, new_ADD_405_U32, new_ADD_405_U33, new_ADD_405_U34,
    new_ADD_405_U35, new_ADD_405_U36, new_ADD_405_U37, new_ADD_405_U38,
    new_ADD_405_U39, new_ADD_405_U40, new_ADD_405_U41, new_ADD_405_U42,
    new_ADD_405_U43, new_ADD_405_U44, new_ADD_405_U45, new_ADD_405_U46,
    new_ADD_405_U47, new_ADD_405_U48, new_ADD_405_U49, new_ADD_405_U50,
    new_ADD_405_U51, new_ADD_405_U52, new_ADD_405_U53, new_ADD_405_U54,
    new_ADD_405_U55, new_ADD_405_U56, new_ADD_405_U57, new_ADD_405_U58,
    new_ADD_405_U59, new_ADD_405_U60, new_ADD_405_U61, new_ADD_405_U62,
    new_ADD_405_U63, new_ADD_405_U64, new_ADD_405_U65, new_ADD_405_U66,
    new_ADD_405_U67, new_ADD_405_U68, new_ADD_405_U69, new_ADD_405_U70,
    new_ADD_405_U71, new_ADD_405_U72, new_ADD_405_U73, new_ADD_405_U74,
    new_ADD_405_U75, new_ADD_405_U76, new_ADD_405_U77, new_ADD_405_U78,
    new_ADD_405_U79, new_ADD_405_U80, new_ADD_405_U81, new_ADD_405_U82,
    new_ADD_405_U83, new_ADD_405_U84, new_ADD_405_U85, new_ADD_405_U86,
    new_ADD_405_U87, new_ADD_405_U88, new_ADD_405_U89, new_ADD_405_U90,
    new_ADD_405_U91, new_ADD_405_U92, new_ADD_405_U93, new_ADD_405_U94,
    new_ADD_405_U95, new_ADD_405_U96, new_ADD_405_U97, new_ADD_405_U98,
    new_ADD_405_U99, new_ADD_405_U100, new_ADD_405_U101, new_ADD_405_U102,
    new_ADD_405_U103, new_ADD_405_U104, new_ADD_405_U105, new_ADD_405_U106,
    new_ADD_405_U107, new_ADD_405_U108, new_ADD_405_U109, new_ADD_405_U110,
    new_ADD_405_U111, new_ADD_405_U112, new_ADD_405_U113, new_ADD_405_U114,
    new_ADD_405_U115, new_ADD_405_U116, new_ADD_405_U117, new_ADD_405_U118,
    new_ADD_405_U119, new_ADD_405_U120, new_ADD_405_U121, new_ADD_405_U122,
    new_ADD_405_U123, new_ADD_405_U124, new_ADD_405_U125, new_ADD_405_U126,
    new_ADD_405_U127, new_ADD_405_U128, new_ADD_405_U129, new_ADD_405_U130,
    new_ADD_405_U131, new_ADD_405_U132, new_ADD_405_U133, new_ADD_405_U134,
    new_ADD_405_U135, new_ADD_405_U136, new_ADD_405_U137, new_ADD_405_U138,
    new_ADD_405_U139, new_ADD_405_U140, new_ADD_405_U141, new_ADD_405_U142,
    new_ADD_405_U143, new_ADD_405_U144, new_ADD_405_U145, new_ADD_405_U146,
    new_ADD_405_U147, new_ADD_405_U148, new_ADD_405_U149, new_ADD_405_U150,
    new_ADD_405_U151, new_ADD_405_U152, new_ADD_405_U153, new_ADD_405_U154,
    new_ADD_405_U155, new_ADD_405_U156, new_ADD_405_U157, new_ADD_405_U158,
    new_ADD_405_U159, new_ADD_405_U160, new_ADD_405_U161, new_ADD_405_U162,
    new_ADD_405_U163, new_ADD_405_U164, new_ADD_405_U165, new_ADD_405_U166,
    new_ADD_405_U167, new_ADD_405_U168, new_ADD_405_U169, new_ADD_405_U170,
    new_ADD_405_U171, new_ADD_405_U172, new_ADD_405_U173, new_ADD_405_U174,
    new_ADD_405_U175, new_ADD_405_U176, new_ADD_405_U177, new_ADD_405_U178,
    new_ADD_405_U179, new_ADD_405_U180, new_ADD_405_U181, new_ADD_405_U182,
    new_ADD_405_U183, new_ADD_405_U184, new_ADD_405_U185, new_ADD_405_U186,
    new_GTE_485_U6, new_GTE_485_U7, new_ADD_515_U4, new_ADD_515_U5,
    new_ADD_515_U6, new_ADD_515_U7, new_ADD_515_U8, new_ADD_515_U9,
    new_ADD_515_U10, new_ADD_515_U11, new_ADD_515_U12, new_ADD_515_U13,
    new_ADD_515_U14, new_ADD_515_U15, new_ADD_515_U16, new_ADD_515_U17,
    new_ADD_515_U18, new_ADD_515_U19, new_ADD_515_U20, new_ADD_515_U21,
    new_ADD_515_U22, new_ADD_515_U23, new_ADD_515_U24, new_ADD_515_U25,
    new_ADD_515_U26, new_ADD_515_U27, new_ADD_515_U28, new_ADD_515_U29,
    new_ADD_515_U30, new_ADD_515_U31, new_ADD_515_U32, new_ADD_515_U33,
    new_ADD_515_U34, new_ADD_515_U35, new_ADD_515_U36, new_ADD_515_U37,
    new_ADD_515_U38, new_ADD_515_U39, new_ADD_515_U40, new_ADD_515_U41,
    new_ADD_515_U42, new_ADD_515_U43, new_ADD_515_U44, new_ADD_515_U45,
    new_ADD_515_U46, new_ADD_515_U47, new_ADD_515_U48, new_ADD_515_U49,
    new_ADD_515_U50, new_ADD_515_U51, new_ADD_515_U52, new_ADD_515_U53,
    new_ADD_515_U54, new_ADD_515_U55, new_ADD_515_U56, new_ADD_515_U57,
    new_ADD_515_U58, new_ADD_515_U59, new_ADD_515_U60, new_ADD_515_U61,
    new_ADD_515_U62, new_ADD_515_U63, new_ADD_515_U64, new_ADD_515_U65,
    new_ADD_515_U66, new_ADD_515_U67, new_ADD_515_U68, new_ADD_515_U69,
    new_ADD_515_U70, new_ADD_515_U71, new_ADD_515_U72, new_ADD_515_U73,
    new_ADD_515_U74, new_ADD_515_U75, new_ADD_515_U76, new_ADD_515_U77,
    new_ADD_515_U78, new_ADD_515_U79, new_ADD_515_U80, new_ADD_515_U81,
    new_ADD_515_U82, new_ADD_515_U83, new_ADD_515_U84, new_ADD_515_U85,
    new_ADD_515_U86, new_ADD_515_U87, new_ADD_515_U88, new_ADD_515_U89,
    new_ADD_515_U90, new_ADD_515_U91, new_ADD_515_U92, new_ADD_515_U93,
    new_ADD_515_U94, new_ADD_515_U95, new_ADD_515_U96, new_ADD_515_U97,
    new_ADD_515_U98, new_ADD_515_U99, new_ADD_515_U100, new_ADD_515_U101,
    new_ADD_515_U102, new_ADD_515_U103, new_ADD_515_U104, new_ADD_515_U105,
    new_ADD_515_U106, new_ADD_515_U107, new_ADD_515_U108, new_ADD_515_U109,
    new_ADD_515_U110, new_ADD_515_U111, new_ADD_515_U112, new_ADD_515_U113,
    new_ADD_515_U114, new_ADD_515_U115, new_ADD_515_U116, new_ADD_515_U117,
    new_ADD_515_U118, new_ADD_515_U119, new_ADD_515_U120, new_ADD_515_U121,
    new_ADD_515_U122, new_ADD_515_U123, new_ADD_515_U124, new_ADD_515_U125,
    new_ADD_515_U126, new_ADD_515_U127, new_ADD_515_U128, new_ADD_515_U129,
    new_ADD_515_U130, new_ADD_515_U131, new_ADD_515_U132, new_ADD_515_U133,
    new_ADD_515_U134, new_ADD_515_U135, new_ADD_515_U136, new_ADD_515_U137,
    new_ADD_515_U138, new_ADD_515_U139, new_ADD_515_U140, new_ADD_515_U141,
    new_ADD_515_U142, new_ADD_515_U143, new_ADD_515_U144, new_ADD_515_U145,
    new_ADD_515_U146, new_ADD_515_U147, new_ADD_515_U148, new_ADD_515_U149,
    new_ADD_515_U150, new_ADD_515_U151, new_not_keyinput0,
    new_not_keyinput1, new_not_keyinput2, new_not_0, new_and_1, new_not_2,
    new_and_3, new_not_Q_0, new_not_Q_1, new_count_state_1,
    new_count_state_2, new_count_state_3, new_y_mux_key0_and_0,
    new_y_mux_key0_and_1, new_y_mux_key0, new_y_mux_key1_and_0,
    new_y_mux_key1_and_1, new_y_mux_key1, new_y_mux_key2_and_0,
    new_y_mux_key2_and_1, new_y_mux_key2, new_y_mux_key3_and_0,
    new_y_mux_key3_and_1, new_y_mux_key3, new__state_1, new__state_2,
    new__state_3, new__state_5, new_s__state_1, new_not_s__state_1,
    new_I0__state_1, new_I1__state_1, new_and_mux__state_1,
    new_and_mux__state_1_2, new_y_mux_4, new_s__state_3,
    new_not_s__state_3, new_I0__state_3, new_I1__state_3,
    new_and_mux__state_3, new_and_mux__state_3_2, new_y_mux_5,
    new_s__state_5, new_not_s__state_5, new_I0__state_5, new_I1__state_5,
    new_and_mux__state_5, new_and_mux__state_5_2, n220, n224, n228, n232,
    n236, n240, n244, n248, n252, n256, n260, n264, n268, n272, n276, n280,
    n284, n288, n292, n296, n300, n304, n308, n312, n316, n320, n324, n328,
    n332, n336, n340, n344, n348, n352, n356, n361, n366, n371, n376, n381,
    n386, n391, n396, n401, n406, n411, n416, n421, n426, n431, n436, n441,
    n446, n451, n456, n461, n466, n471, n476, n481, n486, n491, n496, n501,
    n506, n511, n516, n521, n526, n531, n536, n541, n546, n551, n556, n561,
    n566, n571, n576, n581, n586, n591, n596, n601, n606, n611, n616, n621,
    n626, n631, n636, n641, n646, n651, n656, n661, n666, n671, n676, n681,
    n686, n691, n696, n701, n706, n711, n716, n721, n726, n731, n736, n741,
    n746, n751, n756, n761, n766, n771, n776, n781, n786, n791, n796, n801,
    n806, n811, n816, n821, n826, n831, n836, n841, n846, n851, n856, n861,
    n866, n871, n876, n881, n886, n891, n896, n901, n906, n911, n916, n921,
    n926, n931, n936, n941, n946, n951, n956, n961, n966, n971, n976, n981,
    n986, n991, n996, n1001, n1006, n1011, n1016, n1021, n1026, n1031,
    n1036, n1041, n1046, n1051, n1056, n1061, n1066, n1071, n1076, n1081,
    n1086, n1091, n1096, n1101, n1106, n1111, n1116, n1121, n1126, n1131,
    n1136, n1141, n1146, n1151, n1156, n1161, n1166, n1171, n1176, n1181,
    n1186, n1191, n1196, n1201, n1206, n1211, n1216, n1221, n1226, n1231,
    n1236, n1241, n1246, n1251, n1256, n1261, n1266, n1271, n1276, n1281,
    n1286, n1291, n1296, n1301, n1306, n1311, n1316, n1321, n1326, n1331,
    n1336, n1341, n1346, n1351, n1356, n1361, n1366, n1371, n1376, n1381,
    n1386, n1391, n1396, n1401, n1406, n1411, n1416, n1421, n1426, n1431,
    n1436, n1441, n1446, n1451, n1456, n1461, n1466, n1471, n1476, n1481,
    n1486, n1491, n1496, n1501, n1506, n1511, n1516, n1521, n1526, n1531,
    n1536, n1541, n1546, n1551, n1556, n1561, n1566, n1571, n1576, n1581,
    n1586, n1591, n1596, n1601, n1606, n1611, n1616, n1621, n1626, n1631,
    n1636, n1641, n1646, n1651, n1656, n1661, n1666, n1671, n1676, n1681,
    n1686, n1691, n1696, n1701, n1706, n1711, n1716, n1720, n1724, n1728,
    n1732, n1736, n1740, n1744, n1748, n1752, n1756, n1760, n1764, n1768,
    n1772, n1776, n1780, n1784, n1788, n1792, n1796, n1800, n1804, n1808,
    n1812, n1816, n1820, n1824, n1828, n1832, n1836, n1840, n1844, n1849,
    n1854, n1859, n1864, n1869, n1874, n1879, n1884, n1889, n1894, n1899,
    n1904, n1909, n1914, n1919, n1924, n1929, n1934, n1939, n1944, n1949,
    n1954, n1959, n1964, n1969, n1974, n1979, n1984, n1989, n1994, n1999,
    n2004, n2009, n2014, n2019, n2024, n2029, n2034, n2039, n2044, n2049,
    n2054, n2059, n2064, n2069, n2074, n2079, n2084, n2089, n2094, n2099,
    n2104, n2109, n2114, n2119, n2124, n2129, n2134, n2139, n2144, n2149,
    n2154, n2159, n2164, n2169, n2174, n2179, n2184, n2189, n2194, n2199,
    n2204, n2209, n2214, n2219, n2224, n2229, n2234, n2239, n2244, n2249,
    n2254, n2259, n2264, n2269, n2274, n2279, n2284, n2289, n2294, n2299,
    n2304, n2309, n2314, n2319, n2324, n2329, n2334, n2339, n2344, n2348,
    n2353, n2358, n2363, n2368, n2372, n2376, n2381, n2385, n2390, n18700,
    n18703;
  assign new_ADD_515_U182 = ~new_ADD_515_U101 | ~new_ADD_515_U21;
  assign new_ADD_515_U181 = ~INSTADDRPOINTER_REG_10_ | ~new_ADD_515_U20;
  assign new_ADD_515_U180 = ~new_ADD_515_U102 | ~new_ADD_515_U23;
  assign new_U2352 = ~STATEBS16_REG & ~STATE2_REG_2_;
  assign new_U2353 = new_U4219 & STATE2_REG_2_;
  assign new_U2354 = new_U4253 & new_U4465;
  assign new_U2355 = new_U3221 & new_U2450;
  assign new_U2356 = new_R2238_U6 & new_U4180;
  assign new_U2357 = new_R2167_U17 & new_U5947 & new_U3853;
  assign new_U2358 = new_U2388 & new_U4212;
  assign new_U2359 = STATE2_REG_2_ & new_U3418;
  assign new_U2360 = STATE2_REG_2_ & new_U3401;
  assign new_U2361 = new_U4212 & STATE2_REG_3_;
  assign new_U2362 = new_U2359 & new_U4196;
  assign new_U2363 = new_U2359 & new_U4198;
  assign new_U2364 = new_U3852 & new_U3403;
  assign new_U2365 = new_U4249 & new_U3403;
  assign new_U2366 = new_U3417 & new_U3418 & STATE2_REG_1_;
  assign new_U2367 = new_R2337_U58 & STATE2_REG_1_ & new_U3418;
  assign new_U2368 = new_U4223 & STATE2_REG_0_;
  assign new_U2369 = new_U2362 & new_U4485;
  assign new_U2370 = new_U3401 & new_U3250;
  assign new_U2371 = new_U4210 & new_U4437;
  assign new_U2372 = STATE2_REG_0_ & new_U3403;
  assign new_U2373 = STATE2_REG_3_ & new_U3418;
  assign new_U2374 = new_U2360 & new_U4202;
  assign new_U2375 = new_U2360 & new_U4204;
  assign new_U2376 = new_U5786 & new_U3403;
  assign new_U2377 = new_U3750 & new_U3401;
  assign new_U2378 = new_U2360 & new_U5557;
  assign new_U2379 = new_U2363 & new_U3267;
  assign new_U2380 = new_U2360 & new_U7596;
  assign new_U2381 = new_U2357 & new_U3258;
  assign new_U2382 = new_U2357 & new_U4465;
  assign new_U2383 = new_U4210 & new_U3378;
  assign new_U2384 = STATE2_REG_0_ & new_U3404;
  assign new_U2385 = new_U3404 & new_U3281;
  assign new_U2386 = new_U4211 & new_U3410;
  assign new_U2387 = new_U3872 & new_U4211;
  assign new_U2388 = STATEBS16_REG & new_U4197;
  assign new_U2389 = new_U2452 & new_U7482;
  assign new_U2390 = DATAI_0_ & new_U4212;
  assign new_U2391 = DATAI_1_ & new_U4212;
  assign new_U2392 = DATAI_2_ & new_U4212;
  assign new_U2393 = DATAI_3_ & new_U4212;
  assign new_U2394 = DATAI_4_ & new_U4212;
  assign new_U2395 = DATAI_5_ & new_U4212;
  assign new_U2396 = DATAI_6_ & new_U4212;
  assign new_U2397 = DATAI_7_ & new_U4212;
  assign new_U2398 = DATAI_24_ & new_U2358;
  assign new_U2399 = DATAI_16_ & new_U2358;
  assign new_U2400 = DATAI_25_ & new_U2358;
  assign new_U2401 = DATAI_17_ & new_U2358;
  assign new_U2402 = DATAI_26_ & new_U2358;
  assign new_U2403 = DATAI_18_ & new_U2358;
  assign new_U2404 = DATAI_27_ & new_U2358;
  assign new_U2405 = DATAI_19_ & new_U2358;
  assign new_U2406 = DATAI_28_ & new_U2358;
  assign new_U2407 = DATAI_20_ & new_U2358;
  assign new_U2408 = DATAI_29_ & new_U2358;
  assign new_U2409 = DATAI_21_ & new_U2358;
  assign new_U2410 = DATAI_30_ & new_U2358;
  assign new_U2411 = DATAI_22_ & new_U2358;
  assign new_U2412 = DATAI_31_ & new_U2358;
  assign new_U2413 = DATAI_23_ & new_U2358;
  assign new_U2414 = new_U2361 & new_U3258;
  assign new_U2415 = new_U2361 & new_U3378;
  assign new_U2416 = new_U2361 & new_U3264;
  assign new_U2417 = new_U2361 & new_U3271;
  assign new_U2418 = new_U2361 & new_U3270;
  assign new_U2419 = new_U2361 & new_U3265;
  assign new_U2420 = new_U2361 & new_U4161;
  assign new_U2421 = new_U2361 & new_U4159;
  assign new_U2422 = new_U4211 & new_U5449;
  assign new_U2423 = new_U4211 & new_U4219;
  assign new_U2424 = new_U2384 & new_U3271;
  assign new_U2425 = new_U2368 & new_U2448;
  assign new_U2426 = new_U3877 & new_U3418;
  assign new_U2427 = ~STATE2_REG_1_ & ~STATE2_REG_3_;
  assign new_U2428 = STATE2_REG_2_ & STATE2_REG_1_;
  assign new_U2429 = new_U6354 & new_U3418;
  assign new_U2430 = STATE2_REG_1_ & new_U3374;
  assign new_U2431 = new_U4187 & new_U7482;
  assign new_U2432 = new_U3442 & new_U3347;
  assign new_U2433 = new_U4528 & new_U3442;
  assign new_U2434 = new_U7684 & new_U3347;
  assign new_U2435 = new_U4528 & new_U7684;
  assign new_U2436 = new_U3222 & new_U3288;
  assign new_U2437 = new_U4531 & new_U3288;
  assign new_U2438 = new_R2182_U42 & new_R2182_U25;
  assign new_U2439 = new_R2182_U42 & new_U3303;
  assign new_U2440 = new_R2182_U25 & new_U3304;
  assign new_U2441 = ~new_R2182_U42 & ~new_R2182_U25;
  assign new_U2442 = new_R2182_U33 & new_R2182_U34;
  assign new_U2443 = new_R2182_U33 & new_U3305;
  assign new_U2444 = new_R2182_U34 & new_U3306;
  assign new_U2445 = ~new_R2182_U33 & ~new_R2182_U34;
  assign new_U2446 = STATE2_REG_1_ & new_U3458;
  assign new_U2447 = new_U3565 & new_U2452;
  assign new_U2448 = new_R2167_U17 & new_U3271;
  assign new_U2449 = new_U4482 & new_U3258;
  assign new_U2450 = STATE2_REG_0_ & new_U4388;
  assign new_U2451 = new_U4239 & STATE2_REG_0_;
  assign new_U2452 = new_U4161 & new_U3378 & new_U4388 & new_U3264;
  assign new_U2453 = INSTQUEUERD_ADDR_REG_2_ & INSTQUEUERD_ADDR_REG_1_ & INSTQUEUERD_ADDR_REG_3_ & INSTQUEUERD_ADDR_REG_0_;
  assign new_U2454 = INSTQUEUERD_ADDR_REG_1_ & new_U3253;
  assign new_U2455 = new_U3253 & INSTQUEUERD_ADDR_REG_2_ & INSTQUEUERD_ADDR_REG_3_ & INSTQUEUERD_ADDR_REG_1_;
  assign new_U2456 = INSTQUEUERD_ADDR_REG_0_ & new_U3252;
  assign new_U2457 = new_U3252 & INSTQUEUERD_ADDR_REG_2_ & INSTQUEUERD_ADDR_REG_3_ & INSTQUEUERD_ADDR_REG_0_;
  assign new_U2458 = new_U3495 & new_U4366;
  assign new_U2459 = new_U3251 & INSTQUEUERD_ADDR_REG_1_ & INSTQUEUERD_ADDR_REG_3_ & INSTQUEUERD_ADDR_REG_0_;
  assign new_U2460 = INSTQUEUERD_ADDR_REG_1_ & new_U3251 & new_U3253;
  assign new_U2461 = new_U3494 & new_U3493;
  assign new_U2462 = INSTQUEUERD_ADDR_REG_0_ & new_U3251 & new_U3252;
  assign new_U2463 = new_U3492 & new_U3491;
  assign new_U2464 = INSTQUEUERD_ADDR_REG_3_ & new_U4368;
  assign new_U2465 = new_U3490 & new_U3489;
  assign new_U2466 = new_U3488 & new_U3487;
  assign new_U2467 = new_U4366 & INSTQUEUERD_ADDR_REG_2_ & new_U3257;
  assign new_U2468 = new_U3486 & new_U3485;
  assign new_U2469 = ~INSTQUEUERD_ADDR_REG_3_ & ~INSTQUEUERD_ADDR_REG_2_;
  assign new_U2470 = new_U2469 & INSTQUEUERD_ADDR_REG_1_ & new_U3253;
  assign new_U2471 = new_U2469 & INSTQUEUERD_ADDR_REG_0_ & new_U3252;
  assign new_U2472 = new_U4368 & new_U3257;
  assign new_U2473 = new_U3393 & new_U7668 & new_U7667;
  assign new_U2474 = new_R2144_U49 & new_U3299;
  assign new_U2475 = new_U3441 & new_U3345;
  assign new_U2476 = new_R2144_U8 & new_R2144_U49;
  assign new_U2477 = new_U4516 & new_U2476;
  assign new_U2478 = INSTQUEUEWR_ADDR_REG_2_ & INSTQUEUEWR_ADDR_REG_3_;
  assign new_U2479 = INSTQUEUEWR_ADDR_REG_2_ & new_U3290;
  assign new_U2480 = new_U3302 & new_U4536;
  assign new_U2481 = new_U4512 & new_U2476;
  assign new_U2482 = new_U3314 & new_U4594;
  assign new_U2483 = new_U4513 & new_U2476;
  assign new_U2484 = new_U3321 & new_U4653;
  assign new_U2485 = new_U4514 & new_R2144_U43;
  assign new_U2486 = ~new_R2144_U43 & ~new_R2144_U50;
  assign new_U2487 = new_U2486 & new_U2476;
  assign new_U2488 = ~INSTQUEUEWR_ADDR_REG_0_ & ~INSTQUEUEWR_ADDR_REG_1_;
  assign new_U2489 = new_U3325 & new_U4710;
  assign new_U2490 = new_U7681 & new_U3345;
  assign new_U2491 = new_U4517 & new_U4516;
  assign new_U2492 = new_U3330 & new_U4768;
  assign new_U2493 = new_U4517 & new_U4512;
  assign new_U2494 = new_U3334 & new_U4825;
  assign new_U2495 = new_U4517 & new_U4513;
  assign new_U2496 = new_U3337 & new_U4883;
  assign new_U2497 = new_U4517 & new_U2486;
  assign new_U2498 = new_U3341 & new_U4940;
  assign new_U2499 = new_U4519 & new_U3441;
  assign new_U2500 = new_U3346 & new_U3344;
  assign new_U2501 = new_U4512 & new_U2474;
  assign new_U2502 = new_U3351 & new_U5053;
  assign new_U2503 = new_U4513 & new_U2474;
  assign new_U2504 = new_U3354 & new_U5111;
  assign new_U2505 = new_U2486 & new_U2474;
  assign new_U2506 = new_U3358 & new_U5168;
  assign new_U2507 = new_U4519 & new_U7681;
  assign new_U2508 = ~new_R2144_U49 & ~new_R2144_U8;
  assign new_U2509 = new_U2508 & new_U4516;
  assign new_U2510 = ~INSTQUEUEWR_ADDR_REG_3_ & ~INSTQUEUEWR_ADDR_REG_2_;
  assign new_U2511 = new_U3361 & new_U5226;
  assign new_U2512 = new_U2508 & new_U4512;
  assign new_U2513 = new_U3365 & new_U5283;
  assign new_U2514 = new_U2508 & new_U4513;
  assign new_U2515 = new_U3368 & new_U5341;
  assign new_U2516 = new_U2508 & new_U2486;
  assign new_U2517 = new_U3372 & new_U5398;
  assign new_U2518 = new_U5456 & new_U7688 & new_U7687;
  assign new_U2519 = new_U3732 & new_U5487;
  assign new_U2520 = new_U4207 & new_U3433;
  assign new_U2521 = INSTQUEUERD_ADDR_REG_0_ & new_U3389;
  assign new_U2522 = new_U5471 & new_U5499;
  assign new_U2523 = new_U2522 & new_U2521;
  assign new_U2524 = new_U3253 & new_U3389;
  assign new_U2525 = new_U2522 & new_U2524;
  assign new_U2526 = new_U5507 & INSTQUEUERD_ADDR_REG_0_;
  assign new_U2527 = new_U2522 & new_U2526;
  assign new_U2528 = new_U5507 & new_U3253;
  assign new_U2529 = new_U2522 & new_U2528;
  assign new_U2530 = new_U5471 & new_U3388;
  assign new_U2531 = new_U2530 & new_U2521;
  assign new_U2532 = new_U2530 & new_U2524;
  assign new_U2533 = new_U2530 & new_U2526;
  assign new_U2534 = new_U2530 & new_U2528;
  assign new_U2535 = new_U5499 & new_U3425;
  assign new_U2536 = new_U2535 & new_U2521;
  assign new_U2537 = new_U2535 & new_U2524;
  assign new_U2538 = new_U2535 & new_U2526;
  assign new_U2539 = new_U2535 & new_U2528;
  assign new_U2540 = new_U3425 & new_U3388;
  assign new_U2541 = new_U2521 & new_U2540;
  assign new_U2542 = new_U2524 & new_U2540;
  assign new_U2543 = new_U2526 & new_U2540;
  assign new_U2544 = new_U2528 & new_U2540;
  assign new_U2545 = new_U5468 & new_U7708;
  assign new_U2546 = new_U2545 & new_U2454;
  assign new_U2547 = new_U2545 & new_U3486;
  assign new_U2548 = new_U2545 & new_U4366;
  assign new_U2549 = new_U2545 & new_U2456;
  assign new_U2550 = new_U5468 & new_U3443;
  assign new_U2551 = new_U2550 & new_U2454;
  assign new_U2552 = new_U2550 & new_U3486;
  assign new_U2553 = new_U2550 & new_U4366;
  assign new_U2554 = new_U2550 & new_U2456;
  assign new_U2555 = new_U7708 & new_U3429;
  assign new_U2556 = new_U2555 & new_U2454;
  assign new_U2557 = new_U2555 & new_U3486;
  assign new_U2558 = new_U2555 & new_U4366;
  assign new_U2559 = new_U2555 & new_U2456;
  assign new_U2560 = new_U3443 & new_U3429;
  assign new_U2561 = new_U2560 & new_U2454;
  assign new_U2562 = new_U2560 & new_U3486;
  assign new_U2563 = new_U2560 & new_U4366;
  assign new_U2564 = new_U2560 & new_U2456;
  assign new_U2565 = new_U7053 & new_U4367;
  assign new_U2566 = new_U7053 & new_U2460;
  assign new_U2567 = new_U7053 & new_U2462;
  assign new_U2568 = new_U7053 & new_U4368;
  assign new_U2569 = new_U7053 & INSTQUEUERD_ADDR_REG_2_;
  assign new_U2570 = new_U2569 & new_U3486;
  assign new_U2571 = new_U2569 & new_U2454;
  assign new_U2572 = new_U2569 & new_U2456;
  assign new_U2573 = new_U2569 & new_U4366;
  assign new_U2574 = new_U4367 & new_U3432;
  assign new_U2575 = new_U2460 & new_U3432;
  assign new_U2576 = new_U2462 & new_U3432;
  assign new_U2577 = new_U4368 & new_U3432;
  assign new_U2578 = INSTQUEUERD_ADDR_REG_2_ & new_U3432;
  assign new_U2579 = new_U2578 & new_U3486;
  assign new_U2580 = new_U2578 & new_U2454;
  assign new_U2581 = new_U2578 & new_U2456;
  assign new_U2582 = new_U2578 & new_U4366;
  assign new_U2583 = new_U7778 & new_U4172;
  assign new_U2584 = new_U2583 & new_U2524;
  assign new_U2585 = new_U2583 & new_U2521;
  assign new_U2586 = new_U2583 & new_U2528;
  assign new_U2587 = new_U2583 & new_U2526;
  assign new_U2588 = new_U7778 & new_U3439;
  assign new_U2589 = new_U2588 & new_U2524;
  assign new_U2590 = new_U2588 & new_U2521;
  assign new_U2591 = new_U2588 & new_U2528;
  assign new_U2592 = new_U2588 & new_U2526;
  assign new_U2593 = new_U4172 & new_U3444;
  assign new_U2594 = new_U2593 & new_U2524;
  assign new_U2595 = new_U2593 & new_U2521;
  assign new_U2596 = new_U2593 & new_U2528;
  assign new_U2597 = new_U2593 & new_U2526;
  assign new_U2598 = new_U3444 & new_U3439;
  assign new_U2599 = new_U2598 & new_U2524;
  assign new_U2600 = new_U2598 & new_U2521;
  assign new_U2601 = new_U2598 & new_U2528;
  assign new_U2602 = new_U2598 & new_U2526;
  assign new_U2603 = STATE2_REG_0_ & new_U3376;
  assign new_U2604 = EBX_REG_31_ & new_U2379;
  assign new_U2605 = new_U3518 & new_U3519 & new_U3520 & new_U3521 & new_U2607;
  assign new_U2606 = new_U7492 & new_U3414;
  assign new_U2607 = new_U7660 & new_U7659;
  assign new_U2608 = new_U7775 & new_U7774;
  assign new_U2609 = ~new_U6744 | ~new_U3993;
  assign new_U2610 = ~new_U6741 | ~new_U3992;
  assign new_U2611 = ~new_U6738 | ~new_U3991;
  assign new_U2612 = ~new_U6735 | ~new_U3990;
  assign new_U2613 = ~new_U6844 | ~new_U4014;
  assign new_U2614 = ~new_U6843 | ~new_U6841 | ~new_U6842;
  assign new_U2615 = ~new_U6840 | ~new_U6838 | ~new_U6839;
  assign new_U2616 = ~new_U6837 | ~new_U6835 | ~new_U6836;
  assign new_U2617 = ~new_U6834 | ~new_U6832 | ~new_U6833;
  assign new_U2618 = ~new_U6831 | ~new_U6829 | ~new_U6830;
  assign new_ADD_515_U179 = ~INSTADDRPOINTER_REG_11_ | ~new_ADD_515_U22;
  assign new_U2620 = new_R2144_U145 & new_U6734;
  assign new_U2621 = new_R2144_U145 & new_U6734;
  assign new_U2622 = new_R2144_U145 & new_U6734;
  assign new_U2623 = new_R2144_U145 & new_U6734;
  assign new_U2624 = new_R2144_U145 & new_U6734;
  assign new_U2625 = new_R2144_U145 & new_U6734;
  assign new_U2626 = new_R2144_U145 & new_U6734;
  assign new_U2627 = new_R2144_U145 & new_U6734;
  assign new_U2628 = new_R2144_U145 & new_U6734;
  assign new_U2629 = new_R2144_U145 & new_U6734;
  assign new_U2630 = new_R2144_U145 & new_U6734;
  assign new_U2631 = new_R2144_U145 & new_U6734;
  assign new_U2632 = new_R2144_U145 & new_U6734;
  assign new_U2633 = new_R2144_U145 & new_U6734;
  assign new_U2634 = new_R2144_U11 & new_U6734;
  assign new_U2635 = new_R2144_U37 & new_U6734;
  assign new_U2636 = new_R2144_U38 & new_U6734;
  assign new_U2637 = new_R2144_U39 & new_U6734;
  assign new_U2638 = new_R2144_U40 & new_U6734;
  assign new_U2639 = new_R2144_U41 & new_U6734;
  assign new_U2640 = new_R2144_U42 & new_U6734;
  assign new_U2641 = new_R2144_U30 & new_U6734;
  assign new_U2642 = new_R2144_U80 & new_U6734;
  assign new_U2643 = new_R2144_U10 & new_U6734;
  assign new_U2644 = new_R2144_U9 & new_U6734;
  assign new_U2645 = new_R2144_U45 & new_U6734;
  assign new_U2646 = new_R2144_U47 & new_U6734;
  assign new_U2647 = new_R2144_U8 & new_U6734;
  assign new_U2648 = ~new_U3427 | ~new_U6857;
  assign new_U2649 = new_R2144_U50 & new_U6734;
  assign new_U2650 = STATE2_REG_2_ & new_U6858;
  assign new_U2651 = ~new_U6758 | ~new_U6757 | ~new_U6756;
  assign new_U2652 = ~new_U6759 | ~new_U3997;
  assign new_U2653 = ~new_U6768 | ~new_U3999;
  assign new_U2654 = ~new_U6772 | ~new_U4000;
  assign new_U2655 = ~new_U6776 | ~new_U4001;
  assign new_U2656 = ~new_U6780 | ~new_U4002;
  assign new_U2657 = ~new_U6784 | ~new_U4003;
  assign new_U2658 = ~new_U6788 | ~new_U4004;
  assign new_U2659 = ~new_U6792 | ~new_U4005;
  assign new_U2660 = ~new_U6796 | ~new_U4006;
  assign new_U2661 = ~new_U6800 | ~new_U4007;
  assign new_U2662 = ~new_U6804 | ~new_U4008;
  assign new_U2663 = ~new_U6813 | ~new_U4010;
  assign new_U2664 = ~new_U6817 | ~new_U4011;
  assign new_U2665 = ~new_U6821 | ~new_U4012;
  assign new_U2666 = ~new_U6825 | ~new_U4013;
  assign new_U2667 = ~new_U6747 | ~new_U3994;
  assign new_U2668 = ~new_U6751 | ~new_U3996 | ~new_U6755 | ~new_U6754;
  assign new_U2669 = ~new_U6763 | ~new_U3998 | ~new_U6767 | ~new_U6766;
  assign new_U2670 = ~new_U6808 | ~new_U4009 | ~new_U6812 | ~new_U6811;
  assign new_U2671 = ~new_U6847 | ~new_U4015 | ~new_U6851 | ~new_U6850;
  assign new_U2672 = ~new_U6855 | ~new_U6856 | ~new_U6853 | ~new_U6854 | ~new_U6852;
  assign new_U2673 = ~new_U7446 | ~new_U7445;
  assign new_U2674 = ~new_U7448 | ~new_U7447;
  assign new_U2675 = ~new_U4156 | ~new_U7451;
  assign new_U2676 = ~new_U4157 | ~new_U7454;
  assign new_U2677 = ~new_U7455 | ~new_U7782 | ~new_U7781;
  assign new_U2678 = ~new_U7444 | ~new_U3271;
  assign new_U2679 = ~new_U7393 | ~new_U7392;
  assign new_U2680 = ~new_U7395 | ~new_U7394;
  assign new_U2681 = ~new_U7399 | ~new_U7398;
  assign new_U2682 = ~new_U7401 | ~new_U7400;
  assign new_U2683 = ~new_U7403 | ~new_U7402;
  assign new_U2684 = ~new_U7405 | ~new_U7404;
  assign new_U2685 = ~new_U7407 | ~new_U7406;
  assign new_U2686 = ~new_U7409 | ~new_U7408;
  assign new_U2687 = ~new_U7411 | ~new_U7410;
  assign new_U2688 = ~new_U7413 | ~new_U7412;
  assign new_U2689 = ~new_U7415 | ~new_U7414;
  assign new_U2690 = ~new_U7417 | ~new_U7416;
  assign new_U2691 = ~new_U7421 | ~new_U7420;
  assign new_U2692 = ~new_U7423 | ~new_U7422;
  assign new_U2693 = ~new_U7425 | ~new_U7424;
  assign new_U2694 = ~new_U7427 | ~new_U7426;
  assign new_U2695 = ~new_U7429 | ~new_U7428;
  assign new_U2696 = ~new_U7431 | ~new_U7430;
  assign new_U2697 = ~new_U7433 | ~new_U7432;
  assign new_U2698 = ~new_U7435 | ~new_U7434;
  assign new_U2699 = ~new_U7437 | ~new_U7436;
  assign new_U2700 = ~new_U7439 | ~new_U7438;
  assign new_U2701 = ~new_U7381 | ~new_U7380;
  assign new_U2702 = ~new_U7383 | ~new_U7382;
  assign new_U2703 = ~new_U7385 | ~new_U7384;
  assign new_U2704 = ~new_U7387 | ~new_U7386;
  assign new_U2705 = ~new_U7389 | ~new_U7388;
  assign new_U2706 = ~new_U7391 | ~new_U7390;
  assign new_U2707 = ~new_U7397 | ~new_U7396;
  assign new_U2708 = ~new_U7419 | ~new_U7418;
  assign new_U2709 = ~new_U7441 | ~new_U7440;
  assign new_U2710 = ~new_U7443 | ~new_U7442;
  assign new_U2711 = ~new_U7365 | ~new_U7364;
  assign new_U2712 = ~new_U7367 | ~new_U7366;
  assign new_U2713 = ~new_U4153 | ~new_U4227;
  assign new_U2714 = ~new_U3421 | ~new_U4154 | ~new_U7374 | ~new_U7373;
  assign new_U2715 = ~new_U4227 | ~new_U4155;
  assign new_U2716 = ~new_U7353 | ~new_U7352;
  assign new_U2717 = ~new_U7355 | ~new_U7354;
  assign new_U2718 = ~new_U4149 | ~new_U7356;
  assign new_U2719 = ~new_U4150 | ~new_U7358;
  assign new_U2720 = ~new_U4151 | ~new_U7360;
  assign new_U2721 = ~new_U4152 | ~new_U7362;
  assign new_U2722 = ~new_U4147 | ~new_U4180;
  assign new_U2723 = new_U7224 & new_U7071;
  assign new_U2724 = new_U7241 & new_U7071;
  assign new_U2725 = new_U7258 & new_U7071;
  assign new_U2726 = new_U7608 & new_U7071;
  assign new_U2727 = new_U7290 & new_U7071;
  assign new_U2728 = new_U7307 & new_U7071;
  assign new_U2729 = new_U7324 & new_U7071;
  assign new_U2730 = new_U7341 & new_U7071;
  assign new_U2731 = ~new_U2606 | ~new_U7342;
  assign new_U2732 = new_U7071 & new_U7070;
  assign new_U2733 = new_U7102 & new_U7071;
  assign new_U2734 = new_U7119 & new_U7071;
  assign new_U2735 = new_U7606 & new_U7071;
  assign new_U2736 = new_U7151 & new_U7071;
  assign new_U2737 = new_U7168 & new_U7071;
  assign new_U2738 = new_U7185 & new_U7071;
  assign new_U2739 = new_U7202 & new_U7071;
  assign new_U2740 = INSTQUEUERD_ADDR_REG_4_ & new_U7051;
  assign new_U2741 = ~new_U4066 | ~new_U7084;
  assign new_U2742 = new_U7480 & new_U7479;
  assign new_U2743 = new_U7494 & new_U7458;
  assign new_U2744 = new_U7467 & new_U7466;
  assign new_U2745 = ~new_U7036 | ~new_U7035;
  assign new_U2746 = ~new_U7038 | ~new_U7037;
  assign new_U2747 = ~new_U7040 | ~new_U7039;
  assign new_U2748 = ~new_U7604 | ~new_U7041;
  assign new_U2749 = ~new_U7043 | ~new_U7042;
  assign new_U2750 = ~new_U7045 | ~new_U7044;
  assign new_U2751 = ~new_U4049 | ~new_U7046;
  assign new_U2752 = ~new_U7049 | ~new_U4050 | ~new_U7048;
  assign new_U2753 = new_U6945 & new_U6897;
  assign new_U2754 = new_U6962 & new_U6897;
  assign new_U2755 = new_U6979 & new_U6897;
  assign new_U2756 = new_U7603 & new_U6897;
  assign new_U2757 = new_U7011 & new_U6897;
  assign new_U2758 = new_U7028 & new_U6897;
  assign new_U2759 = new_U6897 & new_U6896;
  assign new_U2760 = new_U6914 & new_U6897;
  assign new_U2761 = ~new_U6916 | ~new_U6915;
  assign new_U2762 = ~new_U6918 | ~new_U6917;
  assign new_U2763 = ~new_U6920 | ~new_U6919;
  assign new_U2764 = ~new_U6922 | ~new_U6921;
  assign new_U2765 = ~new_U6925 | ~new_U6924 | ~new_U6923;
  assign new_U2766 = ~new_U6928 | ~new_U6927 | ~new_U6926;
  assign new_U2767 = ~new_U7030 | ~new_U7031 | ~new_U7029;
  assign new_U2768 = ~new_U7033 | ~new_U7034 | ~new_U7032;
  assign new_U2769 = new_R2144_U145 & new_U4147;
  assign new_U2770 = new_U4147 & new_R2144_U145;
  assign new_U2771 = new_U4147 & new_R2144_U11;
  assign new_U2772 = new_U4147 & new_R2144_U37;
  assign new_U2773 = new_U4147 & new_R2144_U38;
  assign new_U2774 = new_U4147 & new_R2144_U39;
  assign new_U2775 = new_U4147 & new_R2144_U40;
  assign new_U2776 = new_U4147 & new_R2144_U41;
  assign new_U2777 = new_U4147 & new_R2144_U42;
  assign new_U2778 = new_U4147 & new_R2144_U30;
  assign new_U2779 = ~new_U6860 | ~new_U6859;
  assign new_U2780 = ~new_U6862 | ~new_U6861;
  assign new_U2781 = ~new_U6864 | ~new_U6863;
  assign new_U2782 = ~new_U6866 | ~new_U6865;
  assign new_U2783 = ~new_U6868 | ~new_U6867;
  assign new_U2784 = ~new_U6870 | ~new_U6869;
  assign new_U2785 = ~new_U6871 | ~new_U6872 | ~new_U6873;
  assign new_U2786 = ~new_U6874 | ~new_U4016 | ~new_U6875;
  assign new_U2787 = ~new_U6877 | ~new_U6878 | ~new_U6879;
  assign n2390 = ~new_U7486 | ~new_U6605 | ~new_U3419;
  assign n2381 = ~new_U7638 | ~new_U6601;
  assign n2376 = ~new_U6600 | ~new_U6599;
  assign n2368 = ~new_U4231 | ~new_U7757 | ~new_U7756;
  assign n2358 = ~new_U4231 | ~new_U7753 | ~new_U7752;
  assign n2348 = ~new_U6589 | ~new_U4236;
  assign n2334 = ~new_U4228 | ~new_U7745 | ~new_U7744;
  assign n2324 = ~new_U4228 | ~new_U7735 | ~new_U7734;
  assign n2319 = ~new_U6583 | ~new_U6579 | ~new_U3937 | ~new_U6581 | ~new_U3936;
  assign n2314 = ~new_U6576 | ~new_U6572 | ~new_U3935 | ~new_U6574 | ~new_U3934;
  assign n2309 = ~new_U6569 | ~new_U6565 | ~new_U3933 | ~new_U6567 | ~new_U3932;
  assign n2304 = ~new_U6562 | ~new_U6558 | ~new_U3931 | ~new_U6560 | ~new_U3930;
  assign n2299 = ~new_U6555 | ~new_U6551 | ~new_U3929 | ~new_U6553 | ~new_U3928;
  assign n2294 = ~new_U6548 | ~new_U6544 | ~new_U3927 | ~new_U6546 | ~new_U3926;
  assign n2289 = ~new_U6541 | ~new_U6537 | ~new_U3925 | ~new_U6539 | ~new_U3924;
  assign n2284 = ~new_U6534 | ~new_U6530 | ~new_U3923 | ~new_U6532 | ~new_U3922;
  assign n2279 = ~new_U6527 | ~new_U6523 | ~new_U3921 | ~new_U6525 | ~new_U3920;
  assign n2274 = ~new_U6520 | ~new_U6516 | ~new_U3919 | ~new_U6518 | ~new_U3918;
  assign n2269 = ~new_U6513 | ~new_U6509 | ~new_U3917 | ~new_U6511 | ~new_U3916;
  assign n2264 = ~new_U6506 | ~new_U6502 | ~new_U3915 | ~new_U6504 | ~new_U3914;
  assign n2259 = ~new_U6499 | ~new_U6495 | ~new_U3913 | ~new_U3912 | ~new_U6497;
  assign n2254 = ~new_U6492 | ~new_U6488 | ~new_U3911 | ~new_U3910 | ~new_U6490;
  assign n2249 = ~new_U6485 | ~new_U6481 | ~new_U3909 | ~new_U3908 | ~new_U6483;
  assign n2244 = ~new_U6478 | ~new_U3906 | ~new_U3907 | ~new_U6476 | ~new_U6475;
  assign n2239 = ~new_U6471 | ~new_U3904 | ~new_U3905 | ~new_U6469 | ~new_U6468;
  assign n2234 = ~new_U6464 | ~new_U6461 | ~new_U3902 | ~new_U3903 | ~new_U6462;
  assign n2229 = ~new_U6457 | ~new_U6454 | ~new_U3900 | ~new_U3901 | ~new_U6455;
  assign n2224 = ~new_U6450 | ~new_U6447 | ~new_U3898 | ~new_U3899 | ~new_U6448;
  assign n2219 = ~new_U6443 | ~new_U6440 | ~new_U3896 | ~new_U3897 | ~new_U6441;
  assign n2214 = ~new_U6436 | ~new_U6433 | ~new_U3894 | ~new_U3895 | ~new_U6434;
  assign n2209 = ~new_U6429 | ~new_U6426 | ~new_U3892 | ~new_U3893 | ~new_U6427;
  assign n2204 = ~new_U6422 | ~new_U6419 | ~new_U3890 | ~new_U3891 | ~new_U6420;
  assign n2199 = ~new_U6415 | ~new_U6412 | ~new_U3888 | ~new_U3889 | ~new_U6413;
  assign n2194 = ~new_U6408 | ~new_U6405 | ~new_U3886 | ~new_U3887 | ~new_U6406;
  assign n2189 = ~new_U3885 | ~new_U6398 | ~new_U3884 | ~new_U6397;
  assign n2184 = ~new_U6390 | ~new_U6391 | ~new_U3883 | ~new_U3882 | ~new_U6389;
  assign n2179 = ~new_U3881 | ~new_U6382 | ~new_U6381 | ~new_U6380;
  assign n2174 = ~new_U3880 | ~new_U6374 | ~new_U6373 | ~new_U6372;
  assign n2169 = ~new_U3879 | ~new_U6366 | ~new_U6365 | ~new_U6364;
  assign n2164 = ~new_U3878 | ~new_U6358 | ~new_U6357 | ~new_U6356;
  assign n2159 = ~new_U6347 | ~new_U6346;
  assign n2154 = ~new_U6343 | ~new_U6344 | ~new_U6345;
  assign n2149 = ~new_U6340 | ~new_U6341 | ~new_U6342;
  assign n2144 = ~new_U6337 | ~new_U6338 | ~new_U6339;
  assign n2139 = ~new_U6334 | ~new_U6335 | ~new_U6336;
  assign n2134 = ~new_U6331 | ~new_U6332 | ~new_U6333;
  assign n2129 = ~new_U6328 | ~new_U6329 | ~new_U6330;
  assign n2124 = ~new_U6325 | ~new_U6326 | ~new_U6327;
  assign n2119 = ~new_U6322 | ~new_U6323 | ~new_U6324;
  assign n2114 = ~new_U6319 | ~new_U6320 | ~new_U6321;
  assign n2109 = ~new_U6316 | ~new_U6317 | ~new_U6318;
  assign n2104 = ~new_U6313 | ~new_U6314 | ~new_U6315;
  assign n2099 = ~new_U6310 | ~new_U6311 | ~new_U6312;
  assign n2094 = ~new_U6307 | ~new_U6308 | ~new_U6309;
  assign n2089 = ~new_U6304 | ~new_U6305 | ~new_U6306;
  assign n2084 = ~new_U6301 | ~new_U6302 | ~new_U6303;
  assign n2079 = ~new_U6298 | ~new_U6299 | ~new_U6300;
  assign n2074 = ~new_U6295 | ~new_U6296 | ~new_U6297;
  assign n2069 = ~new_U6292 | ~new_U6293 | ~new_U6294;
  assign n2064 = ~new_U6289 | ~new_U6290 | ~new_U6291;
  assign n2059 = ~new_U6286 | ~new_U6287 | ~new_U6288;
  assign n2054 = ~new_U6283 | ~new_U6284 | ~new_U6285;
  assign n2049 = ~new_U6280 | ~new_U6281 | ~new_U6282;
  assign n2044 = ~new_U6277 | ~new_U6278 | ~new_U6279;
  assign n2039 = ~new_U6274 | ~new_U6275 | ~new_U6276;
  assign n2034 = ~new_U6271 | ~new_U6272 | ~new_U6273;
  assign n2029 = ~new_U6268 | ~new_U6269 | ~new_U6270;
  assign n2024 = ~new_U6265 | ~new_U6266 | ~new_U6267;
  assign n2019 = ~new_U6262 | ~new_U6263 | ~new_U6264;
  assign n2014 = ~new_U6259 | ~new_U6260 | ~new_U6261;
  assign n2009 = ~new_U6256 | ~new_U6257 | ~new_U6258;
  assign n2004 = ~new_U6255 | ~new_U6254 | ~new_U6253;
  assign n1999 = ~new_U4164 | ~new_U6250;
  assign n1994 = ~new_U6248 | ~new_U6249 | ~new_U6247 | ~new_U6246;
  assign n1989 = ~new_U6244 | ~new_U6245 | ~new_U6243 | ~new_U6242;
  assign n1984 = ~new_U6240 | ~new_U6241 | ~new_U6239 | ~new_U6238;
  assign n1979 = ~new_U6236 | ~new_U6237 | ~new_U6235 | ~new_U6234;
  assign n1974 = ~new_U6232 | ~new_U6233 | ~new_U6231 | ~new_U6230;
  assign n1969 = ~new_U6228 | ~new_U6229 | ~new_U6227 | ~new_U6226;
  assign n1964 = ~new_U6224 | ~new_U6225 | ~new_U6223 | ~new_U6222;
  assign n1959 = ~new_U6220 | ~new_U6221 | ~new_U6219 | ~new_U6218;
  assign n1954 = ~new_U6216 | ~new_U6217 | ~new_U6215 | ~new_U6214;
  assign n1949 = ~new_U6212 | ~new_U6213 | ~new_U6211 | ~new_U6210;
  assign n1944 = ~new_U6208 | ~new_U6209 | ~new_U6207 | ~new_U6206;
  assign n1939 = ~new_U6204 | ~new_U6205 | ~new_U6203 | ~new_U6202;
  assign n1934 = ~new_U6200 | ~new_U6201 | ~new_U6199 | ~new_U6198;
  assign n1929 = ~new_U6196 | ~new_U6197 | ~new_U6195 | ~new_U6194;
  assign n1924 = ~new_U6192 | ~new_U6193 | ~new_U6191 | ~new_U6190;
  assign n1919 = ~new_U6188 | ~new_U6189 | ~new_U6187;
  assign n1914 = ~new_U6185 | ~new_U6186 | ~new_U6184;
  assign n1909 = ~new_U6182 | ~new_U6183 | ~new_U6181;
  assign n1904 = ~new_U6179 | ~new_U6180 | ~new_U6178;
  assign n1899 = ~new_U6176 | ~new_U6177 | ~new_U6175;
  assign n1894 = ~new_U6173 | ~new_U6174 | ~new_U6172;
  assign n1889 = ~new_U6170 | ~new_U6171 | ~new_U6169;
  assign n1884 = ~new_U6167 | ~new_U6168 | ~new_U6166;
  assign n1879 = ~new_U6164 | ~new_U6165 | ~new_U6163;
  assign n1874 = ~new_U6161 | ~new_U6162 | ~new_U6160;
  assign n1869 = ~new_U6158 | ~new_U6159 | ~new_U6157;
  assign n1864 = ~new_U6155 | ~new_U6156 | ~new_U6154;
  assign n1859 = ~new_U6152 | ~new_U6153 | ~new_U6151;
  assign n1854 = ~new_U6149 | ~new_U6150 | ~new_U6148;
  assign n1849 = ~new_U6147 | ~new_U6146 | ~new_U6145;
  assign n1844 = ~new_U6144 | ~new_U6143 | ~new_U6142;
  assign n1840 = DATAO_REG_31_ & new_U6043;
  assign n1836 = ~new_U3870 | ~new_U6134;
  assign n1832 = ~new_U3869 | ~new_U6131;
  assign n1828 = ~new_U3868 | ~new_U6128;
  assign n1824 = ~new_U3867 | ~new_U6125;
  assign n1820 = ~new_U3866 | ~new_U6122;
  assign n1816 = ~new_U3865 | ~new_U6119;
  assign n1812 = ~new_U3864 | ~new_U6116;
  assign n1808 = ~new_U3863 | ~new_U6113;
  assign n1804 = ~new_U3862 | ~new_U6110;
  assign n1800 = ~new_U3861 | ~new_U6107;
  assign n1796 = ~new_U3860 | ~new_U6104;
  assign n1792 = ~new_U3859 | ~new_U6101;
  assign n1788 = ~new_U3858 | ~new_U6098;
  assign n1784 = ~new_U3857 | ~new_U6095;
  assign n1780 = ~new_U3856 | ~new_U6092;
  assign n1776 = ~new_U6091 | ~new_U6090 | ~new_U6089;
  assign n1772 = ~new_U6088 | ~new_U6087 | ~new_U6086;
  assign n1768 = ~new_U6085 | ~new_U6084 | ~new_U6083;
  assign n1764 = ~new_U6082 | ~new_U6081 | ~new_U6080;
  assign n1760 = ~new_U6079 | ~new_U6078 | ~new_U6077;
  assign n1756 = ~new_U6076 | ~new_U6075 | ~new_U6074;
  assign n1752 = ~new_U6073 | ~new_U6072 | ~new_U6071;
  assign n1748 = ~new_U6070 | ~new_U6069 | ~new_U6068;
  assign n1744 = ~new_U6067 | ~new_U6066 | ~new_U6065;
  assign n1740 = ~new_U6064 | ~new_U6063 | ~new_U6062;
  assign n1736 = ~new_U6061 | ~new_U6060 | ~new_U6059;
  assign n1732 = ~new_U6058 | ~new_U6057 | ~new_U6056;
  assign n1728 = ~new_U6055 | ~new_U6054 | ~new_U6053;
  assign n1724 = ~new_U6052 | ~new_U6051 | ~new_U6050;
  assign n1720 = ~new_U6049 | ~new_U6048 | ~new_U6047;
  assign n1716 = ~new_U6046 | ~new_U6045 | ~new_U6044;
  assign n1711 = ~new_U7528 | ~new_U7530;
  assign n1706 = ~new_U7527 | ~new_U7532;
  assign n1701 = ~new_U7526 | ~new_U7534;
  assign n1696 = ~new_U7525 | ~new_U7536;
  assign n1691 = ~new_U7524 | ~new_U7538;
  assign n1686 = ~new_U7523 | ~new_U7540;
  assign n1681 = ~new_U7522 | ~new_U7542;
  assign n1676 = ~new_U7521 | ~new_U7544;
  assign n1671 = ~new_U7520 | ~new_U7546;
  assign n1666 = ~new_U7519 | ~new_U7548;
  assign n1661 = ~new_U7518 | ~new_U7550;
  assign n1656 = ~new_U7517 | ~new_U7552;
  assign n1651 = ~new_U7516 | ~new_U7554;
  assign n1646 = ~new_U7515 | ~new_U7556;
  assign n1641 = ~new_U7514 | ~new_U7558;
  assign n1636 = ~new_U7513 | ~new_U7560;
  assign n1631 = ~new_U7512 | ~new_U7562;
  assign n1626 = ~new_U7511 | ~new_U7564;
  assign n1621 = ~new_U7510 | ~new_U7566;
  assign n1616 = ~new_U7509 | ~new_U7568;
  assign n1611 = ~new_U7508 | ~new_U7570;
  assign n1606 = ~new_U7507 | ~new_U7572;
  assign n1601 = ~new_U7506 | ~new_U7574;
  assign n1596 = ~new_U7505 | ~new_U7576;
  assign n1591 = ~new_U7504 | ~new_U7578;
  assign n1586 = ~new_U7503 | ~new_U7580;
  assign n1581 = ~new_U7502 | ~new_U7582;
  assign n1576 = ~new_U7501 | ~new_U7584;
  assign n1571 = ~new_U7500 | ~new_U7586;
  assign n1566 = ~new_U7499 | ~new_U7588;
  assign n1561 = ~new_U7498 | ~new_U7590;
  assign n1556 = ~new_U5945 | ~new_U5943 | ~new_U5946 | ~new_U5944 | ~new_U5942;
  assign n1551 = ~new_U5940 | ~new_U5938 | ~new_U5941 | ~new_U5939 | ~new_U5937;
  assign n1546 = ~new_U5935 | ~new_U5933 | ~new_U5936 | ~new_U5934 | ~new_U5932;
  assign n1541 = ~new_U5930 | ~new_U5928 | ~new_U5931 | ~new_U5929 | ~new_U5927;
  assign n1536 = ~new_U5925 | ~new_U5923 | ~new_U5926 | ~new_U5924 | ~new_U5922;
  assign n1531 = ~new_U5920 | ~new_U5918 | ~new_U5921 | ~new_U5919 | ~new_U5917;
  assign n1526 = ~new_U5915 | ~new_U5913 | ~new_U5916 | ~new_U5914 | ~new_U5912;
  assign n1521 = ~new_U5910 | ~new_U5908 | ~new_U5911 | ~new_U5909 | ~new_U5907;
  assign n1516 = ~new_U5905 | ~new_U5903 | ~new_U5906 | ~new_U5904 | ~new_U5902;
  assign n1511 = ~new_U5900 | ~new_U5898 | ~new_U5901 | ~new_U5899 | ~new_U5897;
  assign n1506 = ~new_U5895 | ~new_U5893 | ~new_U5896 | ~new_U5894 | ~new_U5892;
  assign n1501 = ~new_U5890 | ~new_U5888 | ~new_U5891 | ~new_U5889 | ~new_U5887;
  assign n1496 = ~new_U5885 | ~new_U5883 | ~new_U5886 | ~new_U5884 | ~new_U5882;
  assign n1491 = ~new_U5880 | ~new_U5878 | ~new_U5881 | ~new_U5879 | ~new_U5877;
  assign n1486 = ~new_U5875 | ~new_U5873 | ~new_U5876 | ~new_U5874 | ~new_U5872;
  assign n1481 = ~new_U5870 | ~new_U5868 | ~new_U5871 | ~new_U5869 | ~new_U5867;
  assign n1476 = ~new_U5865 | ~new_U5863 | ~new_U5866 | ~new_U5864 | ~new_U5862;
  assign n1471 = ~new_U5860 | ~new_U5858 | ~new_U5861 | ~new_U5859 | ~new_U5857;
  assign n1466 = ~new_U5855 | ~new_U5853 | ~new_U5856 | ~new_U5854 | ~new_U5852;
  assign n1461 = ~new_U5850 | ~new_U5848 | ~new_U5851 | ~new_U5849 | ~new_U5847;
  assign n1456 = ~new_U5845 | ~new_U5843 | ~new_U5846 | ~new_U5844 | ~new_U5842;
  assign n1451 = ~new_U5840 | ~new_U5838 | ~new_U5841 | ~new_U5839 | ~new_U5837;
  assign n1446 = ~new_U5835 | ~new_U5833 | ~new_U5836 | ~new_U5834 | ~new_U5832;
  assign n1441 = ~new_U5830 | ~new_U5828 | ~new_U5831 | ~new_U5829 | ~new_U5827;
  assign n1436 = ~new_U5825 | ~new_U5826 | ~new_U5823 | ~new_U5824 | ~new_U5822;
  assign n1431 = ~new_U5820 | ~new_U5821 | ~new_U5818 | ~new_U5819 | ~new_U5817;
  assign n1426 = ~new_U5815 | ~new_U5816 | ~new_U5813 | ~new_U5814 | ~new_U5812;
  assign n1421 = ~new_U5810 | ~new_U5811 | ~new_U5808 | ~new_U5809 | ~new_U5807;
  assign n1416 = ~new_U5805 | ~new_U5806 | ~new_U5803 | ~new_U5804 | ~new_U5802;
  assign n1411 = ~new_U5800 | ~new_U5801 | ~new_U5798 | ~new_U5799 | ~new_U5797;
  assign n1406 = ~new_U5795 | ~new_U5796 | ~new_U5794 | ~new_U5793 | ~new_U5792;
  assign n1401 = ~new_U5790 | ~new_U5791 | ~new_U5789 | ~new_U5788 | ~new_U5787;
  assign n1396 = ~new_U5777 | ~new_U5775 | ~new_U3849 | ~new_U3847;
  assign n1391 = ~new_U5770 | ~new_U5768 | ~new_U3846 | ~new_U3844;
  assign n1386 = ~new_U5763 | ~new_U5761 | ~new_U3843 | ~new_U3841;
  assign n1381 = ~new_U5756 | ~new_U5754 | ~new_U3840 | ~new_U3838;
  assign n1376 = ~new_U5749 | ~new_U5747 | ~new_U3837 | ~new_U3835;
  assign n1371 = ~new_U5742 | ~new_U5740 | ~new_U3834 | ~new_U3832;
  assign n1366 = ~new_U5735 | ~new_U5733 | ~new_U3831 | ~new_U3829;
  assign n1361 = ~new_U5728 | ~new_U5726 | ~new_U3828 | ~new_U3826;
  assign n1356 = ~new_U5721 | ~new_U5719 | ~new_U3825 | ~new_U3823;
  assign n1351 = ~new_U5714 | ~new_U5712 | ~new_U3822 | ~new_U3820;
  assign n1346 = ~new_U5707 | ~new_U5705 | ~new_U3819 | ~new_U3817;
  assign n1341 = ~new_U5700 | ~new_U5698 | ~new_U3816 | ~new_U3814;
  assign n1336 = ~new_U5693 | ~new_U5691 | ~new_U3813 | ~new_U3811;
  assign n1331 = ~new_U5686 | ~new_U5684 | ~new_U3810 | ~new_U3808;
  assign n1326 = ~new_U5679 | ~new_U5677 | ~new_U3807 | ~new_U3805;
  assign n1321 = ~new_U5672 | ~new_U5670 | ~new_U3804 | ~new_U3802;
  assign n1316 = ~new_U5665 | ~new_U5663 | ~new_U3801 | ~new_U3799;
  assign n1311 = ~new_U5658 | ~new_U5656 | ~new_U3798 | ~new_U3796;
  assign n1306 = ~new_U5651 | ~new_U5649 | ~new_U3795 | ~new_U3793;
  assign n1301 = ~new_U5644 | ~new_U3790 | ~new_U3792;
  assign n1296 = ~new_U5637 | ~new_U3787 | ~new_U3789;
  assign n1291 = ~new_U5630 | ~new_U3784 | ~new_U3786;
  assign n1286 = ~new_U5623 | ~new_U3781 | ~new_U3783;
  assign n1281 = ~new_U5616 | ~new_U3778 | ~new_U3780;
  assign n1276 = ~new_U5609 | ~new_U3775 | ~new_U3777;
  assign n1271 = ~new_U5602 | ~new_U3772 | ~new_U3774;
  assign n1266 = ~new_U5595 | ~new_U3769 | ~new_U3771;
  assign n1261 = ~new_U5588 | ~new_U3766 | ~new_U3768;
  assign n1256 = ~new_U3763 | ~new_U3764;
  assign n1251 = ~new_U3762 | ~new_U3760 | ~new_U3759;
  assign n1246 = ~new_U3758 | ~new_U3756 | ~new_U3755;
  assign n1241 = ~new_U3754 | ~new_U3752 | ~new_U3751;
  assign n1216 = INSTQUEUEWR_ADDR_REG_4_ & new_U5525;
  assign n1186 = ~new_U3718 | ~new_U5448 | ~new_U5447;
  assign n1181 = ~new_U3717 | ~new_U5443 | ~new_U5442;
  assign n1176 = ~new_U3716 | ~new_U5438 | ~new_U5437;
  assign n1171 = ~new_U3715 | ~new_U5433 | ~new_U5432;
  assign n1166 = ~new_U3714 | ~new_U7600 | ~new_U5428;
  assign n1161 = ~new_U3713 | ~new_U5424 | ~new_U5423;
  assign n1156 = ~new_U3712 | ~new_U5419 | ~new_U5418;
  assign n1151 = ~new_U3711 | ~new_U5414 | ~new_U5413;
  assign n1146 = ~new_U3709 | ~new_U5392 | ~new_U5391;
  assign n1141 = ~new_U3708 | ~new_U5387 | ~new_U5386;
  assign n1136 = ~new_U3707 | ~new_U5382 | ~new_U5381;
  assign n1131 = ~new_U3706 | ~new_U5377 | ~new_U5376;
  assign n1126 = ~new_U3705 | ~new_U5372 | ~new_U5371;
  assign n1121 = ~new_U3704 | ~new_U5367 | ~new_U5366;
  assign n1116 = ~new_U3703 | ~new_U5362 | ~new_U5361;
  assign n1111 = ~new_U3702 | ~new_U5357 | ~new_U5356;
  assign n1106 = ~new_U3700 | ~new_U5334 | ~new_U5333;
  assign n1101 = ~new_U3699 | ~new_U5329 | ~new_U5328;
  assign n1096 = ~new_U3698 | ~new_U5324 | ~new_U5323;
  assign n1091 = ~new_U3697 | ~new_U5319 | ~new_U5318;
  assign n1086 = ~new_U3696 | ~new_U5314 | ~new_U5313;
  assign n1081 = ~new_U3695 | ~new_U5309 | ~new_U5308;
  assign n1076 = ~new_U3694 | ~new_U5304 | ~new_U5303;
  assign n1071 = ~new_U3693 | ~new_U5299 | ~new_U5298;
  assign n1066 = ~new_U3691 | ~new_U5277 | ~new_U5276;
  assign n1061 = ~new_U3690 | ~new_U5272 | ~new_U5271;
  assign n1056 = ~new_U3689 | ~new_U5267 | ~new_U5266;
  assign n1051 = ~new_U3688 | ~new_U5262 | ~new_U5261;
  assign n1046 = ~new_U3687 | ~new_U5257 | ~new_U5256;
  assign n1041 = ~new_U3686 | ~new_U5252 | ~new_U5251;
  assign n1036 = ~new_U3685 | ~new_U5247 | ~new_U5246;
  assign n1031 = ~new_U3684 | ~new_U5242 | ~new_U5241;
  assign n1026 = ~new_U3682 | ~new_U5219 | ~new_U5218;
  assign n1021 = ~new_U3681 | ~new_U5214 | ~new_U5213;
  assign n1016 = ~new_U3680 | ~new_U5209 | ~new_U5208;
  assign n1011 = ~new_U3679 | ~new_U5204 | ~new_U5203;
  assign n1006 = ~new_U3678 | ~new_U5199 | ~new_U5198;
  assign n1001 = ~new_U3677 | ~new_U5194 | ~new_U5193;
  assign n996 = ~new_U3676 | ~new_U5189 | ~new_U5188;
  assign n991 = ~new_U3675 | ~new_U5184 | ~new_U5183;
  assign n986 = ~new_U3673 | ~new_U5162 | ~new_U5161;
  assign n981 = ~new_U3672 | ~new_U5157 | ~new_U5156;
  assign n976 = ~new_U3671 | ~new_U5152 | ~new_U5151;
  assign n971 = ~new_U3670 | ~new_U5147 | ~new_U5146;
  assign n966 = ~new_U3669 | ~new_U5142 | ~new_U5141;
  assign n961 = ~new_U3668 | ~new_U5137 | ~new_U5136;
  assign n956 = ~new_U3667 | ~new_U5132 | ~new_U5131;
  assign n951 = ~new_U3666 | ~new_U5127 | ~new_U5126;
  assign n946 = ~new_U3664 | ~new_U5104 | ~new_U5103;
  assign n941 = ~new_U3663 | ~new_U5099 | ~new_U5098;
  assign n936 = ~new_U3662 | ~new_U5094 | ~new_U5093;
  assign n931 = ~new_U3661 | ~new_U5089 | ~new_U5088;
  assign n926 = ~new_U3660 | ~new_U5084 | ~new_U5083;
  assign n921 = ~new_U3659 | ~new_U5079 | ~new_U5078;
  assign n916 = ~new_U3658 | ~new_U5074 | ~new_U5073;
  assign n911 = ~new_U3657 | ~new_U5069 | ~new_U5068;
  assign n906 = ~new_U3655 | ~new_U5047 | ~new_U5046;
  assign n901 = ~new_U3654 | ~new_U5042 | ~new_U5041;
  assign n896 = ~new_U3653 | ~new_U5037 | ~new_U5036;
  assign n891 = ~new_U3652 | ~new_U5032 | ~new_U5031;
  assign n886 = ~new_U3651 | ~new_U5027 | ~new_U5026;
  assign n881 = ~new_U3650 | ~new_U5022 | ~new_U5021;
  assign n876 = ~new_U3649 | ~new_U5017 | ~new_U5016;
  assign n871 = ~new_U3648 | ~new_U5012 | ~new_U5011;
  assign n866 = ~new_U3646 | ~new_U4991 | ~new_U4990;
  assign n861 = ~new_U3645 | ~new_U4986 | ~new_U4985;
  assign n856 = ~new_U3644 | ~new_U4981 | ~new_U4980;
  assign n851 = ~new_U3643 | ~new_U4976 | ~new_U4975;
  assign n846 = ~new_U3642 | ~new_U4971 | ~new_U4970;
  assign n841 = ~new_U3641 | ~new_U4966 | ~new_U4965;
  assign n836 = ~new_U3640 | ~new_U4961 | ~new_U4960;
  assign n831 = ~new_U3639 | ~new_U4956 | ~new_U4955;
  assign n826 = ~new_U3637 | ~new_U4934 | ~new_U4933;
  assign n821 = ~new_U3636 | ~new_U4929 | ~new_U4928;
  assign n816 = ~new_U3635 | ~new_U4924 | ~new_U4923;
  assign n811 = ~new_U3634 | ~new_U4919 | ~new_U4918;
  assign n806 = ~new_U3633 | ~new_U4914 | ~new_U4913;
  assign n801 = ~new_U3632 | ~new_U4909 | ~new_U4908;
  assign n796 = ~new_U3631 | ~new_U4904 | ~new_U4903;
  assign n791 = ~new_U3630 | ~new_U4899 | ~new_U4898;
  assign n786 = ~new_U3628 | ~new_U4876 | ~new_U4875;
  assign n781 = ~new_U3627 | ~new_U4871 | ~new_U4870;
  assign n776 = ~new_U3626 | ~new_U4866 | ~new_U4865;
  assign n771 = ~new_U3625 | ~new_U4861 | ~new_U4860;
  assign n766 = ~new_U3624 | ~new_U4856 | ~new_U4855;
  assign n761 = ~new_U3623 | ~new_U4851 | ~new_U4850;
  assign n756 = ~new_U3622 | ~new_U4846 | ~new_U4845;
  assign n751 = ~new_U3621 | ~new_U4841 | ~new_U4840;
  assign n746 = ~new_U3619 | ~new_U4819 | ~new_U4818;
  assign n741 = ~new_U3618 | ~new_U4814 | ~new_U4813;
  assign n736 = ~new_U3617 | ~new_U4809 | ~new_U4808;
  assign n731 = ~new_U3616 | ~new_U4804 | ~new_U4803;
  assign n726 = ~new_U3615 | ~new_U4799 | ~new_U4798;
  assign n721 = ~new_U3614 | ~new_U4794 | ~new_U4793;
  assign n716 = ~new_U3613 | ~new_U4789 | ~new_U4788;
  assign n711 = ~new_U3612 | ~new_U4784 | ~new_U4783;
  assign n706 = ~new_U3610 | ~new_U4761 | ~new_U4760;
  assign n701 = ~new_U3609 | ~new_U4756 | ~new_U4755;
  assign n696 = ~new_U3608 | ~new_U4751 | ~new_U4750;
  assign n691 = ~new_U3607 | ~new_U4746 | ~new_U4745;
  assign n686 = ~new_U3606 | ~new_U4741 | ~new_U4740;
  assign n681 = ~new_U3605 | ~new_U4736 | ~new_U4735;
  assign n676 = ~new_U3604 | ~new_U4731 | ~new_U4730;
  assign n671 = ~new_U3603 | ~new_U4726 | ~new_U4725;
  assign n666 = ~new_U3601 | ~new_U4704 | ~new_U4703;
  assign n661 = ~new_U3600 | ~new_U4699 | ~new_U4698;
  assign n656 = ~new_U3599 | ~new_U4694 | ~new_U4693;
  assign n651 = ~new_U3598 | ~new_U4689 | ~new_U4688;
  assign n646 = ~new_U3597 | ~new_U4684 | ~new_U4683;
  assign n641 = ~new_U3596 | ~new_U4679 | ~new_U4678;
  assign n636 = ~new_U3595 | ~new_U4674 | ~new_U4673;
  assign n631 = ~new_U3594 | ~new_U4669 | ~new_U4668;
  assign n626 = ~new_U3592 | ~new_U4645 | ~new_U4644;
  assign n621 = ~new_U3591 | ~new_U4640 | ~new_U4639;
  assign n616 = ~new_U3590 | ~new_U4635 | ~new_U4634;
  assign n611 = ~new_U3589 | ~new_U4630 | ~new_U4629;
  assign n606 = ~new_U3588 | ~new_U4625 | ~new_U4624;
  assign n601 = ~new_U3587 | ~new_U4620 | ~new_U4619;
  assign n596 = ~new_U3586 | ~new_U4615 | ~new_U4614;
  assign n591 = ~new_U3585 | ~new_U4610 | ~new_U4609;
  assign n586 = ~new_U3583 | ~new_U4587 | ~new_U4586;
  assign n581 = ~new_U3582 | ~new_U4582 | ~new_U4581;
  assign n576 = ~new_U3581 | ~new_U4577 | ~new_U4576;
  assign n571 = ~new_U3580 | ~new_U4572 | ~new_U4571;
  assign n566 = ~new_U3579 | ~new_U4567 | ~new_U4566;
  assign n561 = ~new_U3578 | ~new_U4562 | ~new_U4561;
  assign n556 = ~new_U3577 | ~new_U4557 | ~new_U4556;
  assign n551 = ~new_U3576 | ~new_U4552 | ~new_U4551;
  assign n546 = ~new_U3574 | ~new_U7678 | ~new_U7677;
  assign n541 = ~new_U4232 | ~new_U4506 | ~new_U4508 | ~new_U4507;
  assign n536 = ~new_U3570 | ~new_U4504;
  assign n526 = DATAWIDTH_REG_31_ & new_U7638;
  assign n521 = DATAWIDTH_REG_30_ & new_U7638;
  assign n516 = DATAWIDTH_REG_29_ & new_U7638;
  assign n511 = DATAWIDTH_REG_28_ & new_U7638;
  assign n506 = DATAWIDTH_REG_27_ & new_U7638;
  assign n501 = DATAWIDTH_REG_26_ & new_U7638;
  assign n496 = DATAWIDTH_REG_25_ & new_U7638;
  assign n491 = DATAWIDTH_REG_24_ & new_U7638;
  assign n486 = DATAWIDTH_REG_23_ & new_U7638;
  assign n481 = DATAWIDTH_REG_22_ & new_U7638;
  assign n476 = DATAWIDTH_REG_21_ & new_U7638;
  assign n471 = DATAWIDTH_REG_20_ & new_U7638;
  assign n466 = DATAWIDTH_REG_19_ & new_U7638;
  assign n461 = DATAWIDTH_REG_18_ & new_U7638;
  assign n456 = DATAWIDTH_REG_17_ & new_U7638;
  assign n451 = DATAWIDTH_REG_16_ & new_U7638;
  assign n446 = DATAWIDTH_REG_15_ & new_U7638;
  assign n441 = DATAWIDTH_REG_14_ & new_U7638;
  assign n436 = DATAWIDTH_REG_13_ & new_U7638;
  assign n431 = DATAWIDTH_REG_12_ & new_U7638;
  assign n426 = DATAWIDTH_REG_11_ & new_U7638;
  assign n421 = DATAWIDTH_REG_10_ & new_U7638;
  assign n416 = DATAWIDTH_REG_9_ & new_U7638;
  assign n411 = DATAWIDTH_REG_8_ & new_U7638;
  assign n406 = DATAWIDTH_REG_7_ & new_U7638;
  assign n401 = DATAWIDTH_REG_6_ & new_U7638;
  assign n396 = DATAWIDTH_REG_5_ & new_U7638;
  assign n391 = DATAWIDTH_REG_4_ & new_U7638;
  assign n386 = DATAWIDTH_REG_3_ & new_U7638;
  assign n381 = DATAWIDTH_REG_2_ & new_U7638;
  assign n366 = ~new_U4363 | ~new_U7635 | ~new_U7634;
  assign n361 = ~new_U3483 | ~new_U7633 | ~new_U7632;
  assign n356 = ~new_U3482 | ~new_U4357;
  assign n352 = ~new_U4344 | ~new_U4343 | ~new_U4342;
  assign n348 = ~new_U4341 | ~new_U4340 | ~new_U4339;
  assign n344 = ~new_U4338 | ~new_U4337 | ~new_U4336;
  assign n340 = ~new_U4335 | ~new_U4334 | ~new_U4333;
  assign n336 = ~new_U4332 | ~new_U4331 | ~new_U4330;
  assign n332 = ~new_U4329 | ~new_U4328 | ~new_U4327;
  assign n328 = ~new_U4326 | ~new_U4325 | ~new_U4324;
  assign n324 = ~new_U4323 | ~new_U4322 | ~new_U4321;
  assign n320 = ~new_U4320 | ~new_U4319 | ~new_U4318;
  assign n316 = ~new_U4317 | ~new_U4316 | ~new_U4315;
  assign n312 = ~new_U4314 | ~new_U4313 | ~new_U4312;
  assign n308 = ~new_U4311 | ~new_U4310 | ~new_U4309;
  assign n304 = ~new_U4308 | ~new_U4307 | ~new_U4306;
  assign n300 = ~new_U4305 | ~new_U4304 | ~new_U4303;
  assign n296 = ~new_U4302 | ~new_U4301 | ~new_U4300;
  assign n292 = ~new_U4299 | ~new_U4298 | ~new_U4297;
  assign n288 = ~new_U4296 | ~new_U4295 | ~new_U4294;
  assign n284 = ~new_U4293 | ~new_U4292 | ~new_U4291;
  assign n280 = ~new_U4290 | ~new_U4289 | ~new_U4288;
  assign n276 = ~new_U4287 | ~new_U4286 | ~new_U4285;
  assign n272 = ~new_U4284 | ~new_U4283 | ~new_U4282;
  assign n268 = ~new_U4281 | ~new_U4280 | ~new_U4279;
  assign n264 = ~new_U4278 | ~new_U4277 | ~new_U4276;
  assign n260 = ~new_U4275 | ~new_U4274 | ~new_U4273;
  assign n256 = ~new_U4272 | ~new_U4271 | ~new_U4270;
  assign n252 = ~new_U4269 | ~new_U4268 | ~new_U4267;
  assign n248 = ~new_U4266 | ~new_U4265 | ~new_U4264;
  assign n244 = ~new_U4263 | ~new_U4262 | ~new_U4261;
  assign n240 = ~new_U4260 | ~new_U4259 | ~new_U4258;
  assign n236 = ~new_U4257 | ~new_U4256 | ~new_U4255;
  assign new_U3214 = ~new_U3986 | ~new_U3987 | ~new_U3989 | ~new_U3988;
  assign new_U3215 = ~new_U3982 | ~new_U3983 | ~new_U3985 | ~new_U3984;
  assign new_U3216 = ~new_U3978 | ~new_U3979 | ~new_U3981 | ~new_U3980;
  assign new_U3217 = ~new_U3974 | ~new_U3975 | ~new_U3977 | ~new_U3976;
  assign new_U3218 = ~new_U3970 | ~new_U3971 | ~new_U3973 | ~new_U3972;
  assign new_U3219 = ~new_U3966 | ~new_U3967 | ~new_U3969 | ~new_U3968;
  assign new_U3220 = ~new_U3962 | ~new_U3963 | ~new_U3965 | ~new_U3964;
  assign new_U3221 = ~new_U3958 | ~new_U3959 | ~new_U3961 | ~new_U3960;
  assign new_U3222 = ~new_U3316 | ~new_U3310;
  assign new_U3223 = ~new_U2432 | ~new_U3222;
  assign new_U3224 = ~new_U2432 | ~new_U4531;
  assign new_U3225 = ~new_U2434 | ~new_U3222;
  assign new_U3226 = ~new_U2434 | ~new_U4531;
  assign new_U3227 = ~new_U2433 | ~new_U3222;
  assign new_U3228 = ~new_U2433 | ~new_U4531;
  assign new_U3229 = ~new_U2435 | ~new_U3222;
  assign new_U3230 = ~new_U2435 | ~new_U4531;
  assign new_U3231 = ~new_U5451 | ~new_U3378 | ~new_U3381;
  assign new_U3232 = ~new_U7074 | ~new_U5452;
  assign new_U3233 = ~new_U4144 | ~new_U4146 | ~new_U7780 | ~new_U7779;
  assign new_U3234 = ~REQUESTPENDING_REG;
  assign new_U3235 = ~STATE_REG_1_;
  assign new_U3236 = ~STATE_REG_1_ | ~new_U3245;
  assign new_U3237 = ~new_U4209 | ~new_U3238;
  assign new_U3238 = ~STATE_REG_2_;
  assign new_U3239 = ~STATE_REG_2_ | ~new_U4209;
  assign new_U3240 = ~REIP_REG_1_;
  assign new_U3241 = ~STATE_REG_1_ | ~new_U3238;
  assign new_U3242 = STATE_REG_1_ | STATE_REG_2_;
  assign new_U3243 = ~HOLD;
  assign new_U3244 = ~READY_N;
  assign new_U3245 = ~STATE_REG_0_;
  assign new_U3246 = ~STATE_REG_0_ | ~new_U3247;
  assign new_U3247 = ~REQUESTPENDING_REG | ~new_U3243;
  assign new_U3248 = HOLD | REQUESTPENDING_REG;
  assign new_U3249 = ~STATE2_REG_1_;
  assign new_U3250 = ~STATE2_REG_2_;
  assign new_U3251 = ~INSTQUEUERD_ADDR_REG_2_;
  assign new_U3252 = ~INSTQUEUERD_ADDR_REG_1_;
  assign new_U3253 = ~INSTQUEUERD_ADDR_REG_0_;
  assign new_U3254 = ~new_U3257 | ~INSTQUEUERD_ADDR_REG_2_ | ~INSTQUEUERD_ADDR_REG_0_ | ~INSTQUEUERD_ADDR_REG_1_;
  assign new_U3255 = INSTQUEUERD_ADDR_REG_2_ | INSTQUEUERD_ADDR_REG_0_ | INSTQUEUERD_ADDR_REG_1_;
  assign new_U3256 = INSTQUEUERD_ADDR_REG_1_ | INSTQUEUERD_ADDR_REG_0_;
  assign new_U3257 = ~INSTQUEUERD_ADDR_REG_3_;
  assign new_U3258 = ~new_U3552 | ~new_U3553 | ~new_U3555 | ~new_U3554;
  assign new_U3259 = ~new_U4484 | ~new_U3245;
  assign new_U3260 = ~new_R2167_U17;
  assign new_U3261 = ~INSTQUEUERD_ADDR_REG_2_ | ~new_U3257;
  assign new_U3262 = ~INSTQUEUERD_ADDR_REG_0_ | ~INSTQUEUERD_ADDR_REG_1_;
  assign new_U3263 = ~new_U3504 | ~new_U3505 | ~new_U3507 | ~new_U3506;
  assign new_U3264 = ~new_U3524 | ~new_U3525 | ~new_U3526 | ~new_U3527 | ~new_U4158;
  assign new_U3265 = ~new_U3542 | ~new_U3543 | ~new_U3545 | ~new_U3544;
  assign new_U3266 = ~new_U3547 | ~new_U3546;
  assign new_U3267 = STATEBS16_REG | READY_N;
  assign new_U3268 = ~new_R2167_U17 | ~new_U4485;
  assign new_U3269 = ~new_U4465 | ~new_U3271;
  assign new_U3270 = ~new_U3496 | ~new_U3497 | ~new_U3499 | ~new_U3498;
  assign new_U3271 = ~new_U3548 | ~new_U3549 | ~new_U3551 | ~new_U3550;
  assign new_U3272 = ~new_U2473 | ~new_U4489;
  assign new_U3273 = ~new_U2389 | ~new_U3270;
  assign new_U3274 = ~new_U4482 | ~new_U4465;
  assign new_U3275 = ~new_U4237 | ~new_U2447;
  assign new_U3276 = ~new_U3265 | ~new_U4161 | ~new_U4448 | ~new_U3378;
  assign new_U3277 = ~new_U3258 | ~new_U3270;
  assign new_U3278 = ~new_U4178 | ~new_U3271;
  assign new_U3279 = ~new_U4244 | ~new_U2431;
  assign new_U3280 = ~new_LT_563_U6 | ~new_U4213 | ~new_U7614 | ~new_U4166 | ~new_U4497;
  assign new_U3281 = ~STATE2_REG_0_;
  assign new_U3282 = ~STATE2_REG_0_ | ~new_U7592;
  assign new_U3283 = ~STATE2_REG_3_;
  assign new_U3284 = ~STATE2_REG_2_ | ~new_U3249;
  assign new_U3285 = STATE2_REG_2_ | STATE2_REG_1_;
  assign new_U3286 = ~STATE2_REG_3_ | ~new_R2167_U17;
  assign new_U3287 = ~new_U4535 | ~new_U3281;
  assign new_U3288 = ~INSTQUEUEWR_ADDR_REG_0_;
  assign new_U3289 = ~INSTQUEUEWR_ADDR_REG_1_;
  assign new_U3290 = ~INSTQUEUEWR_ADDR_REG_3_;
  assign new_U3291 = ~INSTQUEUEWR_ADDR_REG_2_;
  assign new_U3292 = ~INSTQUEUEWR_ADDR_REG_1_ | ~INSTQUEUEWR_ADDR_REG_0_;
  assign new_U3293 = ~new_U4521 | ~new_U2478;
  assign new_U3294 = STATE2_REG_2_ | STATE2_REG_3_;
  assign new_U3295 = ~STATEBS16_REG;
  assign new_U3296 = ~new_R2144_U43;
  assign new_U3297 = ~new_R2144_U50;
  assign new_U3298 = ~new_R2144_U49;
  assign new_U3299 = ~new_R2144_U8;
  assign new_U3300 = ~new_R2144_U50 | ~new_R2144_U43;
  assign new_U3301 = ~new_U3319 | ~new_U3296;
  assign new_U3302 = ~new_U4515 | ~new_U2475;
  assign new_U3303 = ~new_R2182_U25;
  assign new_U3304 = ~new_R2182_U42;
  assign new_U3305 = ~new_R2182_U34;
  assign new_U3306 = ~new_R2182_U33;
  assign new_U3307 = ~new_U4197 | ~new_U3295;
  assign new_U3308 = ~new_U3293 | ~new_U4523;
  assign new_U3309 = ~new_U3293 | ~new_U4532;
  assign new_U3310 = ~INSTQUEUEWR_ADDR_REG_1_ | ~new_U3288;
  assign new_U3311 = ~new_U4530 | ~new_U2478;
  assign new_U3312 = ~new_R2144_U50 | ~new_U3296;
  assign new_U3313 = ~new_R2144_U43 | ~new_U3319;
  assign new_U3314 = ~new_U4588 | ~new_U2475;
  assign new_U3315 = ~new_U3311 | ~new_U4591;
  assign new_U3316 = ~INSTQUEUEWR_ADDR_REG_0_ | ~new_U3289;
  assign new_U3317 = ~new_U4529 | ~new_U2478;
  assign new_U3318 = ~new_R2144_U43 | ~new_U3297;
  assign new_U3319 = ~new_U3312 | ~new_U3318;
  assign new_U3320 = ~new_U4514 | ~new_U3296;
  assign new_U3321 = ~new_U4646 | ~new_U2475;
  assign new_U3322 = ~new_U3317 | ~new_U4649;
  assign new_U3323 = ~new_U3317 | ~new_U4651;
  assign new_U3324 = ~new_U2488 | ~new_U2478;
  assign new_U3325 = ~new_U2485 | ~new_U2475;
  assign new_U3326 = ~new_U3324 | ~new_U4707;
  assign new_U3327 = ~INSTQUEUEWR_ADDR_REG_3_ | ~new_U3291;
  assign new_U3328 = ~new_U4526 | ~new_U4521;
  assign new_U3329 = ~new_R2144_U8 | ~new_U3298;
  assign new_U3330 = ~new_U2490 | ~new_U4515;
  assign new_U3331 = ~new_U3328 | ~new_U4764;
  assign new_U3332 = ~new_U3328 | ~new_U4766;
  assign new_U3333 = ~new_U4526 | ~new_U4530;
  assign new_U3334 = ~new_U2490 | ~new_U4588;
  assign new_U3335 = ~new_U3333 | ~new_U4822;
  assign new_U3336 = ~new_U4526 | ~new_U4529;
  assign new_U3337 = ~new_U2490 | ~new_U4646;
  assign new_U3338 = ~new_U3336 | ~new_U4879;
  assign new_U3339 = ~new_U3336 | ~new_U4881;
  assign new_U3340 = ~new_U4526 | ~new_U2488;
  assign new_U3341 = ~new_U2490 | ~new_U2485;
  assign new_U3342 = ~new_U3340 | ~new_U4937;
  assign new_U3343 = ~new_U2479 | ~new_U4521;
  assign new_U3344 = ~new_U2474 | ~new_U4516;
  assign new_U3345 = ~new_U3344 | ~new_U3329 | ~new_U4518;
  assign new_U3346 = ~new_U2499 | ~new_U4515;
  assign new_U3347 = ~new_U3343 | ~new_U3327 | ~new_U4527;
  assign new_U3348 = ~new_U3343 | ~new_U4993;
  assign new_U3349 = ~new_U3343 | ~new_U4995;
  assign new_U3350 = ~new_U4530 | ~new_U2479;
  assign new_U3351 = ~new_U2499 | ~new_U4588;
  assign new_U3352 = ~new_U3350 | ~new_U5050;
  assign new_U3353 = ~new_U4529 | ~new_U2479;
  assign new_U3354 = ~new_U2499 | ~new_U4646;
  assign new_U3355 = ~new_U3353 | ~new_U5107;
  assign new_U3356 = ~new_U3353 | ~new_U5109;
  assign new_U3357 = ~new_U2488 | ~new_U2479;
  assign new_U3358 = ~new_U2499 | ~new_U2485;
  assign new_U3359 = ~new_U3357 | ~new_U5165;
  assign new_U3360 = ~new_U2510 | ~new_U4521;
  assign new_U3361 = ~new_U2507 | ~new_U4515;
  assign new_U3362 = ~new_U3360 | ~new_U5222;
  assign new_U3363 = ~new_U3360 | ~new_U5224;
  assign new_U3364 = ~new_U2510 | ~new_U4530;
  assign new_U3365 = ~new_U2507 | ~new_U4588;
  assign new_U3366 = ~new_U3364 | ~new_U5280;
  assign new_U3367 = ~new_U2510 | ~new_U4529;
  assign new_U3368 = ~new_U2507 | ~new_U4646;
  assign new_U3369 = ~new_U3367 | ~new_U5337;
  assign new_U3370 = ~new_U3367 | ~new_U5339;
  assign new_U3371 = ~new_U2510 | ~new_U2488;
  assign new_U3372 = ~new_U2507 | ~new_U2485;
  assign new_U3373 = ~new_U3371 | ~new_U5395;
  assign new_U3374 = ~FLUSH_REG;
  assign new_U3375 = ~new_GTE_485_U6;
  assign new_U3376 = ~new_U3271 | ~new_U3265;
  assign new_U3377 = ~new_U3271 | ~new_U3258;
  assign new_U3378 = ~new_U3500 | ~new_U3501 | ~new_U3503 | ~new_U3502;
  assign new_U3379 = ~new_U7616 | ~new_U5478 | ~new_U5477;
  assign new_U3380 = ~new_U4387 | ~new_U3271;
  assign new_U3381 = ~new_U2605 | ~new_U3264;
  assign new_U3382 = ~new_U4482 | ~new_U4387 | ~new_U7482;
  assign new_U3383 = ~new_U3729 | ~new_U4235;
  assign new_U3384 = ~new_U4387 | ~new_U4482 | ~new_U2605 | ~new_U7482 | ~new_U4465;
  assign new_U3385 = ~new_U4388 | ~new_U4437 | ~new_U4159 | ~new_U2605 | ~new_U4448;
  assign new_U3386 = ~new_U4222 | ~new_U4187 | ~new_U4465;
  assign new_U3387 = ~new_U2449 | ~new_U2447;
  assign new_U3388 = ~new_U3431 | ~new_U5498;
  assign new_U3389 = ~new_U3256 | ~new_U3262;
  assign new_U3390 = ~new_LT_589_U6;
  assign new_U3391 = ~new_U5524 | ~new_U4230 | ~new_U3287;
  assign new_U3392 = ~new_U3271 | ~STATE2_REG_0_ | ~new_U3265;
  assign new_U3393 = ~new_U3258 | ~new_U3260;
  assign new_U3394 = ~new_U3264 | ~new_U3378;
  assign new_U3395 = ~new_U2427 | ~new_U3281;
  assign new_U3396 = ~new_U4448 | ~new_U3378;
  assign new_U3397 = ~new_U4241 | ~new_U3265;
  assign new_U3398 = ~new_U4178 | ~new_U2452;
  assign new_U3399 = ~STATE2_REG_2_ | ~new_U3258;
  assign new_U3400 = ~REIP_REG_0_;
  assign new_U3401 = ~new_U3744 | ~new_U5550;
  assign new_U3402 = ~new_U4388 | ~new_U4161;
  assign new_U3403 = ~new_U3851 | ~new_U4236;
  assign new_U3404 = ~new_U6042 | ~new_U6041;
  assign new_U3405 = ~STATE2_REG_0_ | ~new_U4482;
  assign new_U3406 = ~new_U4387 | ~new_U7482;
  assign new_U3407 = ~new_U4194 | ~new_U4465;
  assign new_U3408 = ~new_U4182 | ~new_U2431;
  assign new_U3409 = ~new_U4198 | ~STATE2_REG_0_;
  assign new_U3410 = ~new_U4491 | ~new_U3378;
  assign new_U3411 = ~new_U4223 | ~new_U6141;
  assign new_U3412 = ~STATE2_REG_0_ | ~new_U4204;
  assign new_U3413 = ~new_U4223 | ~new_U6252;
  assign new_U3414 = ~new_U2452 | ~new_U3874 | ~STATE2_REG_0_ | ~new_U4237;
  assign new_U3415 = ~new_U3854 | ~new_U2447;
  assign new_U3416 = ~EBX_REG_31_;
  assign new_U3417 = ~new_R2337_U58;
  assign new_U3418 = ~new_U4216 | ~new_U3875;
  assign new_U3419 = ~new_U4197 | ~new_U3249;
  assign new_U3420 = ~new_U3940 | ~new_U3943 | ~new_U3950 | ~new_U3946;
  assign new_U3421 = ~new_U4194 | ~new_U3258;
  assign new_U3422 = ~CODEFETCH_REG;
  assign new_U3423 = ~READREQUEST_REG;
  assign new_U3424 = ~new_U2447 | ~new_U4486;
  assign new_U3425 = ~new_U3254 | ~new_U5470;
  assign new_U3426 = ~new_U4437 | ~STATE2_REG_2_;
  assign new_U3427 = ~STATEBS16_REG | ~new_U3250;
  assign new_U3428 = ~new_U3221;
  assign new_U3429 = ~new_U5467 | ~new_U5466;
  assign new_U3430 = ~new_U2450 | ~new_U3428;
  assign new_U3431 = ~INSTQUEUERD_ADDR_REG_0_ | ~INSTQUEUERD_ADDR_REG_1_ | ~new_U3251;
  assign new_U3432 = ~new_U3261 | ~new_U7052;
  assign new_U3433 = ~new_U4185 | ~new_U4222;
  assign new_U3434 = ~new_U4238 | ~new_U4219 | ~new_U4388;
  assign new_U3435 = ~new_U4238 | ~new_U4219 | ~new_U3265;
  assign new_U3436 = ~new_U4465 | ~new_U4484;
  assign new_U3437 = ~new_U4065 | ~new_U4063 | ~new_U4062 | ~new_U7081;
  assign new_U3438 = ~new_U4242 | ~new_U4254;
  assign new_U3439 = ~new_U4171 | ~new_U3255;
  assign new_U3440 = ~STATE2_REG_0_ | ~new_U2605;
  assign new_U3441 = ~new_U7680 | ~new_U7679;
  assign new_U3442 = ~new_U7683 | ~new_U7682;
  assign new_U3443 = ~new_U7707 | ~new_U7706;
  assign new_U3444 = ~new_U7777 | ~new_U7776;
  assign new_U3445 = ~new_U7622 | ~new_U7621;
  assign n224 = ~new_U7624 | ~new_U7623;
  assign n228 = ~new_U7626 | ~new_U7625;
  assign n232 = ~new_U7628 | ~new_U7627;
  assign new_U3449 = ~new_U7637 | ~new_U7636;
  assign new_U3450 = new_U3242 & new_U4167;
  assign n371 = ~new_U7640 | ~new_U7639;
  assign n376 = ~new_U7642 | ~new_U7641;
  assign n531 = ~new_U7674 | ~new_U7673;
  assign new_U3454 = new_R2182_U24 & new_U2427 & new_U4203;
  assign n1191 = ~new_U7690 | ~new_U7689;
  assign n1196 = ~new_U7697 | ~new_U7696;
  assign new_U3457 = ~new_U7699 | ~new_U7698;
  assign new_U3458 = ~new_U7702 | ~new_U7701;
  assign n1201 = ~new_U7710 | ~new_U7709;
  assign n1206 = ~new_U7712 | ~new_U7711;
  assign n1211 = ~new_U7716 | ~new_U7715;
  assign n1221 = ~new_U7718 | ~new_U7717;
  assign n1226 = ~new_U7723 | ~new_U7722;
  assign n1231 = ~new_U7725 | ~new_U7724;
  assign n1236 = ~new_U7727 | ~new_U7726;
  assign new_U3466 = new_R2358_U91 & new_U4437;
  assign new_U3467 = ~DATAWIDTH_REG_1_ & ~REIP_REG_1_;
  assign n2329 = ~new_U7743 | ~new_U7742;
  assign n2339 = ~new_U7747 | ~new_U7746;
  assign n2344 = ~new_U7749 | ~new_U7748;
  assign n2353 = ~new_U7751 | ~new_U7750;
  assign n2363 = ~new_U7755 | ~new_U7754;
  assign n2372 = ~new_U7759 | ~new_U7758;
  assign n2385 = ~new_U7761 | ~new_U7760;
  assign new_U3475 = new_R2182_U24 & new_U4203;
  assign new_U3476 = ~new_U7763 | ~new_U7762;
  assign new_U3477 = ~new_U7765 | ~new_U7764;
  assign new_U3478 = ~new_U7767 | ~new_U7766;
  assign new_U3479 = ~new_U7769 | ~new_U7768;
  assign new_U3480 = ~new_U7771 | ~new_U7770;
  assign new_U3481 = STATE_REG_1_ & READY_N;
  assign new_U3482 = new_U4356 & new_U3239;
  assign new_U3483 = new_U4358 & new_U3237;
  assign new_U3484 = REQUESTPENDING_REG & STATE_REG_0_;
  assign new_U3485 = ~INSTQUEUERD_ADDR_REG_2_ & ~INSTQUEUERD_ADDR_REG_3_;
  assign new_U3486 = INSTQUEUERD_ADDR_REG_0_ & INSTQUEUERD_ADDR_REG_1_;
  assign new_U3487 = ~INSTQUEUERD_ADDR_REG_1_ & ~INSTQUEUERD_ADDR_REG_3_;
  assign new_U3488 = INSTQUEUERD_ADDR_REG_0_ & INSTQUEUERD_ADDR_REG_2_;
  assign new_U3489 = ~INSTQUEUERD_ADDR_REG_0_ & ~INSTQUEUERD_ADDR_REG_3_;
  assign new_U3490 = INSTQUEUERD_ADDR_REG_1_ & INSTQUEUERD_ADDR_REG_2_;
  assign new_U3491 = ~INSTQUEUERD_ADDR_REG_1_ & ~INSTQUEUERD_ADDR_REG_2_;
  assign new_U3492 = INSTQUEUERD_ADDR_REG_3_ & INSTQUEUERD_ADDR_REG_0_;
  assign new_U3493 = ~INSTQUEUERD_ADDR_REG_0_ & ~INSTQUEUERD_ADDR_REG_2_;
  assign new_U3494 = INSTQUEUERD_ADDR_REG_3_ & INSTQUEUERD_ADDR_REG_1_;
  assign new_U3495 = INSTQUEUERD_ADDR_REG_3_ & INSTQUEUERD_ADDR_REG_2_;
  assign new_U3496 = new_U4371 & new_U4372 & new_U4374 & new_U4373;
  assign new_U3497 = new_U4375 & new_U4376 & new_U4378 & new_U4377;
  assign new_U3498 = new_U4379 & new_U4380 & new_U4382 & new_U4381;
  assign new_U3499 = new_U4383 & new_U4384 & new_U4386 & new_U4385;
  assign new_U3500 = new_U4421 & new_U4422 & new_U4424 & new_U4423;
  assign new_U3501 = new_U4425 & new_U4426 & new_U4428 & new_U4427;
  assign new_U3502 = new_U4429 & new_U4430 & new_U4432 & new_U4431;
  assign new_U3503 = new_U4433 & new_U4434 & new_U4436 & new_U4435;
  assign new_U3504 = new_U4404 & new_U4405 & new_U4407 & new_U4406;
  assign new_U3505 = new_U4408 & new_U4409 & new_U4411 & new_U4410;
  assign new_U3506 = new_U4412 & new_U4413 & new_U4415 & new_U4414;
  assign new_U3507 = new_U4416 & new_U4417 & new_U4419 & new_U4418;
  assign new_U3508 = ~INSTQUEUERD_ADDR_REG_1_ & ~INSTQUEUERD_ADDR_REG_3_;
  assign new_U3509 = INSTQUEUE_REG_5__5_ & INSTQUEUERD_ADDR_REG_0_;
  assign new_U3510 = ~INSTQUEUERD_ADDR_REG_0_ & ~INSTQUEUERD_ADDR_REG_3_;
  assign new_U3511 = INSTQUEUE_REG_6__5_ & INSTQUEUERD_ADDR_REG_1_;
  assign new_U3512 = INSTQUEUERD_ADDR_REG_3_ & INSTQUEUE_REG_8__5_;
  assign new_U3513 = ~INSTQUEUERD_ADDR_REG_0_ & ~INSTQUEUERD_ADDR_REG_2_;
  assign new_U3514 = INSTQUEUE_REG_10__5_ & INSTQUEUERD_ADDR_REG_3_;
  assign new_U3515 = INSTQUEUE_REG_12__5_ & INSTQUEUERD_ADDR_REG_3_;
  assign new_U3516 = ~INSTQUEUERD_ADDR_REG_1_ & ~INSTQUEUERD_ADDR_REG_2_;
  assign new_U3517 = INSTQUEUE_REG_9__5_ & INSTQUEUERD_ADDR_REG_0_;
  assign new_U3518 = new_U4389 & new_U4390 & new_U4392 & new_U4391;
  assign new_U3519 = new_U4393 & new_U4394 & new_U4396 & new_U4395;
  assign new_U3520 = new_U4397 & new_U4398 & new_U4400 & new_U4399;
  assign new_U3521 = new_U4402 & new_U4401;
  assign new_U3522 = ~INSTQUEUERD_ADDR_REG_2_ & ~INSTQUEUERD_ADDR_REG_3_;
  assign new_U3523 = INSTQUEUE_REG_3__6_ & INSTQUEUERD_ADDR_REG_0_;
  assign new_U3524 = new_U4438 & new_U4439 & new_U4441 & new_U4440;
  assign new_U3525 = new_U4444 & new_U4443 & new_U4442;
  assign new_U3526 = new_U4447 & new_U4446 & new_U4445;
  assign new_U3527 = new_U7663 & new_U7664 & new_U7666 & new_U7665;
  assign new_U3528 = ~INSTQUEUERD_ADDR_REG_2_ & ~INSTQUEUERD_ADDR_REG_3_;
  assign new_U3529 = INSTQUEUE_REG_1__4_ & INSTQUEUERD_ADDR_REG_0_;
  assign new_U3530 = ~INSTQUEUERD_ADDR_REG_0_ & ~INSTQUEUERD_ADDR_REG_1_;
  assign new_U3531 = INSTQUEUE_REG_4__4_ & INSTQUEUERD_ADDR_REG_2_;
  assign new_U3532 = ~INSTQUEUERD_ADDR_REG_0_ & ~INSTQUEUERD_ADDR_REG_1_;
  assign new_U3533 = INSTQUEUE_REG_12__4_ & INSTQUEUERD_ADDR_REG_2_;
  assign new_U3534 = INSTQUEUERD_ADDR_REG_0_ & INSTQUEUERD_ADDR_REG_2_;
  assign new_U3535 = INSTQUEUE_REG_13__4_ & INSTQUEUERD_ADDR_REG_3_;
  assign new_U3536 = ~INSTQUEUERD_ADDR_REG_0_ & ~INSTQUEUERD_ADDR_REG_3_;
  assign new_U3537 = INSTQUEUE_REG_6__4_ & INSTQUEUERD_ADDR_REG_2_;
  assign new_U3538 = INSTQUEUERD_ADDR_REG_1_ & INSTQUEUERD_ADDR_REG_2_;
  assign new_U3539 = INSTQUEUE_REG_14__4_ & INSTQUEUERD_ADDR_REG_3_;
  assign new_U3540 = ~INSTQUEUERD_ADDR_REG_1_ & ~INSTQUEUERD_ADDR_REG_2_;
  assign new_U3541 = INSTQUEUE_REG_9__4_ & INSTQUEUERD_ADDR_REG_3_;
  assign new_U3542 = new_U7643 & new_U7644 & new_U7646 & new_U7645;
  assign new_U3543 = new_U7647 & new_U7648 & new_U7650 & new_U7649;
  assign new_U3544 = new_U7651 & new_U7652 & new_U7654 & new_U7653;
  assign new_U3545 = new_U7655 & new_U7656 & new_U7658 & new_U7657;
  assign new_U3546 = new_U7482 & new_U3378 & new_U3270;
  assign new_U3547 = new_U4388 & new_U4448 & new_U2605;
  assign new_U3548 = new_U4466 & new_U4467 & new_U4469 & new_U4468;
  assign new_U3549 = new_U4470 & new_U4471 & new_U4473 & new_U4472;
  assign new_U3550 = new_U4474 & new_U4475 & new_U4477 & new_U4476;
  assign new_U3551 = new_U4478 & new_U4479 & new_U4481 & new_U4480;
  assign new_U3552 = new_U4449 & new_U4450 & new_U4452 & new_U4451;
  assign new_U3553 = new_U4453 & new_U4454 & new_U4456 & new_U4455;
  assign new_U3554 = new_U4457 & new_U4458 & new_U4460 & new_U4459;
  assign new_U3555 = new_U4461 & new_U4462 & new_U4464 & new_U4463;
  assign new_U3556 = new_U4365 & new_U4196;
  assign new_U3557 = new_U4404 & new_U4405 & new_U4407 & new_U4406;
  assign new_U3558 = new_U4408 & new_U4409 & new_U4411 & new_U4410;
  assign new_U3559 = new_U4412 & new_U4413 & new_U4415 & new_U4414;
  assign new_U3560 = new_U4416 & new_U4417 & new_U4419 & new_U4418;
  assign new_U3561 = new_U4389 & new_U4390 & new_U4392 & new_U4391;
  assign new_U3562 = new_U4393 & new_U4394 & new_U4396 & new_U4395;
  assign new_U3563 = new_U4397 & new_U4398 & new_U4400 & new_U4399;
  assign new_U3564 = new_U4402 & new_U4401;
  assign new_U3565 = new_U4387 & new_U4159;
  assign new_U3566 = new_U4237 & new_U3270;
  assign new_U3567 = new_U7482 & new_U4388 & new_U3271 & new_U3270;
  assign new_U3568 = new_U4205 & new_U3387;
  assign new_U3569 = STATE2_REG_2_ & new_U7591;
  assign new_U3570 = new_U4503 & new_U3284;
  assign new_U3571 = new_U2427 & new_U3244;
  assign new_U3572 = STATE2_REG_3_ & STATE2_REG_0_;
  assign new_U3573 = new_U4234 & new_U4229;
  assign new_U3574 = new_U3573 & new_U4511;
  assign new_U3575 = new_U4212 & new_U4540 & new_U4541;
  assign new_U3576 = new_U4550 & new_U4549 & new_U4548;
  assign new_U3577 = new_U4555 & new_U4554 & new_U4553;
  assign new_U3578 = new_U4560 & new_U4559 & new_U4558;
  assign new_U3579 = new_U4565 & new_U4564 & new_U4563;
  assign new_U3580 = new_U4570 & new_U4569 & new_U4568;
  assign new_U3581 = new_U4575 & new_U4574 & new_U4573;
  assign new_U3582 = new_U4580 & new_U4579 & new_U4578;
  assign new_U3583 = new_U4585 & new_U4584 & new_U4583;
  assign new_U3584 = new_U4212 & new_U4598 & new_U4599;
  assign new_U3585 = new_U4608 & new_U4607 & new_U4606;
  assign new_U3586 = new_U4613 & new_U4612 & new_U4611;
  assign new_U3587 = new_U4618 & new_U4617 & new_U4616;
  assign new_U3588 = new_U4623 & new_U4622 & new_U4621;
  assign new_U3589 = new_U4628 & new_U4627 & new_U4626;
  assign new_U3590 = new_U4633 & new_U4632 & new_U4631;
  assign new_U3591 = new_U4638 & new_U4637 & new_U4636;
  assign new_U3592 = new_U4643 & new_U4642 & new_U4641;
  assign new_U3593 = new_U4212 & new_U4657 & new_U4658;
  assign new_U3594 = new_U4667 & new_U4666 & new_U4665;
  assign new_U3595 = new_U4672 & new_U4671 & new_U4670;
  assign new_U3596 = new_U4677 & new_U4676 & new_U4675;
  assign new_U3597 = new_U4682 & new_U4681 & new_U4680;
  assign new_U3598 = new_U4687 & new_U4686 & new_U4685;
  assign new_U3599 = new_U4692 & new_U4691 & new_U4690;
  assign new_U3600 = new_U4697 & new_U4696 & new_U4695;
  assign new_U3601 = new_U4702 & new_U4701 & new_U4700;
  assign new_U3602 = new_U4212 & new_U4714 & new_U4715;
  assign new_U3603 = new_U4724 & new_U4723 & new_U4722;
  assign new_U3604 = new_U4729 & new_U4728 & new_U4727;
  assign new_U3605 = new_U4734 & new_U4733 & new_U4732;
  assign new_U3606 = new_U4739 & new_U4738 & new_U4737;
  assign new_U3607 = new_U4744 & new_U4743 & new_U4742;
  assign new_U3608 = new_U4749 & new_U4748 & new_U4747;
  assign new_U3609 = new_U4754 & new_U4753 & new_U4752;
  assign new_U3610 = new_U4759 & new_U4758 & new_U4757;
  assign new_U3611 = new_U4212 & new_U4772 & new_U4773;
  assign new_U3612 = new_U4782 & new_U4781 & new_U4780;
  assign new_U3613 = new_U4787 & new_U4786 & new_U4785;
  assign new_U3614 = new_U4792 & new_U4791 & new_U4790;
  assign new_U3615 = new_U4797 & new_U4796 & new_U4795;
  assign new_U3616 = new_U4802 & new_U4801 & new_U4800;
  assign new_U3617 = new_U4807 & new_U4806 & new_U4805;
  assign new_U3618 = new_U4812 & new_U4811 & new_U4810;
  assign new_U3619 = new_U4817 & new_U4816 & new_U4815;
  assign new_U3620 = new_U4212 & new_U4829 & new_U4830;
  assign new_U3621 = new_U4839 & new_U4838 & new_U4837;
  assign new_U3622 = new_U4844 & new_U4843 & new_U4842;
  assign new_U3623 = new_U4849 & new_U4848 & new_U4847;
  assign new_U3624 = new_U4854 & new_U4853 & new_U4852;
  assign new_U3625 = new_U4859 & new_U4858 & new_U4857;
  assign new_U3626 = new_U4864 & new_U4863 & new_U4862;
  assign new_U3627 = new_U4869 & new_U4868 & new_U4867;
  assign new_U3628 = new_U4874 & new_U4873 & new_U4872;
  assign new_U3629 = new_U4212 & new_U4887 & new_U4888;
  assign new_U3630 = new_U4897 & new_U4896 & new_U4895;
  assign new_U3631 = new_U4902 & new_U4901 & new_U4900;
  assign new_U3632 = new_U4907 & new_U4906 & new_U4905;
  assign new_U3633 = new_U4912 & new_U4911 & new_U4910;
  assign new_U3634 = new_U4917 & new_U4916 & new_U4915;
  assign new_U3635 = new_U4922 & new_U4921 & new_U4920;
  assign new_U3636 = new_U4927 & new_U4926 & new_U4925;
  assign new_U3637 = new_U4932 & new_U4931 & new_U4930;
  assign new_U3638 = new_U4212 & new_U4944 & new_U4945;
  assign new_U3639 = new_U4954 & new_U4953 & new_U4952;
  assign new_U3640 = new_U4959 & new_U4958 & new_U4957;
  assign new_U3641 = new_U4964 & new_U4963 & new_U4962;
  assign new_U3642 = new_U4969 & new_U4968 & new_U4967;
  assign new_U3643 = new_U4974 & new_U4973 & new_U4972;
  assign new_U3644 = new_U4979 & new_U4978 & new_U4977;
  assign new_U3645 = new_U4984 & new_U4983 & new_U4982;
  assign new_U3646 = new_U4989 & new_U4988 & new_U4987;
  assign new_U3647 = new_U4212 & new_U5000 & new_U5001;
  assign new_U3648 = new_U5010 & new_U5009 & new_U5008;
  assign new_U3649 = new_U5015 & new_U5014 & new_U5013;
  assign new_U3650 = new_U5020 & new_U5019 & new_U5018;
  assign new_U3651 = new_U5025 & new_U5024 & new_U5023;
  assign new_U3652 = new_U5030 & new_U5029 & new_U5028;
  assign new_U3653 = new_U5035 & new_U5034 & new_U5033;
  assign new_U3654 = new_U5040 & new_U5039 & new_U5038;
  assign new_U3655 = new_U5045 & new_U5044 & new_U5043;
  assign new_U3656 = new_U4212 & new_U5057 & new_U5058;
  assign new_U3657 = new_U5067 & new_U5066 & new_U5065;
  assign new_U3658 = new_U5072 & new_U5071 & new_U5070;
  assign new_U3659 = new_U5077 & new_U5076 & new_U5075;
  assign new_U3660 = new_U5082 & new_U5081 & new_U5080;
  assign new_U3661 = new_U5087 & new_U5086 & new_U5085;
  assign new_U3662 = new_U5092 & new_U5091 & new_U5090;
  assign new_U3663 = new_U5097 & new_U5096 & new_U5095;
  assign new_U3664 = new_U5102 & new_U5101 & new_U5100;
  assign new_U3665 = new_U4212 & new_U5115 & new_U5116;
  assign new_U3666 = new_U5125 & new_U5124 & new_U5123;
  assign new_U3667 = new_U5130 & new_U5129 & new_U5128;
  assign new_U3668 = new_U5135 & new_U5134 & new_U5133;
  assign new_U3669 = new_U5140 & new_U5139 & new_U5138;
  assign new_U3670 = new_U5145 & new_U5144 & new_U5143;
  assign new_U3671 = new_U5150 & new_U5149 & new_U5148;
  assign new_U3672 = new_U5155 & new_U5154 & new_U5153;
  assign new_U3673 = new_U5160 & new_U5159 & new_U5158;
  assign new_U3674 = new_U4212 & new_U5172 & new_U5173;
  assign new_U3675 = new_U5182 & new_U5181 & new_U5180;
  assign new_U3676 = new_U5187 & new_U5186 & new_U5185;
  assign new_U3677 = new_U5192 & new_U5191 & new_U5190;
  assign new_U3678 = new_U5197 & new_U5196 & new_U5195;
  assign new_U3679 = new_U5202 & new_U5201 & new_U5200;
  assign new_U3680 = new_U5207 & new_U5206 & new_U5205;
  assign new_U3681 = new_U5212 & new_U5211 & new_U5210;
  assign new_U3682 = new_U5217 & new_U5216 & new_U5215;
  assign new_U3683 = new_U4212 & new_U5230 & new_U5231;
  assign new_U3684 = new_U5240 & new_U5239 & new_U5238;
  assign new_U3685 = new_U5245 & new_U5244 & new_U5243;
  assign new_U3686 = new_U5250 & new_U5249 & new_U5248;
  assign new_U3687 = new_U5255 & new_U5254 & new_U5253;
  assign new_U3688 = new_U5260 & new_U5259 & new_U5258;
  assign new_U3689 = new_U5265 & new_U5264 & new_U5263;
  assign new_U3690 = new_U5270 & new_U5269 & new_U5268;
  assign new_U3691 = new_U5275 & new_U5274 & new_U5273;
  assign new_U3692 = new_U4212 & new_U5287 & new_U5288;
  assign new_U3693 = new_U5297 & new_U5296 & new_U5295;
  assign new_U3694 = new_U5302 & new_U5301 & new_U5300;
  assign new_U3695 = new_U5307 & new_U5306 & new_U5305;
  assign new_U3696 = new_U5312 & new_U5311 & new_U5310;
  assign new_U3697 = new_U5317 & new_U5316 & new_U5315;
  assign new_U3698 = new_U5322 & new_U5321 & new_U5320;
  assign new_U3699 = new_U5327 & new_U5326 & new_U5325;
  assign new_U3700 = new_U5332 & new_U5331 & new_U5330;
  assign new_U3701 = new_U4212 & new_U5345 & new_U5346;
  assign new_U3702 = new_U5355 & new_U5354 & new_U5353;
  assign new_U3703 = new_U5360 & new_U5359 & new_U5358;
  assign new_U3704 = new_U5365 & new_U5364 & new_U5363;
  assign new_U3705 = new_U5370 & new_U5369 & new_U5368;
  assign new_U3706 = new_U5375 & new_U5374 & new_U5373;
  assign new_U3707 = new_U5380 & new_U5379 & new_U5378;
  assign new_U3708 = new_U5385 & new_U5384 & new_U5383;
  assign new_U3709 = new_U5390 & new_U5389 & new_U5388;
  assign new_U3710 = new_U4212 & new_U5402 & new_U5403;
  assign new_U3711 = new_U5412 & new_U5411 & new_U5410;
  assign new_U3712 = new_U5417 & new_U5416 & new_U5415;
  assign new_U3713 = new_U5422 & new_U5421 & new_U5420;
  assign new_U3714 = new_U5427 & new_U5426 & new_U5425;
  assign new_U3715 = new_U5431 & new_U5430 & new_U5429;
  assign new_U3716 = new_U5436 & new_U5435 & new_U5434;
  assign new_U3717 = new_U5441 & new_U5440 & new_U5439;
  assign new_U3718 = new_U5446 & new_U5445 & new_U5444;
  assign new_U3719 = FLUSH_REG & STATE2_REG_0_;
  assign new_U3720 = new_U4482 & new_U4387;
  assign new_U3721 = new_U4485 & new_U3244;
  assign new_U3722 = new_U4198 & new_U3244;
  assign new_U3723 = new_U7484 & new_U4205;
  assign new_U3724 = new_U5459 & new_U5460;
  assign new_U3725 = new_U3724 & new_U5458;
  assign new_U3726 = new_U3725 & new_U2518;
  assign new_U3727 = new_U5463 & new_U4230;
  assign new_U3728 = new_U5474 & new_U5473;
  assign new_U3729 = new_U4437 & new_U4388;
  assign new_U3730 = new_U5484 & new_U3380;
  assign new_U3731 = new_U5486 & new_U5485;
  assign new_U3732 = new_U3731 & new_U3730 & new_U5488 & new_U7615;
  assign new_U3733 = new_U4251 & new_U3384;
  assign new_U3734 = new_U3266 & new_U2520 & new_U3733 & new_U3398 & new_U3275;
  assign new_U3735 = new_U3736 & new_U5490;
  assign new_U3736 = new_U5493 & new_U5492;
  assign new_U3737 = new_U5501 & new_U7705 & new_U7704;
  assign new_U3738 = new_U5512 & new_U5510;
  assign new_U3739 = new_U5531 & new_U5532;
  assign new_U3740 = new_U5535 & new_U5536;
  assign new_U3741 = new_U5540 & new_U5541;
  assign new_U3742 = new_U5546 & new_U3244;
  assign new_U3743 = new_U3271 & new_U3394;
  assign new_U3744 = new_U5551 & new_U5549;
  assign new_U3745 = new_U5555 & new_U3385 & new_U3386;
  assign new_U3746 = new_U3745 & new_U2520 & new_U5556;
  assign new_U3747 = new_U4174 & new_U3271;
  assign new_U3748 = new_U3435 & new_U3275 & new_U4205;
  assign new_U3749 = new_U5554 & new_U7495;
  assign new_U3750 = new_U7496 & STATE2_REG_2_;
  assign new_U3751 = new_U5559 & new_U5558;
  assign new_U3752 = new_U5561 & new_U5560;
  assign new_U3753 = new_U5563 & new_U5564;
  assign new_U3754 = new_U3753 & new_U5562;
  assign new_U3755 = new_U5566 & new_U5565;
  assign new_U3756 = new_U5568 & new_U5567;
  assign new_U3757 = new_U5570 & new_U5571;
  assign new_U3758 = new_U3757 & new_U5569;
  assign new_U3759 = new_U5573 & new_U5572;
  assign new_U3760 = new_U5575 & new_U5574;
  assign new_U3761 = new_U5577 & new_U5578;
  assign new_U3762 = new_U3761 & new_U5576;
  assign new_U3763 = new_U5582 & new_U5580 & new_U5579;
  assign new_U3764 = new_U5581 & new_U3765 & new_U5583;
  assign new_U3765 = new_U5584 & new_U5585;
  assign new_U3766 = new_U5589 & new_U5587 & new_U5586;
  assign new_U3767 = new_U5591 & new_U5592;
  assign new_U3768 = new_U3767 & new_U5590;
  assign new_U3769 = new_U5596 & new_U5594 & new_U5593;
  assign new_U3770 = new_U5598 & new_U5599;
  assign new_U3771 = new_U3770 & new_U5597;
  assign new_U3772 = new_U5603 & new_U5601 & new_U5600;
  assign new_U3773 = new_U5605 & new_U5606;
  assign new_U3774 = new_U3773 & new_U5604;
  assign new_U3775 = new_U5610 & new_U5608 & new_U5607;
  assign new_U3776 = new_U5612 & new_U5613;
  assign new_U3777 = new_U3776 & new_U5611;
  assign new_U3778 = new_U5617 & new_U5615 & new_U5614;
  assign new_U3779 = new_U5619 & new_U5620;
  assign new_U3780 = new_U3779 & new_U5618;
  assign new_U3781 = new_U5624 & new_U5622 & new_U5621;
  assign new_U3782 = new_U5626 & new_U5627;
  assign new_U3783 = new_U3782 & new_U5625;
  assign new_U3784 = new_U5631 & new_U5629 & new_U5628;
  assign new_U3785 = new_U5633 & new_U5634;
  assign new_U3786 = new_U3785 & new_U5632;
  assign new_U3787 = new_U5638 & new_U5636 & new_U5635;
  assign new_U3788 = new_U5640 & new_U5641;
  assign new_U3789 = new_U3788 & new_U5639;
  assign new_U3790 = new_U5645 & new_U5643 & new_U5642;
  assign new_U3791 = new_U5647 & new_U5648;
  assign new_U3792 = new_U3791 & new_U5646;
  assign new_U3793 = new_U5650 & new_U5652;
  assign new_U3794 = new_U5654 & new_U5655;
  assign new_U3795 = new_U3794 & new_U5653;
  assign new_U3796 = new_U5657 & new_U5659;
  assign new_U3797 = new_U5661 & new_U5662;
  assign new_U3798 = new_U3797 & new_U5660;
  assign new_U3799 = new_U5664 & new_U5666;
  assign new_U3800 = new_U5668 & new_U5669;
  assign new_U3801 = new_U3800 & new_U5667;
  assign new_U3802 = new_U5671 & new_U5673;
  assign new_U3803 = new_U5675 & new_U5676;
  assign new_U3804 = new_U3803 & new_U5674;
  assign new_U3805 = new_U5678 & new_U5680;
  assign new_U3806 = new_U5682 & new_U5683;
  assign new_U3807 = new_U3806 & new_U5681;
  assign new_U3808 = new_U5685 & new_U5687;
  assign new_U3809 = new_U5689 & new_U5690;
  assign new_U3810 = new_U3809 & new_U5688;
  assign new_U3811 = new_U5692 & new_U5694;
  assign new_U3812 = new_U5696 & new_U5697;
  assign new_U3813 = new_U3812 & new_U5695;
  assign new_U3814 = new_U5699 & new_U5701;
  assign new_U3815 = new_U5703 & new_U5704;
  assign new_U3816 = new_U3815 & new_U5702;
  assign new_U3817 = new_U5706 & new_U5708;
  assign new_U3818 = new_U5710 & new_U5711;
  assign new_U3819 = new_U3818 & new_U5709;
  assign new_U3820 = new_U5713 & new_U5715;
  assign new_U3821 = new_U5717 & new_U5718;
  assign new_U3822 = new_U3821 & new_U5716;
  assign new_U3823 = new_U5720 & new_U5722;
  assign new_U3824 = new_U5724 & new_U5725;
  assign new_U3825 = new_U3824 & new_U5723;
  assign new_U3826 = new_U5727 & new_U5729;
  assign new_U3827 = new_U5731 & new_U5732;
  assign new_U3828 = new_U3827 & new_U5730;
  assign new_U3829 = new_U5734 & new_U5736;
  assign new_U3830 = new_U5738 & new_U5739;
  assign new_U3831 = new_U3830 & new_U5737;
  assign new_U3832 = new_U5741 & new_U5743;
  assign new_U3833 = new_U5745 & new_U5746;
  assign new_U3834 = new_U3833 & new_U5744;
  assign new_U3835 = new_U5748 & new_U5750;
  assign new_U3836 = new_U5752 & new_U5753;
  assign new_U3837 = new_U3836 & new_U5751;
  assign new_U3838 = new_U5755 & new_U5757;
  assign new_U3839 = new_U5759 & new_U5760;
  assign new_U3840 = new_U3839 & new_U5758;
  assign new_U3841 = new_U5762 & new_U5764;
  assign new_U3842 = new_U5766 & new_U5767;
  assign new_U3843 = new_U3842 & new_U5765;
  assign new_U3844 = new_U5769 & new_U5771;
  assign new_U3845 = new_U5773 & new_U5774;
  assign new_U3846 = new_U3845 & new_U5772;
  assign new_U3847 = new_U5776 & new_U5778;
  assign new_U3848 = new_U5780 & new_U5781;
  assign new_U3849 = new_U3848 & new_U5779;
  assign new_U3850 = new_U7482 & new_U3270 & new_U3249;
  assign new_U3851 = new_U5782 & new_U3395;
  assign new_U3852 = STATE2_REG_1_ & STATEBS16_REG;
  assign new_U3853 = new_U2368 & new_U3271;
  assign new_U3854 = new_U2449 & STATE2_REG_0_;
  assign new_U3855 = new_U4196 & new_U2368;
  assign new_U3856 = new_U6093 & new_U6094;
  assign new_U3857 = new_U6096 & new_U6097;
  assign new_U3858 = new_U6099 & new_U6100;
  assign new_U3859 = new_U6102 & new_U6103;
  assign new_U3860 = new_U6105 & new_U6106;
  assign new_U3861 = new_U6108 & new_U6109;
  assign new_U3862 = new_U6111 & new_U6112;
  assign new_U3863 = new_U6114 & new_U6115;
  assign new_U3864 = new_U6117 & new_U6118;
  assign new_U3865 = new_U6120 & new_U6121;
  assign new_U3866 = new_U6123 & new_U6124;
  assign new_U3867 = new_U6126 & new_U6127;
  assign new_U3868 = new_U6129 & new_U6130;
  assign new_U3869 = new_U6132 & new_U6133;
  assign new_U3870 = new_U6135 & new_U6136;
  assign new_U3871 = new_U6139 & new_U6138;
  assign new_U3872 = new_U2605 & new_U3378;
  assign new_U3873 = new_U7482 & STATE2_REG_0_ & new_U3258;
  assign new_U3874 = new_U4387 & new_U4159;
  assign new_U3875 = new_U6350 & new_U4229 & new_U4232;
  assign new_U3876 = ~READY_N & ~STATEBS16_REG;
  assign new_U3877 = new_U4482 & new_U4174;
  assign new_U3878 = new_U6359 & new_U6362 & new_U6363 & new_U6361 & new_U6360;
  assign new_U3879 = new_U6367 & new_U6370 & new_U6371 & new_U6369 & new_U6368;
  assign new_U3880 = new_U6375 & new_U6378 & new_U6379 & new_U6377 & new_U6376;
  assign new_U3881 = new_U6383 & new_U6386 & new_U6387 & new_U6385 & new_U6384;
  assign new_U3882 = new_U6388 & new_U4215;
  assign new_U3883 = new_U6394 & new_U6395 & new_U6393 & new_U6392;
  assign new_U3884 = new_U6396 & new_U4215;
  assign new_U3885 = new_U6399 & new_U6402 & new_U6403 & new_U6401 & new_U6400;
  assign new_U3886 = new_U6404 & new_U4215;
  assign new_U3887 = new_U6409 & new_U6410 & new_U6407;
  assign new_U3888 = new_U6411 & new_U4215;
  assign new_U3889 = new_U6416 & new_U6417 & new_U6414;
  assign new_U3890 = new_U6418 & new_U4215;
  assign new_U3891 = new_U6423 & new_U6424 & new_U6421;
  assign new_U3892 = new_U6425 & new_U4215;
  assign new_U3893 = new_U6430 & new_U6431 & new_U6428;
  assign new_U3894 = new_U6432 & new_U4215;
  assign new_U3895 = new_U6437 & new_U6438 & new_U6435;
  assign new_U3896 = new_U6439 & new_U4215;
  assign new_U3897 = new_U6444 & new_U6445 & new_U6442;
  assign new_U3898 = new_U6446 & new_U4215;
  assign new_U3899 = new_U6451 & new_U6452 & new_U6449;
  assign new_U3900 = new_U6453 & new_U4215;
  assign new_U3901 = new_U6458 & new_U6459 & new_U6456;
  assign new_U3902 = new_U6460 & new_U4215;
  assign new_U3903 = new_U6465 & new_U6466 & new_U6463;
  assign new_U3904 = new_U6467 & new_U4215;
  assign new_U3905 = new_U6472 & new_U6473 & new_U6470;
  assign new_U3906 = new_U6474 & new_U4215;
  assign new_U3907 = new_U6479 & new_U6480 & new_U6477;
  assign new_U3908 = new_U4215 & new_U6482;
  assign new_U3909 = new_U6486 & new_U6487 & new_U6484;
  assign new_U3910 = new_U4215 & new_U6489;
  assign new_U3911 = new_U6493 & new_U6494 & new_U6491;
  assign new_U3912 = new_U4215 & new_U6496;
  assign new_U3913 = new_U6500 & new_U6501 & new_U6498;
  assign new_U3914 = new_U6505 & new_U6503;
  assign new_U3915 = new_U6507 & new_U6508;
  assign new_U3916 = new_U6512 & new_U6510;
  assign new_U3917 = new_U6514 & new_U6515;
  assign new_U3918 = new_U6519 & new_U6517;
  assign new_U3919 = new_U6521 & new_U6522;
  assign new_U3920 = new_U6526 & new_U6524;
  assign new_U3921 = new_U6528 & new_U6529;
  assign new_U3922 = new_U6533 & new_U6531;
  assign new_U3923 = new_U6535 & new_U6536;
  assign new_U3924 = new_U6540 & new_U6538;
  assign new_U3925 = new_U6542 & new_U6543;
  assign new_U3926 = new_U6547 & new_U6545;
  assign new_U3927 = new_U6549 & new_U6550;
  assign new_U3928 = new_U6554 & new_U6552;
  assign new_U3929 = new_U6556 & new_U6557;
  assign new_U3930 = new_U6561 & new_U6559;
  assign new_U3931 = new_U6563 & new_U6564;
  assign new_U3932 = new_U6568 & new_U6566;
  assign new_U3933 = new_U6570 & new_U6571;
  assign new_U3934 = new_U6575 & new_U6573;
  assign new_U3935 = new_U6577 & new_U6578;
  assign new_U3936 = new_U6582 & new_U6580;
  assign new_U3937 = new_U6584 & new_U6585;
  assign new_U3938 = ~DATAWIDTH_REG_5_ & ~DATAWIDTH_REG_4_ & ~DATAWIDTH_REG_2_ & ~DATAWIDTH_REG_3_;
  assign new_U3939 = ~DATAWIDTH_REG_9_ & ~DATAWIDTH_REG_8_ & ~DATAWIDTH_REG_6_ & ~DATAWIDTH_REG_7_;
  assign new_U3940 = new_U3939 & new_U3938;
  assign new_U3941 = ~DATAWIDTH_REG_13_ & ~DATAWIDTH_REG_12_ & ~DATAWIDTH_REG_10_ & ~DATAWIDTH_REG_11_;
  assign new_U3942 = ~DATAWIDTH_REG_17_ & ~DATAWIDTH_REG_16_ & ~DATAWIDTH_REG_14_ & ~DATAWIDTH_REG_15_;
  assign new_U3943 = new_U3942 & new_U3941;
  assign new_U3944 = ~DATAWIDTH_REG_21_ & ~DATAWIDTH_REG_20_ & ~DATAWIDTH_REG_18_ & ~DATAWIDTH_REG_19_;
  assign new_U3945 = ~DATAWIDTH_REG_25_ & ~DATAWIDTH_REG_24_ & ~DATAWIDTH_REG_22_ & ~DATAWIDTH_REG_23_;
  assign new_U3946 = new_U3945 & new_U3944;
  assign new_U3947 = ~DATAWIDTH_REG_26_ & ~DATAWIDTH_REG_27_;
  assign new_U3948 = ~DATAWIDTH_REG_28_ & ~DATAWIDTH_REG_29_;
  assign new_U3949 = ~DATAWIDTH_REG_30_ & ~DATAWIDTH_REG_31_;
  assign new_U3950 = new_U3947 & new_U3948 & new_U3949 & new_U6586;
  assign new_U3951 = ~DATAWIDTH_REG_1_ & ~REIP_REG_0_ & ~DATAWIDTH_REG_0_;
  assign new_U3952 = STATE2_REG_2_ & new_U3244;
  assign new_U3953 = new_U6596 & new_U3285;
  assign new_U3954 = ~READY_N & ~STATE2_REG_0_;
  assign new_U3955 = new_U6590 & new_U3294 & new_U3395;
  assign new_U3956 = STATE2_REG_2_ & new_U3274;
  assign new_U3957 = new_U4223 & new_U4194;
  assign new_U3958 = new_U6606 & new_U6607 & new_U6609 & new_U6608;
  assign new_U3959 = new_U6610 & new_U6611 & new_U6613 & new_U6612;
  assign new_U3960 = new_U6614 & new_U6615 & new_U6617 & new_U6616;
  assign new_U3961 = new_U6618 & new_U6619 & new_U6621 & new_U6620;
  assign new_U3962 = new_U6622 & new_U6623 & new_U6625 & new_U6624;
  assign new_U3963 = new_U6626 & new_U6627 & new_U6629 & new_U6628;
  assign new_U3964 = new_U6630 & new_U6631 & new_U6633 & new_U6632;
  assign new_U3965 = new_U6634 & new_U6635 & new_U6637 & new_U6636;
  assign new_U3966 = new_U6638 & new_U6639 & new_U6641 & new_U6640;
  assign new_U3967 = new_U6642 & new_U6643 & new_U6645 & new_U6644;
  assign new_U3968 = new_U6646 & new_U6647 & new_U6649 & new_U6648;
  assign new_U3969 = new_U6650 & new_U6651 & new_U6653 & new_U6652;
  assign new_U3970 = new_U6654 & new_U6655 & new_U6657 & new_U6656;
  assign new_U3971 = new_U6658 & new_U6659 & new_U6661 & new_U6660;
  assign new_U3972 = new_U6662 & new_U6663 & new_U6665 & new_U6664;
  assign new_U3973 = new_U6666 & new_U6667 & new_U7601 & new_U6668;
  assign new_U3974 = new_U6669 & new_U6670 & new_U6672 & new_U6671;
  assign new_U3975 = new_U6673 & new_U6674 & new_U6676 & new_U6675;
  assign new_U3976 = new_U6677 & new_U6678 & new_U6680 & new_U6679;
  assign new_U3977 = new_U6681 & new_U6682 & new_U6684 & new_U6683;
  assign new_U3978 = new_U6685 & new_U6686 & new_U6688 & new_U6687;
  assign new_U3979 = new_U6689 & new_U6690 & new_U6692 & new_U6691;
  assign new_U3980 = new_U6693 & new_U6694 & new_U6696 & new_U6695;
  assign new_U3981 = new_U6697 & new_U6698 & new_U6700 & new_U6699;
  assign new_U3982 = new_U6701 & new_U6702 & new_U6704 & new_U6703;
  assign new_U3983 = new_U6705 & new_U6706 & new_U6708 & new_U6707;
  assign new_U3984 = new_U6709 & new_U6710 & new_U6712 & new_U6711;
  assign new_U3985 = new_U6713 & new_U6714 & new_U6716 & new_U6715;
  assign new_U3986 = new_U6717 & new_U6718 & new_U6720 & new_U6719;
  assign new_U3987 = new_U6721 & new_U6722 & new_U6724 & new_U6723;
  assign new_U3988 = new_U6725 & new_U6726 & new_U6728 & new_U6727;
  assign new_U3989 = new_U6729 & new_U6730 & new_U6732 & new_U6731;
  assign new_U3990 = new_U6737 & new_U6736;
  assign new_U3991 = new_U6740 & new_U6739;
  assign new_U3992 = new_U6743 & new_U6742;
  assign new_U3993 = new_U6746 & new_U6745;
  assign new_U3994 = new_U6748 & new_U3995;
  assign new_U3995 = new_U6750 & new_U6749;
  assign new_U3996 = new_U6752 & new_U6753;
  assign new_U3997 = new_U6762 & new_U6760 & new_U6761;
  assign new_U3998 = new_U6764 & new_U6765;
  assign new_U3999 = new_U6771 & new_U6769 & new_U6770;
  assign new_U4000 = new_U6775 & new_U6773 & new_U6774;
  assign new_U4001 = new_U6779 & new_U6777 & new_U6778;
  assign new_U4002 = new_U6783 & new_U6781 & new_U6782;
  assign new_U4003 = new_U6787 & new_U6785 & new_U6786;
  assign new_U4004 = new_U6791 & new_U6789 & new_U6790;
  assign new_U4005 = new_U6795 & new_U6793 & new_U6794;
  assign new_U4006 = new_U6799 & new_U6797 & new_U6798;
  assign new_U4007 = new_U6803 & new_U6801 & new_U6802;
  assign new_U4008 = new_U6807 & new_U6805 & new_U6806;
  assign new_U4009 = new_U6809 & new_U6810;
  assign new_U4010 = new_U6816 & new_U6814 & new_U6815;
  assign new_U4011 = new_U6820 & new_U6818 & new_U6819;
  assign new_U4012 = new_U6824 & new_U6822 & new_U6823;
  assign new_U4013 = new_U6828 & new_U6826 & new_U6827;
  assign new_U4014 = new_U6846 & new_U6845;
  assign new_U4015 = new_U6848 & new_U6849;
  assign new_U4016 = new_U3270 & new_U7482 & new_U6876;
  assign new_U4017 = new_U6880 & new_U6881 & new_U6883 & new_U6882;
  assign new_U4018 = new_U6884 & new_U6885 & new_U6887 & new_U6886;
  assign new_U4019 = new_U6888 & new_U6889 & new_U6891 & new_U6890;
  assign new_U4020 = new_U6892 & new_U6893 & new_U6895 & new_U6894;
  assign new_U4021 = new_U6898 & new_U6899 & new_U6901 & new_U6900;
  assign new_U4022 = new_U6902 & new_U6903 & new_U6905 & new_U6904;
  assign new_U4023 = new_U6906 & new_U6907 & new_U6909 & new_U6908;
  assign new_U4024 = new_U6910 & new_U6911 & new_U6913 & new_U6912;
  assign new_U4025 = new_U6929 & new_U6930 & new_U6932 & new_U6931;
  assign new_U4026 = new_U6933 & new_U6934 & new_U6936 & new_U6935;
  assign new_U4027 = new_U6937 & new_U6938 & new_U6940 & new_U6939;
  assign new_U4028 = new_U6941 & new_U6942 & new_U6944 & new_U6943;
  assign new_U4029 = new_U6946 & new_U6947 & new_U6949 & new_U6948;
  assign new_U4030 = new_U6950 & new_U6951 & new_U6953 & new_U6952;
  assign new_U4031 = new_U6954 & new_U6955 & new_U6957 & new_U6956;
  assign new_U4032 = new_U6958 & new_U6959 & new_U6961 & new_U6960;
  assign new_U4033 = new_U6963 & new_U6964 & new_U6966 & new_U6965;
  assign new_U4034 = new_U6967 & new_U6968 & new_U6970 & new_U6969;
  assign new_U4035 = new_U6971 & new_U6972 & new_U6974 & new_U6973;
  assign new_U4036 = new_U6975 & new_U6976 & new_U6978 & new_U6977;
  assign new_U4037 = new_U6980 & new_U6981 & new_U6983 & new_U6982;
  assign new_U4038 = new_U6984 & new_U6985 & new_U6987 & new_U6986;
  assign new_U4039 = new_U6988 & new_U6989 & new_U6991 & new_U6990;
  assign new_U4040 = new_U6992 & new_U6993 & new_U7602 & new_U6994;
  assign new_U4041 = new_U6995 & new_U6996 & new_U6998 & new_U6997;
  assign new_U4042 = new_U6999 & new_U7000 & new_U7002 & new_U7001;
  assign new_U4043 = new_U7003 & new_U7004 & new_U7006 & new_U7005;
  assign new_U4044 = new_U7007 & new_U7008 & new_U7010 & new_U7009;
  assign new_U4045 = new_U7012 & new_U7013 & new_U7015 & new_U7014;
  assign new_U4046 = new_U7016 & new_U7017 & new_U7019 & new_U7018;
  assign new_U4047 = new_U7020 & new_U7021 & new_U7023 & new_U7022;
  assign new_U4048 = new_U7024 & new_U7025 & new_U7027 & new_U7026;
  assign new_U4049 = new_U7047 & new_U3430;
  assign new_U4050 = STATE2_REG_0_ & new_U7050;
  assign new_U4051 = new_U7054 & new_U7055 & new_U7057 & new_U7056;
  assign new_U4052 = new_U7058 & new_U7059 & new_U7061 & new_U7060;
  assign new_U4053 = new_U7062 & new_U7063 & new_U7065 & new_U7064;
  assign new_U4054 = new_U7066 & new_U7067 & new_U7069 & new_U7068;
  assign new_U4055 = new_U4244 & STATE2_REG_0_;
  assign new_U4056 = new_U4389 & new_U4391 & new_U4393 & new_U4392;
  assign new_U4057 = new_U4396 & new_U4395 & new_U4394;
  assign new_U4058 = new_U4397 & new_U4398 & new_U4400 & new_U4399;
  assign new_U4059 = new_U4402 & new_U4401;
  assign new_U4060 = new_U4388 & new_U3378;
  assign new_U4061 = STATE2_REG_0_ & new_U3271;
  assign new_U4062 = new_U7078 & new_U7077;
  assign new_U4063 = new_U7461 & new_U7460 & new_U3421;
  assign new_U4064 = new_U7462 & new_U7463 & new_U7464;
  assign new_U4065 = new_U4064 & new_U2606 & new_U7465;
  assign new_U4066 = new_U7085 & new_U7083;
  assign new_U4067 = new_U7086 & new_U7087 & new_U7089 & new_U7088;
  assign new_U4068 = new_U7090 & new_U7091 & new_U7093 & new_U7092;
  assign new_U4069 = new_U7094 & new_U7095 & new_U7097 & new_U7096;
  assign new_U4070 = new_U7098 & new_U7099 & new_U7101 & new_U7100;
  assign new_U4071 = new_U7103 & new_U7104 & new_U7106 & new_U7105;
  assign new_U4072 = new_U7107 & new_U7108 & new_U7110 & new_U7109;
  assign new_U4073 = new_U7111 & new_U7112 & new_U7114 & new_U7113;
  assign new_U4074 = new_U7115 & new_U7116 & new_U7118 & new_U7117;
  assign new_U4075 = new_U7120 & new_U7121 & new_U7123 & new_U7122;
  assign new_U4076 = new_U7124 & new_U7125 & new_U7127 & new_U7126;
  assign new_U4077 = new_U7128 & new_U7129 & new_U7131 & new_U7130;
  assign new_U4078 = new_U7133 & new_U7132;
  assign new_U4079 = new_U4078 & new_U7605 & new_U7134;
  assign new_U4080 = new_U7135 & new_U7136 & new_U7138 & new_U7137;
  assign new_U4081 = new_U7139 & new_U7140 & new_U7142 & new_U7141;
  assign new_U4082 = new_U7143 & new_U7144 & new_U7146 & new_U7145;
  assign new_U4083 = new_U7147 & new_U7148 & new_U7150 & new_U7149;
  assign new_U4084 = new_U7152 & new_U7153 & new_U7155 & new_U7154;
  assign new_U4085 = new_U7156 & new_U7157 & new_U7159 & new_U7158;
  assign new_U4086 = new_U7160 & new_U7161 & new_U7163 & new_U7162;
  assign new_U4087 = new_U7164 & new_U7165 & new_U7167 & new_U7166;
  assign new_U4088 = new_U7169 & new_U7170 & new_U7172 & new_U7171;
  assign new_U4089 = new_U7173 & new_U7174 & new_U7176 & new_U7175;
  assign new_U4090 = new_U7177 & new_U7178 & new_U7180 & new_U7179;
  assign new_U4091 = new_U7181 & new_U7182 & new_U7184 & new_U7183;
  assign new_U4092 = new_U7186 & new_U7187 & new_U7189 & new_U7188;
  assign new_U4093 = new_U7190 & new_U7191 & new_U7193 & new_U7192;
  assign new_U4094 = new_U7194 & new_U7195 & new_U7197 & new_U7196;
  assign new_U4095 = new_U7198 & new_U7199 & new_U7201 & new_U7200;
  assign new_U4096 = new_U7203 & new_U3251;
  assign new_U4097 = new_U7204 & new_U7203;
  assign new_U4098 = new_U7205 & new_U3252;
  assign new_U4099 = new_U7077 & new_U3414;
  assign new_U4100 = new_U7206 & new_U7205;
  assign new_U4101 = new_U7461 & new_U4100 & new_U7460;
  assign new_U4102 = new_U4101 & new_U4099 & new_U7078 & new_U3421;
  assign new_U4103 = new_U7462 & new_U7464 & new_U7474 & new_U7468;
  assign new_U4104 = new_U7475 & new_U7476 & new_U7493 & new_U7477;
  assign new_U4105 = new_U7078 & new_U7077;
  assign new_U4106 = new_U7461 & new_U7460 & new_U3421;
  assign new_U4107 = new_U7462 & new_U7463 & new_U7464;
  assign new_U4108 = new_U4107 & new_U2606 & new_U2608 & new_U7465;
  assign new_U4109 = new_U7208 & new_U7209 & new_U7211 & new_U7210;
  assign new_U4110 = new_U7212 & new_U7213 & new_U7215 & new_U7214;
  assign new_U4111 = new_U7216 & new_U7217 & new_U7219 & new_U7218;
  assign new_U4112 = new_U7220 & new_U7221 & new_U7223 & new_U7222;
  assign new_U4113 = new_U7225 & new_U7226 & new_U7228 & new_U7227;
  assign new_U4114 = new_U7229 & new_U7230 & new_U7232 & new_U7231;
  assign new_U4115 = new_U7233 & new_U7234 & new_U7236 & new_U7235;
  assign new_U4116 = new_U7237 & new_U7238 & new_U7240 & new_U7239;
  assign new_U4117 = new_U7242 & new_U7243 & new_U7245 & new_U7244;
  assign new_U4118 = new_U7246 & new_U7247 & new_U7249 & new_U7248;
  assign new_U4119 = new_U7250 & new_U7251 & new_U7253 & new_U7252;
  assign new_U4120 = new_U7254 & new_U7255 & new_U7257 & new_U7256;
  assign new_U4121 = new_U7259 & new_U7260 & new_U7262 & new_U7261;
  assign new_U4122 = new_U7263 & new_U7264 & new_U7266 & new_U7265;
  assign new_U4123 = new_U7267 & new_U7268 & new_U7270 & new_U7269;
  assign new_U4124 = new_U7271 & new_U7272 & new_U7607 & new_U7273;
  assign new_U4125 = new_U7274 & new_U7275 & new_U7277 & new_U7276;
  assign new_U4126 = new_U7278 & new_U7279 & new_U7281 & new_U7280;
  assign new_U4127 = new_U7282 & new_U7283 & new_U7285 & new_U7284;
  assign new_U4128 = new_U7286 & new_U7287 & new_U7289 & new_U7288;
  assign new_U4129 = new_U7291 & new_U7292 & new_U7294 & new_U7293;
  assign new_U4130 = new_U7295 & new_U7296 & new_U7298 & new_U7297;
  assign new_U4131 = new_U7299 & new_U7300 & new_U7302 & new_U7301;
  assign new_U4132 = new_U7303 & new_U7304 & new_U7306 & new_U7305;
  assign new_U4133 = new_U7308 & new_U7309 & new_U7311 & new_U7310;
  assign new_U4134 = new_U7312 & new_U7313 & new_U7315 & new_U7314;
  assign new_U4135 = new_U7316 & new_U7317 & new_U7319 & new_U7318;
  assign new_U4136 = new_U7320 & new_U7321 & new_U7323 & new_U7322;
  assign new_U4137 = new_U7325 & new_U7326 & new_U7328 & new_U7327;
  assign new_U4138 = new_U7329 & new_U7330 & new_U7332 & new_U7331;
  assign new_U4139 = new_U7333 & new_U7334 & new_U7336 & new_U7335;
  assign new_U4140 = new_U7337 & new_U7338 & new_U7340 & new_U7339;
  assign new_U4141 = new_U3271 & new_U3406;
  assign new_U4142 = new_U3270 & new_U3378;
  assign new_U4143 = new_U4251 & new_U7345 & new_U7346;
  assign new_U4144 = new_U4143 & new_U7347;
  assign new_U4145 = STATE2_REG_0_ & new_U2427;
  assign new_U4146 = new_U4145 & new_U7348;
  assign new_U4147 = new_U3258 & new_U4161;
  assign new_U4148 = STATE2_REG_0_ & new_U4161;
  assign new_U4149 = new_U7357 & STATE2_REG_0_;
  assign new_U4150 = new_U7359 & new_U2603;
  assign new_U4151 = new_U7361 & STATE2_REG_0_;
  assign new_U4152 = new_U7363 & new_U2603;
  assign new_U4153 = new_U7370 & new_U7371;
  assign new_U4154 = new_U3440 & new_U7372;
  assign new_U4155 = new_U7375 & new_U7377 & new_U7376;
  assign new_U4156 = new_U7450 & new_U7449;
  assign new_U4157 = new_U7453 & new_U7452;
  assign new_U4158 = new_U7662 & new_U7661;
  assign new_U4159 = ~new_U3557 | ~new_U3558 | ~new_U3560 | ~new_U3559;
  assign new_U4160 = ~new_U3727 | ~new_U5462;
  assign new_U4161 = ~new_U3561 | ~new_U3562 | ~new_U3563 | ~new_U3564 | ~new_U2607;
  assign new_U4162 = ~INSTADDRPOINTER_REG_31_;
  assign new_U4163 = new_U7714 & new_U7713;
  assign new_U4164 = new_U7733 & new_U7732;
  assign new_U4165 = ~new_U2368 | ~new_U3272;
  assign new_U4166 = ~new_U4496 | ~new_U3378;
  assign new_U4167 = ~BS16_N;
  assign new_U4168 = ~new_U3955 | ~new_U4216;
  assign new_U4169 = ~new_U4216 | ~new_U3419;
  assign new_U4170 = ~new_U3726 | ~new_U7686 | ~new_U7685;
  assign new_U4171 = ~INSTQUEUERD_ADDR_REG_2_ | ~new_U3256;
  assign new_U4172 = ~new_U3439;
  assign new_U4173 = ~HOLD | ~new_U3244;
  assign new_U4174 = ~new_U3399;
  assign new_U4175 = ~new_U3427;
  assign new_U4176 = ~new_U3426;
  assign new_U4177 = ~new_U3380;
  assign new_U4178 = ~new_U3277;
  assign new_U4179 = ~new_U3436;
  assign new_U4180 = ~new_U3392;
  assign new_U4181 = ~new_U3421;
  assign new_U4182 = ~new_U3407;
  assign new_U4183 = ~new_U4253 | ~new_U3258;
  assign new_U4184 = ~new_U4448 | ~new_U2605;
  assign new_U4185 = ~new_U3383;
  assign new_U4186 = ~new_U3412;
  assign new_U4187 = ~new_U3276;
  assign new_U4188 = ~new_U3408;
  assign new_U4189 = ~new_U3409;
  assign new_U4190 = ~new_U3415;
  assign new_U4191 = ~new_U3395;
  assign new_U4192 = ~new_U3414;
  assign new_U4193 = ~new_U4185 | ~new_U3873 | ~new_U4177;
  assign new_U4194 = ~new_U3405;
  assign new_U4195 = ~new_U3430;
  assign new_U4196 = ~new_U3269;
  assign new_U4197 = ~new_U3294;
  assign new_U4198 = ~new_U3377;
  assign new_U4199 = ~new_U3433;
  assign new_U4200 = ~new_U3434;
  assign new_U4201 = ~new_U3435;
  assign new_U4202 = ~new_U3387;
  assign new_U4203 = ~new_U3275;
  assign new_U4204 = ~new_U3279;
  assign new_U4205 = ~new_U3566 | ~new_U2431;
  assign new_U4206 = ~new_U3386;
  assign new_U4207 = ~new_U4437 | ~new_U3258;
  assign new_U4208 = ~new_U3420;
  assign new_U4209 = ~new_U3236;
  assign new_U4210 = ~new_U3413;
  assign new_U4211 = ~new_U3411;
  assign new_U4212 = ~new_U3287;
  assign new_U4213 = ~new_LT_563_1260_U6;
  assign new_U4214 = ~new_U3307;
  assign new_U4215 = ~new_U4243 | ~new_U3418;
  assign new_U4216 = ~new_U4223 | ~new_U7488;
  assign new_U4217 = ~new_U2362 | ~new_U3259;
  assign new_U4218 = ~new_U2363 | ~new_U4365;
  assign new_U4219 = ~new_U3394;
  assign new_U4220 = ~new_U3239;
  assign new_U4221 = ~new_U3237;
  assign new_U4222 = ~new_U3382;
  assign new_U4223 = ~new_U3284;
  assign new_U4224 = ~new_U3385;
  assign new_U4225 = ~new_U4166;
  assign new_U4226 = ~new_U3344;
  assign new_U4227 = ~new_U4465 | ~new_U7369;
  assign new_U4228 = ~new_U3951 | ~new_U4208;
  assign new_U4229 = ~new_U3572 | ~new_U4249;
  assign new_U4230 = ~new_U3719 | ~new_U2428;
  assign new_U4231 = ~new_U4352 | ~new_U3245;
  assign new_U4232 = ~new_U2352 | ~STATE2_REG_1_ | ~new_U3281;
  assign new_U4233 = ~new_U2428 | ~new_U3390;
  assign new_U4234 = ~STATE2_REG_0_ | ~READY_N | ~new_U3250;
  assign new_U4235 = ~new_U3381;
  assign new_U4236 = ~new_U2448 | ~new_U3850 | ~new_U2451 | ~new_U2353;
  assign new_U4237 = ~new_U3274;
  assign new_U4238 = ~new_U3384;
  assign new_U4239 = ~new_U3402;
  assign new_U4240 = ~new_U3286;
  assign new_U4241 = ~new_U3396;
  assign new_U4242 = ~new_U3406;
  assign new_U4243 = ~new_U3419;
  assign new_U4244 = ~new_U3278;
  assign new_U4245 = ~new_U3376;
  assign new_U4246 = ~new_U3241;
  assign new_U4247 = ~new_U3268;
  assign new_U4248 = ~new_U3393;
  assign new_U4249 = ~new_U3285;
  assign new_U4250 = ~new_U3273;
  assign new_U4251 = ~new_U4224 | ~new_U4387;
  assign new_U4252 = ~new_U3398;
  assign new_U4253 = ~new_U3440;
  assign new_U4254 = ~new_U3397;
  assign new_U4255 = ~REIP_REG_31_ | ~new_U4221;
  assign new_U4256 = ~REIP_REG_30_ | ~new_U4220;
  assign new_U4257 = ~ADDRESS_REG_29_ | ~new_U3236;
  assign new_U4258 = ~REIP_REG_30_ | ~new_U4221;
  assign new_U4259 = ~REIP_REG_29_ | ~new_U4220;
  assign new_U4260 = ~ADDRESS_REG_28_ | ~new_U3236;
  assign new_U4261 = ~REIP_REG_29_ | ~new_U4221;
  assign new_U4262 = ~REIP_REG_28_ | ~new_U4220;
  assign new_U4263 = ~ADDRESS_REG_27_ | ~new_U3236;
  assign new_U4264 = ~REIP_REG_28_ | ~new_U4221;
  assign new_U4265 = ~REIP_REG_27_ | ~new_U4220;
  assign new_U4266 = ~ADDRESS_REG_26_ | ~new_U3236;
  assign new_U4267 = ~REIP_REG_27_ | ~new_U4221;
  assign new_U4268 = ~REIP_REG_26_ | ~new_U4220;
  assign new_U4269 = ~ADDRESS_REG_25_ | ~new_U3236;
  assign new_U4270 = ~REIP_REG_26_ | ~new_U4221;
  assign new_U4271 = ~REIP_REG_25_ | ~new_U4220;
  assign new_U4272 = ~ADDRESS_REG_24_ | ~new_U3236;
  assign new_U4273 = ~REIP_REG_25_ | ~new_U4221;
  assign new_U4274 = ~REIP_REG_24_ | ~new_U4220;
  assign new_U4275 = ~ADDRESS_REG_23_ | ~new_U3236;
  assign new_U4276 = ~REIP_REG_24_ | ~new_U4221;
  assign new_U4277 = ~REIP_REG_23_ | ~new_U4220;
  assign new_U4278 = ~ADDRESS_REG_22_ | ~new_U3236;
  assign new_U4279 = ~REIP_REG_23_ | ~new_U4221;
  assign new_U4280 = ~REIP_REG_22_ | ~new_U4220;
  assign new_U4281 = ~ADDRESS_REG_21_ | ~new_U3236;
  assign new_U4282 = ~REIP_REG_22_ | ~new_U4221;
  assign new_U4283 = ~REIP_REG_21_ | ~new_U4220;
  assign new_U4284 = ~ADDRESS_REG_20_ | ~new_U3236;
  assign new_U4285 = ~REIP_REG_21_ | ~new_U4221;
  assign new_U4286 = ~REIP_REG_20_ | ~new_U4220;
  assign new_U4287 = ~ADDRESS_REG_19_ | ~new_U3236;
  assign new_U4288 = ~REIP_REG_20_ | ~new_U4221;
  assign new_U4289 = ~REIP_REG_19_ | ~new_U4220;
  assign new_U4290 = ~ADDRESS_REG_18_ | ~new_U3236;
  assign new_U4291 = ~REIP_REG_19_ | ~new_U4221;
  assign new_U4292 = ~REIP_REG_18_ | ~new_U4220;
  assign new_U4293 = ~ADDRESS_REG_17_ | ~new_U3236;
  assign new_U4294 = ~REIP_REG_18_ | ~new_U4221;
  assign new_U4295 = ~REIP_REG_17_ | ~new_U4220;
  assign new_U4296 = ~ADDRESS_REG_16_ | ~new_U3236;
  assign new_U4297 = ~REIP_REG_17_ | ~new_U4221;
  assign new_U4298 = ~REIP_REG_16_ | ~new_U4220;
  assign new_U4299 = ~ADDRESS_REG_15_ | ~new_U3236;
  assign new_U4300 = ~REIP_REG_16_ | ~new_U4221;
  assign new_U4301 = ~REIP_REG_15_ | ~new_U4220;
  assign new_U4302 = ~ADDRESS_REG_14_ | ~new_U3236;
  assign new_U4303 = ~REIP_REG_15_ | ~new_U4221;
  assign new_U4304 = ~REIP_REG_14_ | ~new_U4220;
  assign new_U4305 = ~ADDRESS_REG_13_ | ~new_U3236;
  assign new_U4306 = ~REIP_REG_14_ | ~new_U4221;
  assign new_U4307 = ~REIP_REG_13_ | ~new_U4220;
  assign new_U4308 = ~ADDRESS_REG_12_ | ~new_U3236;
  assign new_U4309 = ~REIP_REG_13_ | ~new_U4221;
  assign new_U4310 = ~REIP_REG_12_ | ~new_U4220;
  assign new_U4311 = ~ADDRESS_REG_11_ | ~new_U3236;
  assign new_U4312 = ~REIP_REG_12_ | ~new_U4221;
  assign new_U4313 = ~REIP_REG_11_ | ~new_U4220;
  assign new_U4314 = ~ADDRESS_REG_10_ | ~new_U3236;
  assign new_U4315 = ~REIP_REG_11_ | ~new_U4221;
  assign new_U4316 = ~REIP_REG_10_ | ~new_U4220;
  assign new_U4317 = ~ADDRESS_REG_9_ | ~new_U3236;
  assign new_U4318 = ~REIP_REG_10_ | ~new_U4221;
  assign new_U4319 = ~REIP_REG_9_ | ~new_U4220;
  assign new_U4320 = ~ADDRESS_REG_8_ | ~new_U3236;
  assign new_U4321 = ~REIP_REG_9_ | ~new_U4221;
  assign new_U4322 = ~REIP_REG_8_ | ~new_U4220;
  assign new_U4323 = ~ADDRESS_REG_7_ | ~new_U3236;
  assign new_U4324 = ~REIP_REG_8_ | ~new_U4221;
  assign new_U4325 = ~REIP_REG_7_ | ~new_U4220;
  assign new_U4326 = ~ADDRESS_REG_6_ | ~new_U3236;
  assign new_U4327 = ~REIP_REG_7_ | ~new_U4221;
  assign new_U4328 = ~REIP_REG_6_ | ~new_U4220;
  assign new_U4329 = ~ADDRESS_REG_5_ | ~new_U3236;
  assign new_U4330 = ~REIP_REG_6_ | ~new_U4221;
  assign new_U4331 = ~REIP_REG_5_ | ~new_U4220;
  assign new_U4332 = ~ADDRESS_REG_4_ | ~new_U3236;
  assign new_U4333 = ~REIP_REG_5_ | ~new_U4221;
  assign new_U4334 = ~REIP_REG_4_ | ~new_U4220;
  assign new_U4335 = ~ADDRESS_REG_3_ | ~new_U3236;
  assign new_U4336 = ~REIP_REG_4_ | ~new_U4221;
  assign new_U4337 = ~REIP_REG_3_ | ~new_U4220;
  assign new_U4338 = ~ADDRESS_REG_2_ | ~new_U3236;
  assign new_U4339 = ~REIP_REG_3_ | ~new_U4221;
  assign new_U4340 = ~REIP_REG_2_ | ~new_U4220;
  assign new_U4341 = ~ADDRESS_REG_1_ | ~new_U3236;
  assign new_U4342 = ~REIP_REG_2_ | ~new_U4221;
  assign new_U4343 = ~REIP_REG_1_ | ~new_U4220;
  assign new_U4344 = ~ADDRESS_REG_0_ | ~new_U3236;
  assign new_U4345 = ~new_U3247;
  assign new_U4346 = ~new_U4345 | ~new_U3244;
  assign new_U4347 = ~NA_N | ~new_U4246;
  assign new_U4348 = ~new_U3248;
  assign new_U4349 = ~new_U4348 | ~new_U3244;
  assign new_U4350 = STATE_REG_0_ | NA_N;
  assign new_U4351 = ~new_U7611 | ~new_U7610 | ~new_U4350;
  assign new_U4352 = ~new_U3242;
  assign new_U4353 = ~new_U4352 | ~HOLD | ~new_U3234;
  assign new_U4354 = ~new_U3481 | ~new_U3248;
  assign new_U4355 = ~new_U4354 | ~new_U4353;
  assign new_U4356 = ~new_U4355 | ~STATE_REG_0_ | ~new_U4347;
  assign new_U4357 = ~STATE_REG_2_ | ~new_U4351;
  assign new_U4358 = ~READY_N | ~new_U4209;
  assign new_U4359 = ~new_U3484 | ~new_U7613;
  assign new_U4360 = ~STATE_REG_2_ | ~new_U3247;
  assign new_U4361 = ~NA_N | ~new_U3245;
  assign new_U4362 = ~new_U4361 | ~new_U4360;
  assign new_U4363 = ~new_U4362 | ~new_U3235;
  assign new_U4364 = ~new_U4167 | ~new_U3242;
  assign new_U4365 = ~new_U3267;
  assign new_U4366 = ~new_U3256;
  assign new_U4367 = ~new_U3431;
  assign new_U4368 = ~new_U3255;
  assign new_U4369 = ~new_U3261;
  assign new_U4370 = ~new_U3254;
  assign new_U4371 = ~INSTQUEUE_REG_7__3_ | ~new_U4370;
  assign new_U4372 = ~INSTQUEUE_REG_0__3_ | ~new_U2472;
  assign new_U4373 = ~INSTQUEUE_REG_1__3_ | ~new_U2471;
  assign new_U4374 = ~INSTQUEUE_REG_2__3_ | ~new_U2470;
  assign new_U4375 = ~INSTQUEUE_REG_3__3_ | ~new_U2468;
  assign new_U4376 = ~INSTQUEUE_REG_4__3_ | ~new_U2467;
  assign new_U4377 = ~INSTQUEUE_REG_5__3_ | ~new_U2466;
  assign new_U4378 = ~INSTQUEUE_REG_6__3_ | ~new_U2465;
  assign new_U4379 = ~INSTQUEUE_REG_8__3_ | ~new_U2464;
  assign new_U4380 = ~INSTQUEUE_REG_9__3_ | ~new_U2463;
  assign new_U4381 = ~INSTQUEUE_REG_10__3_ | ~new_U2461;
  assign new_U4382 = ~INSTQUEUE_REG_11__3_ | ~new_U2459;
  assign new_U4383 = ~INSTQUEUE_REG_12__3_ | ~new_U2458;
  assign new_U4384 = ~INSTQUEUE_REG_13__3_ | ~new_U2457;
  assign new_U4385 = ~INSTQUEUE_REG_14__3_ | ~new_U2455;
  assign new_U4386 = ~INSTQUEUE_REG_15__3_ | ~new_U2453;
  assign new_U4387 = ~new_U3270;
  assign new_U4388 = ~new_U3265;
  assign new_U4389 = ~INSTQUEUERD_ADDR_REG_0_ | ~INSTQUEUE_REG_7__5_ | ~INSTQUEUERD_ADDR_REG_1_ | ~INSTQUEUERD_ADDR_REG_2_ | ~new_U3257;
  assign new_U4390 = ~new_U4368 | ~INSTQUEUE_REG_0__5_ | ~new_U3257;
  assign new_U4391 = ~new_U3252 | ~INSTQUEUERD_ADDR_REG_0_ | ~INSTQUEUE_REG_1__5_ | ~new_U2469;
  assign new_U4392 = ~new_U3253 | ~INSTQUEUERD_ADDR_REG_1_ | ~INSTQUEUE_REG_2__5_ | ~new_U2469;
  assign new_U4393 = ~new_U3257 | ~INSTQUEUERD_ADDR_REG_2_ | ~INSTQUEUE_REG_4__5_ | ~new_U4366;
  assign new_U4394 = ~new_U3509 | ~new_U3508 | ~INSTQUEUERD_ADDR_REG_2_;
  assign new_U4395 = ~new_U3511 | ~new_U3510 | ~INSTQUEUERD_ADDR_REG_2_;
  assign new_U4396 = ~new_U3512 | ~new_U4368;
  assign new_U4397 = ~new_U3514 | ~new_U3513 | ~INSTQUEUERD_ADDR_REG_1_;
  assign new_U4398 = ~INSTQUEUERD_ADDR_REG_3_ | ~INSTQUEUE_REG_11__5_ | ~INSTQUEUERD_ADDR_REG_0_ | ~INSTQUEUERD_ADDR_REG_1_ | ~new_U3251;
  assign new_U4399 = ~new_U3515 | ~new_U4366 | ~INSTQUEUERD_ADDR_REG_2_;
  assign new_U4400 = ~INSTQUEUERD_ADDR_REG_3_ | ~INSTQUEUE_REG_13__5_ | ~INSTQUEUERD_ADDR_REG_0_ | ~INSTQUEUERD_ADDR_REG_2_ | ~new_U3252;
  assign new_U4401 = ~INSTQUEUERD_ADDR_REG_3_ | ~INSTQUEUE_REG_14__5_ | ~INSTQUEUERD_ADDR_REG_1_ | ~INSTQUEUERD_ADDR_REG_2_ | ~new_U3253;
  assign new_U4402 = ~INSTQUEUERD_ADDR_REG_3_ | ~INSTQUEUE_REG_15__5_ | ~INSTQUEUERD_ADDR_REG_0_ | ~INSTQUEUERD_ADDR_REG_1_ | ~INSTQUEUERD_ADDR_REG_2_;
  assign new_U4403 = ~new_U4161;
  assign new_U4404 = ~INSTQUEUE_REG_7__2_ | ~new_U4370;
  assign new_U4405 = ~INSTQUEUE_REG_0__2_ | ~new_U2472;
  assign new_U4406 = ~INSTQUEUE_REG_1__2_ | ~new_U2471;
  assign new_U4407 = ~INSTQUEUE_REG_2__2_ | ~new_U2470;
  assign new_U4408 = ~INSTQUEUE_REG_3__2_ | ~new_U2468;
  assign new_U4409 = ~INSTQUEUE_REG_4__2_ | ~new_U2467;
  assign new_U4410 = ~INSTQUEUE_REG_5__2_ | ~new_U2466;
  assign new_U4411 = ~INSTQUEUE_REG_6__2_ | ~new_U2465;
  assign new_U4412 = ~INSTQUEUE_REG_8__2_ | ~new_U2464;
  assign new_U4413 = ~INSTQUEUE_REG_9__2_ | ~new_U2463;
  assign new_U4414 = ~INSTQUEUE_REG_10__2_ | ~new_U2461;
  assign new_U4415 = ~INSTQUEUE_REG_11__2_ | ~new_U2459;
  assign new_U4416 = ~INSTQUEUE_REG_12__2_ | ~new_U2458;
  assign new_U4417 = ~INSTQUEUE_REG_13__2_ | ~new_U2457;
  assign new_U4418 = ~INSTQUEUE_REG_14__2_ | ~new_U2455;
  assign new_U4419 = ~INSTQUEUE_REG_15__2_ | ~new_U2453;
  assign new_U4420 = ~new_U4159;
  assign new_U4421 = ~INSTQUEUE_REG_7__7_ | ~new_U4370;
  assign new_U4422 = ~INSTQUEUE_REG_0__7_ | ~new_U2472;
  assign new_U4423 = ~INSTQUEUE_REG_1__7_ | ~new_U2471;
  assign new_U4424 = ~INSTQUEUE_REG_2__7_ | ~new_U2470;
  assign new_U4425 = ~INSTQUEUE_REG_3__7_ | ~new_U2468;
  assign new_U4426 = ~INSTQUEUE_REG_4__7_ | ~new_U2467;
  assign new_U4427 = ~INSTQUEUE_REG_5__7_ | ~new_U2466;
  assign new_U4428 = ~INSTQUEUE_REG_6__7_ | ~new_U2465;
  assign new_U4429 = ~INSTQUEUE_REG_8__7_ | ~new_U2464;
  assign new_U4430 = ~INSTQUEUE_REG_9__7_ | ~new_U2463;
  assign new_U4431 = ~INSTQUEUE_REG_10__7_ | ~new_U2461;
  assign new_U4432 = ~INSTQUEUE_REG_11__7_ | ~new_U2459;
  assign new_U4433 = ~INSTQUEUE_REG_12__7_ | ~new_U2458;
  assign new_U4434 = ~INSTQUEUE_REG_13__7_ | ~new_U2457;
  assign new_U4435 = ~INSTQUEUE_REG_14__7_ | ~new_U2455;
  assign new_U4436 = ~INSTQUEUE_REG_15__7_ | ~new_U2453;
  assign new_U4437 = ~new_U3378;
  assign new_U4438 = ~INSTQUEUE_REG_7__6_ | ~new_U3486 | ~new_U4369;
  assign new_U4439 = ~new_U2456 | ~INSTQUEUE_REG_1__6_ | ~new_U2469;
  assign new_U4440 = ~new_U2454 | ~INSTQUEUE_REG_2__6_ | ~new_U2469;
  assign new_U4441 = ~new_U4369 | ~INSTQUEUE_REG_4__6_ | ~new_U4366;
  assign new_U4442 = ~INSTQUEUE_REG_5__6_ | ~new_U2456 | ~new_U4369;
  assign new_U4443 = ~INSTQUEUE_REG_6__6_ | ~new_U2454 | ~new_U4369;
  assign new_U4444 = ~new_U3495 | ~INSTQUEUE_REG_12__6_ | ~new_U4366;
  assign new_U4445 = ~INSTQUEUE_REG_13__6_ | ~new_U3495 | ~new_U2456;
  assign new_U4446 = ~INSTQUEUE_REG_14__6_ | ~new_U3495 | ~new_U2454;
  assign new_U4447 = ~INSTQUEUE_REG_15__6_ | ~new_U3495 | ~new_U3486;
  assign new_U4448 = ~new_U3264;
  assign new_U4449 = ~INSTQUEUE_REG_7__1_ | ~new_U4370;
  assign new_U4450 = ~INSTQUEUE_REG_0__1_ | ~new_U2472;
  assign new_U4451 = ~INSTQUEUE_REG_1__1_ | ~new_U2471;
  assign new_U4452 = ~INSTQUEUE_REG_2__1_ | ~new_U2470;
  assign new_U4453 = ~INSTQUEUE_REG_3__1_ | ~new_U2468;
  assign new_U4454 = ~INSTQUEUE_REG_4__1_ | ~new_U2467;
  assign new_U4455 = ~INSTQUEUE_REG_5__1_ | ~new_U2466;
  assign new_U4456 = ~INSTQUEUE_REG_6__1_ | ~new_U2465;
  assign new_U4457 = ~INSTQUEUE_REG_8__1_ | ~new_U2464;
  assign new_U4458 = ~INSTQUEUE_REG_9__1_ | ~new_U2463;
  assign new_U4459 = ~INSTQUEUE_REG_10__1_ | ~new_U2461;
  assign new_U4460 = ~INSTQUEUE_REG_11__1_ | ~new_U2459;
  assign new_U4461 = ~INSTQUEUE_REG_12__1_ | ~new_U2458;
  assign new_U4462 = ~INSTQUEUE_REG_13__1_ | ~new_U2457;
  assign new_U4463 = ~INSTQUEUE_REG_14__1_ | ~new_U2455;
  assign new_U4464 = ~INSTQUEUE_REG_15__1_ | ~new_U2453;
  assign new_U4465 = ~new_U3258;
  assign new_U4466 = ~INSTQUEUE_REG_7__0_ | ~new_U4370;
  assign new_U4467 = ~INSTQUEUE_REG_0__0_ | ~new_U2472;
  assign new_U4468 = ~INSTQUEUE_REG_1__0_ | ~new_U2471;
  assign new_U4469 = ~INSTQUEUE_REG_2__0_ | ~new_U2470;
  assign new_U4470 = ~INSTQUEUE_REG_3__0_ | ~new_U2468;
  assign new_U4471 = ~INSTQUEUE_REG_4__0_ | ~new_U2467;
  assign new_U4472 = ~INSTQUEUE_REG_5__0_ | ~new_U2466;
  assign new_U4473 = ~INSTQUEUE_REG_6__0_ | ~new_U2465;
  assign new_U4474 = ~INSTQUEUE_REG_8__0_ | ~new_U2464;
  assign new_U4475 = ~INSTQUEUE_REG_9__0_ | ~new_U2463;
  assign new_U4476 = ~INSTQUEUE_REG_10__0_ | ~new_U2461;
  assign new_U4477 = ~INSTQUEUE_REG_11__0_ | ~new_U2459;
  assign new_U4478 = ~INSTQUEUE_REG_12__0_ | ~new_U2458;
  assign new_U4479 = ~INSTQUEUE_REG_13__0_ | ~new_U2457;
  assign new_U4480 = ~INSTQUEUE_REG_14__0_ | ~new_U2455;
  assign new_U4481 = ~INSTQUEUE_REG_15__0_ | ~new_U2453;
  assign new_U4482 = ~new_U3271;
  assign new_U4483 = ~STATE_REG_2_ | ~new_U3235;
  assign new_U4484 = ~new_U3241 | ~new_U4483;
  assign new_U4485 = ~new_U3259;
  assign new_U4486 = ~new_U4465 | ~new_U3375;
  assign new_U4487 = ~new_U3424;
  assign new_U4488 = ~new_U3274 | ~new_U3259 | ~new_U3377;
  assign new_U4489 = ~new_U4488 | ~new_U3244;
  assign new_U4490 = ~new_U3272;
  assign new_U4491 = ~new_U4448 | ~new_U4161;
  assign new_U4492 = ~new_U4184 | ~new_U3273;
  assign new_U4493 = ~new_U4492 | ~new_U3567;
  assign new_U4494 = ~new_U3568 | ~new_U4493;
  assign new_U4495 = ~new_U4203 | ~new_U3375;
  assign new_U4496 = ~new_U4495 | ~new_U7670 | ~new_U7669;
  assign new_U4497 = ~new_U2448 | ~new_U4250;
  assign new_U4498 = MORE_REG | FLUSH_REG;
  assign new_U4499 = ~new_U3280;
  assign new_U4500 = ~new_U4499 | ~new_U3249;
  assign new_U4501 = ~STATE2_REG_1_ | ~READY_N;
  assign new_U4502 = ~new_U3282;
  assign new_U4503 = ~STATE2_REG_1_ | ~new_U7676 | ~new_U7675;
  assign new_U4504 = ~STATE2_REG_2_ | ~new_U3282;
  assign new_U4505 = ~new_U7592 | ~new_U4234;
  assign new_U4506 = ~new_U3571 | ~new_U4502;
  assign new_U4507 = ~STATE2_REG_1_ | ~new_U4505;
  assign new_U4508 = ~new_U2368 | ~new_U7592;
  assign new_U4509 = ~new_U4240 | ~new_U4249;
  assign new_U4510 = ~new_U7592 | ~new_U4233;
  assign new_U4511 = ~new_U2368 | ~new_U3280;
  assign new_U4512 = ~new_U3312;
  assign new_U4513 = ~new_U3318;
  assign new_U4514 = ~new_U3319;
  assign new_U4515 = ~new_U3301;
  assign new_U4516 = ~new_U3300;
  assign new_U4517 = ~new_U3329;
  assign new_U4518 = ~new_R2144_U8 | ~new_U3300;
  assign new_U4519 = ~new_U3345;
  assign new_U4520 = ~new_U3302;
  assign new_U4521 = ~new_U3292;
  assign new_U4522 = ~new_U3293;
  assign new_U4523 = ~new_U2438 | ~new_U2442;
  assign new_U4524 = ~new_U3308;
  assign new_U4525 = ~new_U3343;
  assign new_U4526 = ~new_U3327;
  assign new_U4527 = ~INSTQUEUEWR_ADDR_REG_3_ | ~new_U3292;
  assign new_U4528 = ~new_U3347;
  assign new_U4529 = ~new_U3316;
  assign new_U4530 = ~new_U3310;
  assign new_U4531 = ~new_U3222;
  assign new_U4532 = ~new_U2432 | ~new_U2436;
  assign new_U4533 = ~new_U3309;
  assign new_U4534 = ~STATE2_REG_1_ | ~new_U3250;
  assign new_U4535 = ~new_U3286 | ~new_U4534 | ~new_U3284;
  assign new_U4536 = ~new_U4516 | ~new_U2476;
  assign new_U4537 = ~new_U2480 | ~new_U2358;
  assign new_U4538 = ~new_U3307 | ~new_U4537;
  assign new_U4539 = ~new_U4524 | ~new_U4538;
  assign new_U4540 = ~STATE2_REG_3_ | ~new_U3293;
  assign new_U4541 = ~new_U4533 | ~STATE2_REG_2_;
  assign new_U4542 = ~new_U4539 | ~new_U3575;
  assign new_U4543 = ~new_U2480 | ~new_U2388;
  assign new_U4544 = ~new_U3307 | ~new_U4543;
  assign new_U4545 = ~new_U4544 | ~new_U3308;
  assign new_U4546 = ~STATE2_REG_2_ | ~new_U3309;
  assign new_U4547 = ~new_U4546 | ~new_U4545;
  assign new_U4548 = ~new_U2415 | ~new_U4522;
  assign new_U4549 = ~new_U2413 | ~new_U2477;
  assign new_U4550 = ~new_U2412 | ~new_U4520;
  assign new_U4551 = ~new_U2397 | ~new_U4547;
  assign new_U4552 = ~INSTQUEUE_REG_15__7_ | ~new_U4542;
  assign new_U4553 = ~new_U2416 | ~new_U4522;
  assign new_U4554 = ~new_U2411 | ~new_U2477;
  assign new_U4555 = ~new_U2410 | ~new_U4520;
  assign new_U4556 = ~new_U2396 | ~new_U4547;
  assign new_U4557 = ~INSTQUEUE_REG_15__6_ | ~new_U4542;
  assign new_U4558 = ~new_U2420 | ~new_U4522;
  assign new_U4559 = ~new_U2409 | ~new_U2477;
  assign new_U4560 = ~new_U2408 | ~new_U4520;
  assign new_U4561 = ~new_U2395 | ~new_U4547;
  assign new_U4562 = ~INSTQUEUE_REG_15__5_ | ~new_U4542;
  assign new_U4563 = ~new_U2419 | ~new_U4522;
  assign new_U4564 = ~new_U2407 | ~new_U2477;
  assign new_U4565 = ~new_U2406 | ~new_U4520;
  assign new_U4566 = ~new_U2394 | ~new_U4547;
  assign new_U4567 = ~INSTQUEUE_REG_15__4_ | ~new_U4542;
  assign new_U4568 = ~new_U2418 | ~new_U4522;
  assign new_U4569 = ~new_U2405 | ~new_U2477;
  assign new_U4570 = ~new_U2404 | ~new_U4520;
  assign new_U4571 = ~new_U2393 | ~new_U4547;
  assign new_U4572 = ~INSTQUEUE_REG_15__3_ | ~new_U4542;
  assign new_U4573 = ~new_U2421 | ~new_U4522;
  assign new_U4574 = ~new_U2403 | ~new_U2477;
  assign new_U4575 = ~new_U2402 | ~new_U4520;
  assign new_U4576 = ~new_U2392 | ~new_U4547;
  assign new_U4577 = ~INSTQUEUE_REG_15__2_ | ~new_U4542;
  assign new_U4578 = ~new_U2414 | ~new_U4522;
  assign new_U4579 = ~new_U2401 | ~new_U2477;
  assign new_U4580 = ~new_U2400 | ~new_U4520;
  assign new_U4581 = ~new_U2391 | ~new_U4547;
  assign new_U4582 = ~INSTQUEUE_REG_15__1_ | ~new_U4542;
  assign new_U4583 = ~new_U2417 | ~new_U4522;
  assign new_U4584 = ~new_U2399 | ~new_U2477;
  assign new_U4585 = ~new_U2398 | ~new_U4520;
  assign new_U4586 = ~new_U2390 | ~new_U4547;
  assign new_U4587 = ~INSTQUEUE_REG_15__0_ | ~new_U4542;
  assign new_U4588 = ~new_U3313;
  assign new_U4589 = ~new_U3314;
  assign new_U4590 = ~new_U3311;
  assign new_U4591 = ~new_U2443 | ~new_U2438;
  assign new_U4592 = ~new_U3315;
  assign new_U4593 = ~new_U3223;
  assign new_U4594 = ~new_U4512 | ~new_U2476;
  assign new_U4595 = ~new_U2482 | ~new_U2358;
  assign new_U4596 = ~new_U3307 | ~new_U4595;
  assign new_U4597 = ~new_U4592 | ~new_U4596;
  assign new_U4598 = ~STATE2_REG_3_ | ~new_U3311;
  assign new_U4599 = ~STATE2_REG_2_ | ~new_U3223;
  assign new_U4600 = ~new_U4597 | ~new_U3584;
  assign new_U4601 = ~new_U2482 | ~new_U2388;
  assign new_U4602 = ~new_U3307 | ~new_U4601;
  assign new_U4603 = ~new_U4602 | ~new_U3315;
  assign new_U4604 = ~STATE2_REG_2_ | ~new_U4593;
  assign new_U4605 = ~new_U4604 | ~new_U4603;
  assign new_U4606 = ~new_U4590 | ~new_U2415;
  assign new_U4607 = ~new_U2481 | ~new_U2413;
  assign new_U4608 = ~new_U4589 | ~new_U2412;
  assign new_U4609 = ~new_U2397 | ~new_U4605;
  assign new_U4610 = ~INSTQUEUE_REG_14__7_ | ~new_U4600;
  assign new_U4611 = ~new_U4590 | ~new_U2416;
  assign new_U4612 = ~new_U2481 | ~new_U2411;
  assign new_U4613 = ~new_U4589 | ~new_U2410;
  assign new_U4614 = ~new_U2396 | ~new_U4605;
  assign new_U4615 = ~INSTQUEUE_REG_14__6_ | ~new_U4600;
  assign new_U4616 = ~new_U4590 | ~new_U2420;
  assign new_U4617 = ~new_U2481 | ~new_U2409;
  assign new_U4618 = ~new_U4589 | ~new_U2408;
  assign new_U4619 = ~new_U2395 | ~new_U4605;
  assign new_U4620 = ~INSTQUEUE_REG_14__5_ | ~new_U4600;
  assign new_U4621 = ~new_U4590 | ~new_U2419;
  assign new_U4622 = ~new_U2481 | ~new_U2407;
  assign new_U4623 = ~new_U4589 | ~new_U2406;
  assign new_U4624 = ~new_U2394 | ~new_U4605;
  assign new_U4625 = ~INSTQUEUE_REG_14__4_ | ~new_U4600;
  assign new_U4626 = ~new_U4590 | ~new_U2418;
  assign new_U4627 = ~new_U2481 | ~new_U2405;
  assign new_U4628 = ~new_U4589 | ~new_U2404;
  assign new_U4629 = ~new_U2393 | ~new_U4605;
  assign new_U4630 = ~INSTQUEUE_REG_14__3_ | ~new_U4600;
  assign new_U4631 = ~new_U4590 | ~new_U2421;
  assign new_U4632 = ~new_U2481 | ~new_U2403;
  assign new_U4633 = ~new_U4589 | ~new_U2402;
  assign new_U4634 = ~new_U2392 | ~new_U4605;
  assign new_U4635 = ~INSTQUEUE_REG_14__2_ | ~new_U4600;
  assign new_U4636 = ~new_U4590 | ~new_U2414;
  assign new_U4637 = ~new_U2481 | ~new_U2401;
  assign new_U4638 = ~new_U4589 | ~new_U2400;
  assign new_U4639 = ~new_U2391 | ~new_U4605;
  assign new_U4640 = ~INSTQUEUE_REG_14__1_ | ~new_U4600;
  assign new_U4641 = ~new_U4590 | ~new_U2417;
  assign new_U4642 = ~new_U2481 | ~new_U2399;
  assign new_U4643 = ~new_U4589 | ~new_U2398;
  assign new_U4644 = ~new_U2390 | ~new_U4605;
  assign new_U4645 = ~INSTQUEUE_REG_14__0_ | ~new_U4600;
  assign new_U4646 = ~new_U3320;
  assign new_U4647 = ~new_U3321;
  assign new_U4648 = ~new_U3317;
  assign new_U4649 = ~new_U2444 | ~new_U2438;
  assign new_U4650 = ~new_U3322;
  assign new_U4651 = ~new_U2437 | ~new_U2432;
  assign new_U4652 = ~new_U3323;
  assign new_U4653 = ~new_U4513 | ~new_U2476;
  assign new_U4654 = ~new_U2484 | ~new_U2358;
  assign new_U4655 = ~new_U3307 | ~new_U4654;
  assign new_U4656 = ~new_U4650 | ~new_U4655;
  assign new_U4657 = ~STATE2_REG_3_ | ~new_U3317;
  assign new_U4658 = ~new_U4652 | ~STATE2_REG_2_;
  assign new_U4659 = ~new_U4656 | ~new_U3593;
  assign new_U4660 = ~new_U2484 | ~new_U2388;
  assign new_U4661 = ~new_U3307 | ~new_U4660;
  assign new_U4662 = ~new_U4661 | ~new_U3322;
  assign new_U4663 = ~STATE2_REG_2_ | ~new_U3323;
  assign new_U4664 = ~new_U4663 | ~new_U4662;
  assign new_U4665 = ~new_U4648 | ~new_U2415;
  assign new_U4666 = ~new_U2483 | ~new_U2413;
  assign new_U4667 = ~new_U4647 | ~new_U2412;
  assign new_U4668 = ~new_U2397 | ~new_U4664;
  assign new_U4669 = ~INSTQUEUE_REG_13__7_ | ~new_U4659;
  assign new_U4670 = ~new_U4648 | ~new_U2416;
  assign new_U4671 = ~new_U2483 | ~new_U2411;
  assign new_U4672 = ~new_U4647 | ~new_U2410;
  assign new_U4673 = ~new_U2396 | ~new_U4664;
  assign new_U4674 = ~INSTQUEUE_REG_13__6_ | ~new_U4659;
  assign new_U4675 = ~new_U4648 | ~new_U2420;
  assign new_U4676 = ~new_U2483 | ~new_U2409;
  assign new_U4677 = ~new_U4647 | ~new_U2408;
  assign new_U4678 = ~new_U2395 | ~new_U4664;
  assign new_U4679 = ~INSTQUEUE_REG_13__5_ | ~new_U4659;
  assign new_U4680 = ~new_U4648 | ~new_U2419;
  assign new_U4681 = ~new_U2483 | ~new_U2407;
  assign new_U4682 = ~new_U4647 | ~new_U2406;
  assign new_U4683 = ~new_U2394 | ~new_U4664;
  assign new_U4684 = ~INSTQUEUE_REG_13__4_ | ~new_U4659;
  assign new_U4685 = ~new_U4648 | ~new_U2418;
  assign new_U4686 = ~new_U2483 | ~new_U2405;
  assign new_U4687 = ~new_U4647 | ~new_U2404;
  assign new_U4688 = ~new_U2393 | ~new_U4664;
  assign new_U4689 = ~INSTQUEUE_REG_13__3_ | ~new_U4659;
  assign new_U4690 = ~new_U4648 | ~new_U2421;
  assign new_U4691 = ~new_U2483 | ~new_U2403;
  assign new_U4692 = ~new_U4647 | ~new_U2402;
  assign new_U4693 = ~new_U2392 | ~new_U4664;
  assign new_U4694 = ~INSTQUEUE_REG_13__2_ | ~new_U4659;
  assign new_U4695 = ~new_U4648 | ~new_U2414;
  assign new_U4696 = ~new_U2483 | ~new_U2401;
  assign new_U4697 = ~new_U4647 | ~new_U2400;
  assign new_U4698 = ~new_U2391 | ~new_U4664;
  assign new_U4699 = ~INSTQUEUE_REG_13__1_ | ~new_U4659;
  assign new_U4700 = ~new_U4648 | ~new_U2417;
  assign new_U4701 = ~new_U2483 | ~new_U2399;
  assign new_U4702 = ~new_U4647 | ~new_U2398;
  assign new_U4703 = ~new_U2390 | ~new_U4664;
  assign new_U4704 = ~INSTQUEUE_REG_13__0_ | ~new_U4659;
  assign new_U4705 = ~new_U3325;
  assign new_U4706 = ~new_U3324;
  assign new_U4707 = ~new_U2445 | ~new_U2438;
  assign new_U4708 = ~new_U3326;
  assign new_U4709 = ~new_U3224;
  assign new_U4710 = ~new_U2486 | ~new_U2476;
  assign new_U4711 = ~new_U2489 | ~new_U2358;
  assign new_U4712 = ~new_U3307 | ~new_U4711;
  assign new_U4713 = ~new_U4708 | ~new_U4712;
  assign new_U4714 = ~STATE2_REG_3_ | ~new_U3324;
  assign new_U4715 = ~STATE2_REG_2_ | ~new_U3224;
  assign new_U4716 = ~new_U4713 | ~new_U3602;
  assign new_U4717 = ~new_U2489 | ~new_U2388;
  assign new_U4718 = ~new_U3307 | ~new_U4717;
  assign new_U4719 = ~new_U4718 | ~new_U3326;
  assign new_U4720 = ~STATE2_REG_2_ | ~new_U4709;
  assign new_U4721 = ~new_U4720 | ~new_U4719;
  assign new_U4722 = ~new_U4706 | ~new_U2415;
  assign new_U4723 = ~new_U2487 | ~new_U2413;
  assign new_U4724 = ~new_U4705 | ~new_U2412;
  assign new_U4725 = ~new_U2397 | ~new_U4721;
  assign new_U4726 = ~INSTQUEUE_REG_12__7_ | ~new_U4716;
  assign new_U4727 = ~new_U4706 | ~new_U2416;
  assign new_U4728 = ~new_U2487 | ~new_U2411;
  assign new_U4729 = ~new_U4705 | ~new_U2410;
  assign new_U4730 = ~new_U2396 | ~new_U4721;
  assign new_U4731 = ~INSTQUEUE_REG_12__6_ | ~new_U4716;
  assign new_U4732 = ~new_U4706 | ~new_U2420;
  assign new_U4733 = ~new_U2487 | ~new_U2409;
  assign new_U4734 = ~new_U4705 | ~new_U2408;
  assign new_U4735 = ~new_U2395 | ~new_U4721;
  assign new_U4736 = ~INSTQUEUE_REG_12__5_ | ~new_U4716;
  assign new_U4737 = ~new_U4706 | ~new_U2419;
  assign new_U4738 = ~new_U2487 | ~new_U2407;
  assign new_U4739 = ~new_U4705 | ~new_U2406;
  assign new_U4740 = ~new_U2394 | ~new_U4721;
  assign new_U4741 = ~INSTQUEUE_REG_12__4_ | ~new_U4716;
  assign new_U4742 = ~new_U4706 | ~new_U2418;
  assign new_U4743 = ~new_U2487 | ~new_U2405;
  assign new_U4744 = ~new_U4705 | ~new_U2404;
  assign new_U4745 = ~new_U2393 | ~new_U4721;
  assign new_U4746 = ~INSTQUEUE_REG_12__3_ | ~new_U4716;
  assign new_U4747 = ~new_U4706 | ~new_U2421;
  assign new_U4748 = ~new_U2487 | ~new_U2403;
  assign new_U4749 = ~new_U4705 | ~new_U2402;
  assign new_U4750 = ~new_U2392 | ~new_U4721;
  assign new_U4751 = ~INSTQUEUE_REG_12__2_ | ~new_U4716;
  assign new_U4752 = ~new_U4706 | ~new_U2414;
  assign new_U4753 = ~new_U2487 | ~new_U2401;
  assign new_U4754 = ~new_U4705 | ~new_U2400;
  assign new_U4755 = ~new_U2391 | ~new_U4721;
  assign new_U4756 = ~INSTQUEUE_REG_12__1_ | ~new_U4716;
  assign new_U4757 = ~new_U4706 | ~new_U2417;
  assign new_U4758 = ~new_U2487 | ~new_U2399;
  assign new_U4759 = ~new_U4705 | ~new_U2398;
  assign new_U4760 = ~new_U2390 | ~new_U4721;
  assign new_U4761 = ~INSTQUEUE_REG_12__0_ | ~new_U4716;
  assign new_U4762 = ~new_U3330;
  assign new_U4763 = ~new_U3328;
  assign new_U4764 = ~new_U2440 | ~new_U2442;
  assign new_U4765 = ~new_U3331;
  assign new_U4766 = ~new_U2434 | ~new_U2436;
  assign new_U4767 = ~new_U3332;
  assign new_U4768 = ~new_U4517 | ~new_U4516;
  assign new_U4769 = ~new_U2492 | ~new_U2358;
  assign new_U4770 = ~new_U3307 | ~new_U4769;
  assign new_U4771 = ~new_U4765 | ~new_U4770;
  assign new_U4772 = ~STATE2_REG_3_ | ~new_U3328;
  assign new_U4773 = ~new_U4767 | ~STATE2_REG_2_;
  assign new_U4774 = ~new_U4771 | ~new_U3611;
  assign new_U4775 = ~new_U2492 | ~new_U2388;
  assign new_U4776 = ~new_U3307 | ~new_U4775;
  assign new_U4777 = ~new_U4776 | ~new_U3331;
  assign new_U4778 = ~STATE2_REG_2_ | ~new_U3332;
  assign new_U4779 = ~new_U4778 | ~new_U4777;
  assign new_U4780 = ~new_U4763 | ~new_U2415;
  assign new_U4781 = ~new_U2491 | ~new_U2413;
  assign new_U4782 = ~new_U4762 | ~new_U2412;
  assign new_U4783 = ~new_U2397 | ~new_U4779;
  assign new_U4784 = ~INSTQUEUE_REG_11__7_ | ~new_U4774;
  assign new_U4785 = ~new_U4763 | ~new_U2416;
  assign new_U4786 = ~new_U2491 | ~new_U2411;
  assign new_U4787 = ~new_U4762 | ~new_U2410;
  assign new_U4788 = ~new_U2396 | ~new_U4779;
  assign new_U4789 = ~INSTQUEUE_REG_11__6_ | ~new_U4774;
  assign new_U4790 = ~new_U4763 | ~new_U2420;
  assign new_U4791 = ~new_U2491 | ~new_U2409;
  assign new_U4792 = ~new_U4762 | ~new_U2408;
  assign new_U4793 = ~new_U2395 | ~new_U4779;
  assign new_U4794 = ~INSTQUEUE_REG_11__5_ | ~new_U4774;
  assign new_U4795 = ~new_U4763 | ~new_U2419;
  assign new_U4796 = ~new_U2491 | ~new_U2407;
  assign new_U4797 = ~new_U4762 | ~new_U2406;
  assign new_U4798 = ~new_U2394 | ~new_U4779;
  assign new_U4799 = ~INSTQUEUE_REG_11__4_ | ~new_U4774;
  assign new_U4800 = ~new_U4763 | ~new_U2418;
  assign new_U4801 = ~new_U2491 | ~new_U2405;
  assign new_U4802 = ~new_U4762 | ~new_U2404;
  assign new_U4803 = ~new_U2393 | ~new_U4779;
  assign new_U4804 = ~INSTQUEUE_REG_11__3_ | ~new_U4774;
  assign new_U4805 = ~new_U4763 | ~new_U2421;
  assign new_U4806 = ~new_U2491 | ~new_U2403;
  assign new_U4807 = ~new_U4762 | ~new_U2402;
  assign new_U4808 = ~new_U2392 | ~new_U4779;
  assign new_U4809 = ~INSTQUEUE_REG_11__2_ | ~new_U4774;
  assign new_U4810 = ~new_U4763 | ~new_U2414;
  assign new_U4811 = ~new_U2491 | ~new_U2401;
  assign new_U4812 = ~new_U4762 | ~new_U2400;
  assign new_U4813 = ~new_U2391 | ~new_U4779;
  assign new_U4814 = ~INSTQUEUE_REG_11__1_ | ~new_U4774;
  assign new_U4815 = ~new_U4763 | ~new_U2417;
  assign new_U4816 = ~new_U2491 | ~new_U2399;
  assign new_U4817 = ~new_U4762 | ~new_U2398;
  assign new_U4818 = ~new_U2390 | ~new_U4779;
  assign new_U4819 = ~INSTQUEUE_REG_11__0_ | ~new_U4774;
  assign new_U4820 = ~new_U3334;
  assign new_U4821 = ~new_U3333;
  assign new_U4822 = ~new_U2440 | ~new_U2443;
  assign new_U4823 = ~new_U3335;
  assign new_U4824 = ~new_U3225;
  assign new_U4825 = ~new_U4517 | ~new_U4512;
  assign new_U4826 = ~new_U2494 | ~new_U2358;
  assign new_U4827 = ~new_U3307 | ~new_U4826;
  assign new_U4828 = ~new_U4823 | ~new_U4827;
  assign new_U4829 = ~STATE2_REG_3_ | ~new_U3333;
  assign new_U4830 = ~STATE2_REG_2_ | ~new_U3225;
  assign new_U4831 = ~new_U4828 | ~new_U3620;
  assign new_U4832 = ~new_U2494 | ~new_U2388;
  assign new_U4833 = ~new_U3307 | ~new_U4832;
  assign new_U4834 = ~new_U4833 | ~new_U3335;
  assign new_U4835 = ~STATE2_REG_2_ | ~new_U4824;
  assign new_U4836 = ~new_U4835 | ~new_U4834;
  assign new_U4837 = ~new_U4821 | ~new_U2415;
  assign new_U4838 = ~new_U2493 | ~new_U2413;
  assign new_U4839 = ~new_U4820 | ~new_U2412;
  assign new_U4840 = ~new_U2397 | ~new_U4836;
  assign new_U4841 = ~INSTQUEUE_REG_10__7_ | ~new_U4831;
  assign new_U4842 = ~new_U4821 | ~new_U2416;
  assign new_U4843 = ~new_U2493 | ~new_U2411;
  assign new_U4844 = ~new_U4820 | ~new_U2410;
  assign new_U4845 = ~new_U2396 | ~new_U4836;
  assign new_U4846 = ~INSTQUEUE_REG_10__6_ | ~new_U4831;
  assign new_U4847 = ~new_U4821 | ~new_U2420;
  assign new_U4848 = ~new_U2493 | ~new_U2409;
  assign new_U4849 = ~new_U4820 | ~new_U2408;
  assign new_U4850 = ~new_U2395 | ~new_U4836;
  assign new_U4851 = ~INSTQUEUE_REG_10__5_ | ~new_U4831;
  assign new_U4852 = ~new_U4821 | ~new_U2419;
  assign new_U4853 = ~new_U2493 | ~new_U2407;
  assign new_U4854 = ~new_U4820 | ~new_U2406;
  assign new_U4855 = ~new_U2394 | ~new_U4836;
  assign new_U4856 = ~INSTQUEUE_REG_10__4_ | ~new_U4831;
  assign new_U4857 = ~new_U4821 | ~new_U2418;
  assign new_U4858 = ~new_U2493 | ~new_U2405;
  assign new_U4859 = ~new_U4820 | ~new_U2404;
  assign new_U4860 = ~new_U2393 | ~new_U4836;
  assign new_U4861 = ~INSTQUEUE_REG_10__3_ | ~new_U4831;
  assign new_U4862 = ~new_U4821 | ~new_U2421;
  assign new_U4863 = ~new_U2493 | ~new_U2403;
  assign new_U4864 = ~new_U4820 | ~new_U2402;
  assign new_U4865 = ~new_U2392 | ~new_U4836;
  assign new_U4866 = ~INSTQUEUE_REG_10__2_ | ~new_U4831;
  assign new_U4867 = ~new_U4821 | ~new_U2414;
  assign new_U4868 = ~new_U2493 | ~new_U2401;
  assign new_U4869 = ~new_U4820 | ~new_U2400;
  assign new_U4870 = ~new_U2391 | ~new_U4836;
  assign new_U4871 = ~INSTQUEUE_REG_10__1_ | ~new_U4831;
  assign new_U4872 = ~new_U4821 | ~new_U2417;
  assign new_U4873 = ~new_U2493 | ~new_U2399;
  assign new_U4874 = ~new_U4820 | ~new_U2398;
  assign new_U4875 = ~new_U2390 | ~new_U4836;
  assign new_U4876 = ~INSTQUEUE_REG_10__0_ | ~new_U4831;
  assign new_U4877 = ~new_U3337;
  assign new_U4878 = ~new_U3336;
  assign new_U4879 = ~new_U2440 | ~new_U2444;
  assign new_U4880 = ~new_U3338;
  assign new_U4881 = ~new_U2434 | ~new_U2437;
  assign new_U4882 = ~new_U3339;
  assign new_U4883 = ~new_U4517 | ~new_U4513;
  assign new_U4884 = ~new_U2496 | ~new_U2358;
  assign new_U4885 = ~new_U3307 | ~new_U4884;
  assign new_U4886 = ~new_U4880 | ~new_U4885;
  assign new_U4887 = ~STATE2_REG_3_ | ~new_U3336;
  assign new_U4888 = ~new_U4882 | ~STATE2_REG_2_;
  assign new_U4889 = ~new_U4886 | ~new_U3629;
  assign new_U4890 = ~new_U2496 | ~new_U2388;
  assign new_U4891 = ~new_U3307 | ~new_U4890;
  assign new_U4892 = ~new_U4891 | ~new_U3338;
  assign new_U4893 = ~STATE2_REG_2_ | ~new_U3339;
  assign new_U4894 = ~new_U4893 | ~new_U4892;
  assign new_U4895 = ~new_U4878 | ~new_U2415;
  assign new_U4896 = ~new_U2495 | ~new_U2413;
  assign new_U4897 = ~new_U4877 | ~new_U2412;
  assign new_U4898 = ~new_U2397 | ~new_U4894;
  assign new_U4899 = ~INSTQUEUE_REG_9__7_ | ~new_U4889;
  assign new_U4900 = ~new_U4878 | ~new_U2416;
  assign new_U4901 = ~new_U2495 | ~new_U2411;
  assign new_U4902 = ~new_U4877 | ~new_U2410;
  assign new_U4903 = ~new_U2396 | ~new_U4894;
  assign new_U4904 = ~INSTQUEUE_REG_9__6_ | ~new_U4889;
  assign new_U4905 = ~new_U4878 | ~new_U2420;
  assign new_U4906 = ~new_U2495 | ~new_U2409;
  assign new_U4907 = ~new_U4877 | ~new_U2408;
  assign new_U4908 = ~new_U2395 | ~new_U4894;
  assign new_U4909 = ~INSTQUEUE_REG_9__5_ | ~new_U4889;
  assign new_U4910 = ~new_U4878 | ~new_U2419;
  assign new_U4911 = ~new_U2495 | ~new_U2407;
  assign new_U4912 = ~new_U4877 | ~new_U2406;
  assign new_U4913 = ~new_U2394 | ~new_U4894;
  assign new_U4914 = ~INSTQUEUE_REG_9__4_ | ~new_U4889;
  assign new_U4915 = ~new_U4878 | ~new_U2418;
  assign new_U4916 = ~new_U2495 | ~new_U2405;
  assign new_U4917 = ~new_U4877 | ~new_U2404;
  assign new_U4918 = ~new_U2393 | ~new_U4894;
  assign new_U4919 = ~INSTQUEUE_REG_9__3_ | ~new_U4889;
  assign new_U4920 = ~new_U4878 | ~new_U2421;
  assign new_U4921 = ~new_U2495 | ~new_U2403;
  assign new_U4922 = ~new_U4877 | ~new_U2402;
  assign new_U4923 = ~new_U2392 | ~new_U4894;
  assign new_U4924 = ~INSTQUEUE_REG_9__2_ | ~new_U4889;
  assign new_U4925 = ~new_U4878 | ~new_U2414;
  assign new_U4926 = ~new_U2495 | ~new_U2401;
  assign new_U4927 = ~new_U4877 | ~new_U2400;
  assign new_U4928 = ~new_U2391 | ~new_U4894;
  assign new_U4929 = ~INSTQUEUE_REG_9__1_ | ~new_U4889;
  assign new_U4930 = ~new_U4878 | ~new_U2417;
  assign new_U4931 = ~new_U2495 | ~new_U2399;
  assign new_U4932 = ~new_U4877 | ~new_U2398;
  assign new_U4933 = ~new_U2390 | ~new_U4894;
  assign new_U4934 = ~INSTQUEUE_REG_9__0_ | ~new_U4889;
  assign new_U4935 = ~new_U3341;
  assign new_U4936 = ~new_U3340;
  assign new_U4937 = ~new_U2440 | ~new_U2445;
  assign new_U4938 = ~new_U3342;
  assign new_U4939 = ~new_U3226;
  assign new_U4940 = ~new_U4517 | ~new_U2486;
  assign new_U4941 = ~new_U2498 | ~new_U2358;
  assign new_U4942 = ~new_U3307 | ~new_U4941;
  assign new_U4943 = ~new_U4938 | ~new_U4942;
  assign new_U4944 = ~STATE2_REG_3_ | ~new_U3340;
  assign new_U4945 = ~STATE2_REG_2_ | ~new_U3226;
  assign new_U4946 = ~new_U4943 | ~new_U3638;
  assign new_U4947 = ~new_U2498 | ~new_U2388;
  assign new_U4948 = ~new_U3307 | ~new_U4947;
  assign new_U4949 = ~new_U4948 | ~new_U3342;
  assign new_U4950 = ~STATE2_REG_2_ | ~new_U4939;
  assign new_U4951 = ~new_U4950 | ~new_U4949;
  assign new_U4952 = ~new_U4936 | ~new_U2415;
  assign new_U4953 = ~new_U2497 | ~new_U2413;
  assign new_U4954 = ~new_U4935 | ~new_U2412;
  assign new_U4955 = ~new_U2397 | ~new_U4951;
  assign new_U4956 = ~INSTQUEUE_REG_8__7_ | ~new_U4946;
  assign new_U4957 = ~new_U4936 | ~new_U2416;
  assign new_U4958 = ~new_U2497 | ~new_U2411;
  assign new_U4959 = ~new_U4935 | ~new_U2410;
  assign new_U4960 = ~new_U2396 | ~new_U4951;
  assign new_U4961 = ~INSTQUEUE_REG_8__6_ | ~new_U4946;
  assign new_U4962 = ~new_U4936 | ~new_U2420;
  assign new_U4963 = ~new_U2497 | ~new_U2409;
  assign new_U4964 = ~new_U4935 | ~new_U2408;
  assign new_U4965 = ~new_U2395 | ~new_U4951;
  assign new_U4966 = ~INSTQUEUE_REG_8__5_ | ~new_U4946;
  assign new_U4967 = ~new_U4936 | ~new_U2419;
  assign new_U4968 = ~new_U2497 | ~new_U2407;
  assign new_U4969 = ~new_U4935 | ~new_U2406;
  assign new_U4970 = ~new_U2394 | ~new_U4951;
  assign new_U4971 = ~INSTQUEUE_REG_8__4_ | ~new_U4946;
  assign new_U4972 = ~new_U4936 | ~new_U2418;
  assign new_U4973 = ~new_U2497 | ~new_U2405;
  assign new_U4974 = ~new_U4935 | ~new_U2404;
  assign new_U4975 = ~new_U2393 | ~new_U4951;
  assign new_U4976 = ~INSTQUEUE_REG_8__3_ | ~new_U4946;
  assign new_U4977 = ~new_U4936 | ~new_U2421;
  assign new_U4978 = ~new_U2497 | ~new_U2403;
  assign new_U4979 = ~new_U4935 | ~new_U2402;
  assign new_U4980 = ~new_U2392 | ~new_U4951;
  assign new_U4981 = ~INSTQUEUE_REG_8__2_ | ~new_U4946;
  assign new_U4982 = ~new_U4936 | ~new_U2414;
  assign new_U4983 = ~new_U2497 | ~new_U2401;
  assign new_U4984 = ~new_U4935 | ~new_U2400;
  assign new_U4985 = ~new_U2391 | ~new_U4951;
  assign new_U4986 = ~INSTQUEUE_REG_8__1_ | ~new_U4946;
  assign new_U4987 = ~new_U4936 | ~new_U2417;
  assign new_U4988 = ~new_U2497 | ~new_U2399;
  assign new_U4989 = ~new_U4935 | ~new_U2398;
  assign new_U4990 = ~new_U2390 | ~new_U4951;
  assign new_U4991 = ~INSTQUEUE_REG_8__0_ | ~new_U4946;
  assign new_U4992 = ~new_U3346;
  assign new_U4993 = ~new_U2439 | ~new_U2442;
  assign new_U4994 = ~new_U3348;
  assign new_U4995 = ~new_U2433 | ~new_U2436;
  assign new_U4996 = ~new_U3349;
  assign new_U4997 = ~new_U2500 | ~new_U2358;
  assign new_U4998 = ~new_U3307 | ~new_U4997;
  assign new_U4999 = ~new_U4994 | ~new_U4998;
  assign new_U5000 = ~STATE2_REG_3_ | ~new_U3343;
  assign new_U5001 = ~new_U4996 | ~STATE2_REG_2_;
  assign new_U5002 = ~new_U4999 | ~new_U3647;
  assign new_U5003 = ~new_U2500 | ~new_U2388;
  assign new_U5004 = ~new_U3307 | ~new_U5003;
  assign new_U5005 = ~new_U5004 | ~new_U3348;
  assign new_U5006 = ~STATE2_REG_2_ | ~new_U3349;
  assign new_U5007 = ~new_U5006 | ~new_U5005;
  assign new_U5008 = ~new_U4525 | ~new_U2415;
  assign new_U5009 = ~new_U4226 | ~new_U2413;
  assign new_U5010 = ~new_U4992 | ~new_U2412;
  assign new_U5011 = ~new_U2397 | ~new_U5007;
  assign new_U5012 = ~INSTQUEUE_REG_7__7_ | ~new_U5002;
  assign new_U5013 = ~new_U4525 | ~new_U2416;
  assign new_U5014 = ~new_U4226 | ~new_U2411;
  assign new_U5015 = ~new_U4992 | ~new_U2410;
  assign new_U5016 = ~new_U2396 | ~new_U5007;
  assign new_U5017 = ~INSTQUEUE_REG_7__6_ | ~new_U5002;
  assign new_U5018 = ~new_U4525 | ~new_U2420;
  assign new_U5019 = ~new_U4226 | ~new_U2409;
  assign new_U5020 = ~new_U4992 | ~new_U2408;
  assign new_U5021 = ~new_U2395 | ~new_U5007;
  assign new_U5022 = ~INSTQUEUE_REG_7__5_ | ~new_U5002;
  assign new_U5023 = ~new_U4525 | ~new_U2419;
  assign new_U5024 = ~new_U4226 | ~new_U2407;
  assign new_U5025 = ~new_U4992 | ~new_U2406;
  assign new_U5026 = ~new_U2394 | ~new_U5007;
  assign new_U5027 = ~INSTQUEUE_REG_7__4_ | ~new_U5002;
  assign new_U5028 = ~new_U4525 | ~new_U2418;
  assign new_U5029 = ~new_U4226 | ~new_U2405;
  assign new_U5030 = ~new_U4992 | ~new_U2404;
  assign new_U5031 = ~new_U2393 | ~new_U5007;
  assign new_U5032 = ~INSTQUEUE_REG_7__3_ | ~new_U5002;
  assign new_U5033 = ~new_U4525 | ~new_U2421;
  assign new_U5034 = ~new_U4226 | ~new_U2403;
  assign new_U5035 = ~new_U4992 | ~new_U2402;
  assign new_U5036 = ~new_U2392 | ~new_U5007;
  assign new_U5037 = ~INSTQUEUE_REG_7__2_ | ~new_U5002;
  assign new_U5038 = ~new_U4525 | ~new_U2414;
  assign new_U5039 = ~new_U4226 | ~new_U2401;
  assign new_U5040 = ~new_U4992 | ~new_U2400;
  assign new_U5041 = ~new_U2391 | ~new_U5007;
  assign new_U5042 = ~INSTQUEUE_REG_7__1_ | ~new_U5002;
  assign new_U5043 = ~new_U4525 | ~new_U2417;
  assign new_U5044 = ~new_U4226 | ~new_U2399;
  assign new_U5045 = ~new_U4992 | ~new_U2398;
  assign new_U5046 = ~new_U2390 | ~new_U5007;
  assign new_U5047 = ~INSTQUEUE_REG_7__0_ | ~new_U5002;
  assign new_U5048 = ~new_U3351;
  assign new_U5049 = ~new_U3350;
  assign new_U5050 = ~new_U2439 | ~new_U2443;
  assign new_U5051 = ~new_U3352;
  assign new_U5052 = ~new_U3227;
  assign new_U5053 = ~new_U4512 | ~new_U2474;
  assign new_U5054 = ~new_U2502 | ~new_U2358;
  assign new_U5055 = ~new_U3307 | ~new_U5054;
  assign new_U5056 = ~new_U5051 | ~new_U5055;
  assign new_U5057 = ~STATE2_REG_3_ | ~new_U3350;
  assign new_U5058 = ~STATE2_REG_2_ | ~new_U3227;
  assign new_U5059 = ~new_U5056 | ~new_U3656;
  assign new_U5060 = ~new_U2502 | ~new_U2388;
  assign new_U5061 = ~new_U3307 | ~new_U5060;
  assign new_U5062 = ~new_U5061 | ~new_U3352;
  assign new_U5063 = ~STATE2_REG_2_ | ~new_U5052;
  assign new_U5064 = ~new_U5063 | ~new_U5062;
  assign new_U5065 = ~new_U5049 | ~new_U2415;
  assign new_U5066 = ~new_U2501 | ~new_U2413;
  assign new_U5067 = ~new_U5048 | ~new_U2412;
  assign new_U5068 = ~new_U2397 | ~new_U5064;
  assign new_U5069 = ~INSTQUEUE_REG_6__7_ | ~new_U5059;
  assign new_U5070 = ~new_U5049 | ~new_U2416;
  assign new_U5071 = ~new_U2501 | ~new_U2411;
  assign new_U5072 = ~new_U5048 | ~new_U2410;
  assign new_U5073 = ~new_U2396 | ~new_U5064;
  assign new_U5074 = ~INSTQUEUE_REG_6__6_ | ~new_U5059;
  assign new_U5075 = ~new_U5049 | ~new_U2420;
  assign new_U5076 = ~new_U2501 | ~new_U2409;
  assign new_U5077 = ~new_U5048 | ~new_U2408;
  assign new_U5078 = ~new_U2395 | ~new_U5064;
  assign new_U5079 = ~INSTQUEUE_REG_6__5_ | ~new_U5059;
  assign new_U5080 = ~new_U5049 | ~new_U2419;
  assign new_U5081 = ~new_U2501 | ~new_U2407;
  assign new_U5082 = ~new_U5048 | ~new_U2406;
  assign new_U5083 = ~new_U2394 | ~new_U5064;
  assign new_U5084 = ~INSTQUEUE_REG_6__4_ | ~new_U5059;
  assign new_U5085 = ~new_U5049 | ~new_U2418;
  assign new_U5086 = ~new_U2501 | ~new_U2405;
  assign new_U5087 = ~new_U5048 | ~new_U2404;
  assign new_U5088 = ~new_U2393 | ~new_U5064;
  assign new_U5089 = ~INSTQUEUE_REG_6__3_ | ~new_U5059;
  assign new_U5090 = ~new_U5049 | ~new_U2421;
  assign new_U5091 = ~new_U2501 | ~new_U2403;
  assign new_U5092 = ~new_U5048 | ~new_U2402;
  assign new_U5093 = ~new_U2392 | ~new_U5064;
  assign new_U5094 = ~INSTQUEUE_REG_6__2_ | ~new_U5059;
  assign new_U5095 = ~new_U5049 | ~new_U2414;
  assign new_U5096 = ~new_U2501 | ~new_U2401;
  assign new_U5097 = ~new_U5048 | ~new_U2400;
  assign new_U5098 = ~new_U2391 | ~new_U5064;
  assign new_U5099 = ~INSTQUEUE_REG_6__1_ | ~new_U5059;
  assign new_U5100 = ~new_U5049 | ~new_U2417;
  assign new_U5101 = ~new_U2501 | ~new_U2399;
  assign new_U5102 = ~new_U5048 | ~new_U2398;
  assign new_U5103 = ~new_U2390 | ~new_U5064;
  assign new_U5104 = ~INSTQUEUE_REG_6__0_ | ~new_U5059;
  assign new_U5105 = ~new_U3354;
  assign new_U5106 = ~new_U3353;
  assign new_U5107 = ~new_U2439 | ~new_U2444;
  assign new_U5108 = ~new_U3355;
  assign new_U5109 = ~new_U2433 | ~new_U2437;
  assign new_U5110 = ~new_U3356;
  assign new_U5111 = ~new_U4513 | ~new_U2474;
  assign new_U5112 = ~new_U2504 | ~new_U2358;
  assign new_U5113 = ~new_U3307 | ~new_U5112;
  assign new_U5114 = ~new_U5108 | ~new_U5113;
  assign new_U5115 = ~STATE2_REG_3_ | ~new_U3353;
  assign new_U5116 = ~new_U5110 | ~STATE2_REG_2_;
  assign new_U5117 = ~new_U5114 | ~new_U3665;
  assign new_U5118 = ~new_U2504 | ~new_U2388;
  assign new_U5119 = ~new_U3307 | ~new_U5118;
  assign new_U5120 = ~new_U5119 | ~new_U3355;
  assign new_U5121 = ~STATE2_REG_2_ | ~new_U3356;
  assign new_U5122 = ~new_U5121 | ~new_U5120;
  assign new_U5123 = ~new_U5106 | ~new_U2415;
  assign new_U5124 = ~new_U2503 | ~new_U2413;
  assign new_U5125 = ~new_U5105 | ~new_U2412;
  assign new_U5126 = ~new_U2397 | ~new_U5122;
  assign new_U5127 = ~INSTQUEUE_REG_5__7_ | ~new_U5117;
  assign new_U5128 = ~new_U5106 | ~new_U2416;
  assign new_U5129 = ~new_U2503 | ~new_U2411;
  assign new_U5130 = ~new_U5105 | ~new_U2410;
  assign new_U5131 = ~new_U2396 | ~new_U5122;
  assign new_U5132 = ~INSTQUEUE_REG_5__6_ | ~new_U5117;
  assign new_U5133 = ~new_U5106 | ~new_U2420;
  assign new_U5134 = ~new_U2503 | ~new_U2409;
  assign new_U5135 = ~new_U5105 | ~new_U2408;
  assign new_U5136 = ~new_U2395 | ~new_U5122;
  assign new_U5137 = ~INSTQUEUE_REG_5__5_ | ~new_U5117;
  assign new_U5138 = ~new_U5106 | ~new_U2419;
  assign new_U5139 = ~new_U2503 | ~new_U2407;
  assign new_U5140 = ~new_U5105 | ~new_U2406;
  assign new_U5141 = ~new_U2394 | ~new_U5122;
  assign new_U5142 = ~INSTQUEUE_REG_5__4_ | ~new_U5117;
  assign new_U5143 = ~new_U5106 | ~new_U2418;
  assign new_U5144 = ~new_U2503 | ~new_U2405;
  assign new_U5145 = ~new_U5105 | ~new_U2404;
  assign new_U5146 = ~new_U2393 | ~new_U5122;
  assign new_U5147 = ~INSTQUEUE_REG_5__3_ | ~new_U5117;
  assign new_U5148 = ~new_U5106 | ~new_U2421;
  assign new_U5149 = ~new_U2503 | ~new_U2403;
  assign new_U5150 = ~new_U5105 | ~new_U2402;
  assign new_U5151 = ~new_U2392 | ~new_U5122;
  assign new_U5152 = ~INSTQUEUE_REG_5__2_ | ~new_U5117;
  assign new_U5153 = ~new_U5106 | ~new_U2414;
  assign new_U5154 = ~new_U2503 | ~new_U2401;
  assign new_U5155 = ~new_U5105 | ~new_U2400;
  assign new_U5156 = ~new_U2391 | ~new_U5122;
  assign new_U5157 = ~INSTQUEUE_REG_5__1_ | ~new_U5117;
  assign new_U5158 = ~new_U5106 | ~new_U2417;
  assign new_U5159 = ~new_U2503 | ~new_U2399;
  assign new_U5160 = ~new_U5105 | ~new_U2398;
  assign new_U5161 = ~new_U2390 | ~new_U5122;
  assign new_U5162 = ~INSTQUEUE_REG_5__0_ | ~new_U5117;
  assign new_U5163 = ~new_U3358;
  assign new_U5164 = ~new_U3357;
  assign new_U5165 = ~new_U2439 | ~new_U2445;
  assign new_U5166 = ~new_U3359;
  assign new_U5167 = ~new_U3228;
  assign new_U5168 = ~new_U2486 | ~new_U2474;
  assign new_U5169 = ~new_U2506 | ~new_U2358;
  assign new_U5170 = ~new_U3307 | ~new_U5169;
  assign new_U5171 = ~new_U5166 | ~new_U5170;
  assign new_U5172 = ~STATE2_REG_3_ | ~new_U3357;
  assign new_U5173 = ~STATE2_REG_2_ | ~new_U3228;
  assign new_U5174 = ~new_U5171 | ~new_U3674;
  assign new_U5175 = ~new_U2506 | ~new_U2388;
  assign new_U5176 = ~new_U3307 | ~new_U5175;
  assign new_U5177 = ~new_U5176 | ~new_U3359;
  assign new_U5178 = ~STATE2_REG_2_ | ~new_U5167;
  assign new_U5179 = ~new_U5178 | ~new_U5177;
  assign new_U5180 = ~new_U5164 | ~new_U2415;
  assign new_U5181 = ~new_U2505 | ~new_U2413;
  assign new_U5182 = ~new_U5163 | ~new_U2412;
  assign new_U5183 = ~new_U2397 | ~new_U5179;
  assign new_U5184 = ~INSTQUEUE_REG_4__7_ | ~new_U5174;
  assign new_U5185 = ~new_U5164 | ~new_U2416;
  assign new_U5186 = ~new_U2505 | ~new_U2411;
  assign new_U5187 = ~new_U5163 | ~new_U2410;
  assign new_U5188 = ~new_U2396 | ~new_U5179;
  assign new_U5189 = ~INSTQUEUE_REG_4__6_ | ~new_U5174;
  assign new_U5190 = ~new_U5164 | ~new_U2420;
  assign new_U5191 = ~new_U2505 | ~new_U2409;
  assign new_U5192 = ~new_U5163 | ~new_U2408;
  assign new_U5193 = ~new_U2395 | ~new_U5179;
  assign new_U5194 = ~INSTQUEUE_REG_4__5_ | ~new_U5174;
  assign new_U5195 = ~new_U5164 | ~new_U2419;
  assign new_U5196 = ~new_U2505 | ~new_U2407;
  assign new_U5197 = ~new_U5163 | ~new_U2406;
  assign new_U5198 = ~new_U2394 | ~new_U5179;
  assign new_U5199 = ~INSTQUEUE_REG_4__4_ | ~new_U5174;
  assign new_U5200 = ~new_U5164 | ~new_U2418;
  assign new_U5201 = ~new_U2505 | ~new_U2405;
  assign new_U5202 = ~new_U5163 | ~new_U2404;
  assign new_U5203 = ~new_U2393 | ~new_U5179;
  assign new_U5204 = ~INSTQUEUE_REG_4__3_ | ~new_U5174;
  assign new_U5205 = ~new_U5164 | ~new_U2421;
  assign new_U5206 = ~new_U2505 | ~new_U2403;
  assign new_U5207 = ~new_U5163 | ~new_U2402;
  assign new_U5208 = ~new_U2392 | ~new_U5179;
  assign new_U5209 = ~INSTQUEUE_REG_4__2_ | ~new_U5174;
  assign new_U5210 = ~new_U5164 | ~new_U2414;
  assign new_U5211 = ~new_U2505 | ~new_U2401;
  assign new_U5212 = ~new_U5163 | ~new_U2400;
  assign new_U5213 = ~new_U2391 | ~new_U5179;
  assign new_U5214 = ~INSTQUEUE_REG_4__1_ | ~new_U5174;
  assign new_U5215 = ~new_U5164 | ~new_U2417;
  assign new_U5216 = ~new_U2505 | ~new_U2399;
  assign new_U5217 = ~new_U5163 | ~new_U2398;
  assign new_U5218 = ~new_U2390 | ~new_U5179;
  assign new_U5219 = ~INSTQUEUE_REG_4__0_ | ~new_U5174;
  assign new_U5220 = ~new_U3361;
  assign new_U5221 = ~new_U3360;
  assign new_U5222 = ~new_U2441 | ~new_U2442;
  assign new_U5223 = ~new_U3362;
  assign new_U5224 = ~new_U2435 | ~new_U2436;
  assign new_U5225 = ~new_U3363;
  assign new_U5226 = ~new_U2508 | ~new_U4516;
  assign new_U5227 = ~new_U2511 | ~new_U2358;
  assign new_U5228 = ~new_U3307 | ~new_U5227;
  assign new_U5229 = ~new_U5223 | ~new_U5228;
  assign new_U5230 = ~STATE2_REG_3_ | ~new_U3360;
  assign new_U5231 = ~new_U5225 | ~STATE2_REG_2_;
  assign new_U5232 = ~new_U5229 | ~new_U3683;
  assign new_U5233 = ~new_U2511 | ~new_U2388;
  assign new_U5234 = ~new_U3307 | ~new_U5233;
  assign new_U5235 = ~new_U5234 | ~new_U3362;
  assign new_U5236 = ~STATE2_REG_2_ | ~new_U3363;
  assign new_U5237 = ~new_U5236 | ~new_U5235;
  assign new_U5238 = ~new_U5221 | ~new_U2415;
  assign new_U5239 = ~new_U2509 | ~new_U2413;
  assign new_U5240 = ~new_U5220 | ~new_U2412;
  assign new_U5241 = ~new_U2397 | ~new_U5237;
  assign new_U5242 = ~INSTQUEUE_REG_3__7_ | ~new_U5232;
  assign new_U5243 = ~new_U5221 | ~new_U2416;
  assign new_U5244 = ~new_U2509 | ~new_U2411;
  assign new_U5245 = ~new_U5220 | ~new_U2410;
  assign new_U5246 = ~new_U2396 | ~new_U5237;
  assign new_U5247 = ~INSTQUEUE_REG_3__6_ | ~new_U5232;
  assign new_U5248 = ~new_U5221 | ~new_U2420;
  assign new_U5249 = ~new_U2509 | ~new_U2409;
  assign new_U5250 = ~new_U5220 | ~new_U2408;
  assign new_U5251 = ~new_U2395 | ~new_U5237;
  assign new_U5252 = ~INSTQUEUE_REG_3__5_ | ~new_U5232;
  assign new_U5253 = ~new_U5221 | ~new_U2419;
  assign new_U5254 = ~new_U2509 | ~new_U2407;
  assign new_U5255 = ~new_U5220 | ~new_U2406;
  assign new_U5256 = ~new_U2394 | ~new_U5237;
  assign new_U5257 = ~INSTQUEUE_REG_3__4_ | ~new_U5232;
  assign new_U5258 = ~new_U5221 | ~new_U2418;
  assign new_U5259 = ~new_U2509 | ~new_U2405;
  assign new_U5260 = ~new_U5220 | ~new_U2404;
  assign new_U5261 = ~new_U2393 | ~new_U5237;
  assign new_U5262 = ~INSTQUEUE_REG_3__3_ | ~new_U5232;
  assign new_U5263 = ~new_U5221 | ~new_U2421;
  assign new_U5264 = ~new_U2509 | ~new_U2403;
  assign new_U5265 = ~new_U5220 | ~new_U2402;
  assign new_U5266 = ~new_U2392 | ~new_U5237;
  assign new_U5267 = ~INSTQUEUE_REG_3__2_ | ~new_U5232;
  assign new_U5268 = ~new_U5221 | ~new_U2414;
  assign new_U5269 = ~new_U2509 | ~new_U2401;
  assign new_U5270 = ~new_U5220 | ~new_U2400;
  assign new_U5271 = ~new_U2391 | ~new_U5237;
  assign new_U5272 = ~INSTQUEUE_REG_3__1_ | ~new_U5232;
  assign new_U5273 = ~new_U5221 | ~new_U2417;
  assign new_U5274 = ~new_U2509 | ~new_U2399;
  assign new_U5275 = ~new_U5220 | ~new_U2398;
  assign new_U5276 = ~new_U2390 | ~new_U5237;
  assign new_U5277 = ~INSTQUEUE_REG_3__0_ | ~new_U5232;
  assign new_U5278 = ~new_U3365;
  assign new_U5279 = ~new_U3364;
  assign new_U5280 = ~new_U2441 | ~new_U2443;
  assign new_U5281 = ~new_U3366;
  assign new_U5282 = ~new_U3229;
  assign new_U5283 = ~new_U2508 | ~new_U4512;
  assign new_U5284 = ~new_U2513 | ~new_U2358;
  assign new_U5285 = ~new_U3307 | ~new_U5284;
  assign new_U5286 = ~new_U5281 | ~new_U5285;
  assign new_U5287 = ~STATE2_REG_3_ | ~new_U3364;
  assign new_U5288 = ~STATE2_REG_2_ | ~new_U3229;
  assign new_U5289 = ~new_U5286 | ~new_U3692;
  assign new_U5290 = ~new_U2513 | ~new_U2388;
  assign new_U5291 = ~new_U3307 | ~new_U5290;
  assign new_U5292 = ~new_U5291 | ~new_U3366;
  assign new_U5293 = ~STATE2_REG_2_ | ~new_U5282;
  assign new_U5294 = ~new_U5293 | ~new_U5292;
  assign new_U5295 = ~new_U5279 | ~new_U2415;
  assign new_U5296 = ~new_U2512 | ~new_U2413;
  assign new_U5297 = ~new_U5278 | ~new_U2412;
  assign new_U5298 = ~new_U2397 | ~new_U5294;
  assign new_U5299 = ~INSTQUEUE_REG_2__7_ | ~new_U5289;
  assign new_U5300 = ~new_U5279 | ~new_U2416;
  assign new_U5301 = ~new_U2512 | ~new_U2411;
  assign new_U5302 = ~new_U5278 | ~new_U2410;
  assign new_U5303 = ~new_U2396 | ~new_U5294;
  assign new_U5304 = ~INSTQUEUE_REG_2__6_ | ~new_U5289;
  assign new_U5305 = ~new_U5279 | ~new_U2420;
  assign new_U5306 = ~new_U2512 | ~new_U2409;
  assign new_U5307 = ~new_U5278 | ~new_U2408;
  assign new_U5308 = ~new_U2395 | ~new_U5294;
  assign new_U5309 = ~INSTQUEUE_REG_2__5_ | ~new_U5289;
  assign new_U5310 = ~new_U5279 | ~new_U2419;
  assign new_U5311 = ~new_U2512 | ~new_U2407;
  assign new_U5312 = ~new_U5278 | ~new_U2406;
  assign new_U5313 = ~new_U2394 | ~new_U5294;
  assign new_U5314 = ~INSTQUEUE_REG_2__4_ | ~new_U5289;
  assign new_U5315 = ~new_U5279 | ~new_U2418;
  assign new_U5316 = ~new_U2512 | ~new_U2405;
  assign new_U5317 = ~new_U5278 | ~new_U2404;
  assign new_U5318 = ~new_U2393 | ~new_U5294;
  assign new_U5319 = ~INSTQUEUE_REG_2__3_ | ~new_U5289;
  assign new_U5320 = ~new_U5279 | ~new_U2421;
  assign new_U5321 = ~new_U2512 | ~new_U2403;
  assign new_U5322 = ~new_U5278 | ~new_U2402;
  assign new_U5323 = ~new_U2392 | ~new_U5294;
  assign new_U5324 = ~INSTQUEUE_REG_2__2_ | ~new_U5289;
  assign new_U5325 = ~new_U5279 | ~new_U2414;
  assign new_U5326 = ~new_U2512 | ~new_U2401;
  assign new_U5327 = ~new_U5278 | ~new_U2400;
  assign new_U5328 = ~new_U2391 | ~new_U5294;
  assign new_U5329 = ~INSTQUEUE_REG_2__1_ | ~new_U5289;
  assign new_U5330 = ~new_U5279 | ~new_U2417;
  assign new_U5331 = ~new_U2512 | ~new_U2399;
  assign new_U5332 = ~new_U5278 | ~new_U2398;
  assign new_U5333 = ~new_U2390 | ~new_U5294;
  assign new_U5334 = ~INSTQUEUE_REG_2__0_ | ~new_U5289;
  assign new_U5335 = ~new_U3368;
  assign new_U5336 = ~new_U3367;
  assign new_U5337 = ~new_U2441 | ~new_U2444;
  assign new_U5338 = ~new_U3369;
  assign new_U5339 = ~new_U2435 | ~new_U2437;
  assign new_U5340 = ~new_U3370;
  assign new_U5341 = ~new_U2508 | ~new_U4513;
  assign new_U5342 = ~new_U2515 | ~new_U2358;
  assign new_U5343 = ~new_U3307 | ~new_U5342;
  assign new_U5344 = ~new_U5338 | ~new_U5343;
  assign new_U5345 = ~STATE2_REG_3_ | ~new_U3367;
  assign new_U5346 = ~new_U5340 | ~STATE2_REG_2_;
  assign new_U5347 = ~new_U5344 | ~new_U3701;
  assign new_U5348 = ~new_U2515 | ~new_U2388;
  assign new_U5349 = ~new_U3307 | ~new_U5348;
  assign new_U5350 = ~new_U5349 | ~new_U3369;
  assign new_U5351 = ~STATE2_REG_2_ | ~new_U3370;
  assign new_U5352 = ~new_U5351 | ~new_U5350;
  assign new_U5353 = ~new_U5336 | ~new_U2415;
  assign new_U5354 = ~new_U2514 | ~new_U2413;
  assign new_U5355 = ~new_U5335 | ~new_U2412;
  assign new_U5356 = ~new_U2397 | ~new_U5352;
  assign new_U5357 = ~INSTQUEUE_REG_1__7_ | ~new_U5347;
  assign new_U5358 = ~new_U5336 | ~new_U2416;
  assign new_U5359 = ~new_U2514 | ~new_U2411;
  assign new_U5360 = ~new_U5335 | ~new_U2410;
  assign new_U5361 = ~new_U2396 | ~new_U5352;
  assign new_U5362 = ~INSTQUEUE_REG_1__6_ | ~new_U5347;
  assign new_U5363 = ~new_U5336 | ~new_U2420;
  assign new_U5364 = ~new_U2514 | ~new_U2409;
  assign new_U5365 = ~new_U5335 | ~new_U2408;
  assign new_U5366 = ~new_U2395 | ~new_U5352;
  assign new_U5367 = ~INSTQUEUE_REG_1__5_ | ~new_U5347;
  assign new_U5368 = ~new_U5336 | ~new_U2419;
  assign new_U5369 = ~new_U2514 | ~new_U2407;
  assign new_U5370 = ~new_U5335 | ~new_U2406;
  assign new_U5371 = ~new_U2394 | ~new_U5352;
  assign new_U5372 = ~INSTQUEUE_REG_1__4_ | ~new_U5347;
  assign new_U5373 = ~new_U5336 | ~new_U2418;
  assign new_U5374 = ~new_U2514 | ~new_U2405;
  assign new_U5375 = ~new_U5335 | ~new_U2404;
  assign new_U5376 = ~new_U2393 | ~new_U5352;
  assign new_U5377 = ~INSTQUEUE_REG_1__3_ | ~new_U5347;
  assign new_U5378 = ~new_U5336 | ~new_U2421;
  assign new_U5379 = ~new_U2514 | ~new_U2403;
  assign new_U5380 = ~new_U5335 | ~new_U2402;
  assign new_U5381 = ~new_U2392 | ~new_U5352;
  assign new_U5382 = ~INSTQUEUE_REG_1__2_ | ~new_U5347;
  assign new_U5383 = ~new_U5336 | ~new_U2414;
  assign new_U5384 = ~new_U2514 | ~new_U2401;
  assign new_U5385 = ~new_U5335 | ~new_U2400;
  assign new_U5386 = ~new_U2391 | ~new_U5352;
  assign new_U5387 = ~INSTQUEUE_REG_1__1_ | ~new_U5347;
  assign new_U5388 = ~new_U5336 | ~new_U2417;
  assign new_U5389 = ~new_U2514 | ~new_U2399;
  assign new_U5390 = ~new_U5335 | ~new_U2398;
  assign new_U5391 = ~new_U2390 | ~new_U5352;
  assign new_U5392 = ~INSTQUEUE_REG_1__0_ | ~new_U5347;
  assign new_U5393 = ~new_U3372;
  assign new_U5394 = ~new_U3371;
  assign new_U5395 = ~new_U2441 | ~new_U2445;
  assign new_U5396 = ~new_U3373;
  assign new_U5397 = ~new_U3230;
  assign new_U5398 = ~new_U2508 | ~new_U2486;
  assign new_U5399 = ~new_U2517 | ~new_U2358;
  assign new_U5400 = ~new_U3307 | ~new_U5399;
  assign new_U5401 = ~new_U5396 | ~new_U5400;
  assign new_U5402 = ~STATE2_REG_3_ | ~new_U3371;
  assign new_U5403 = ~STATE2_REG_2_ | ~new_U3230;
  assign new_U5404 = ~new_U5401 | ~new_U3710;
  assign new_U5405 = ~new_U2517 | ~new_U2388;
  assign new_U5406 = ~new_U3307 | ~new_U5405;
  assign new_U5407 = ~new_U5406 | ~new_U3373;
  assign new_U5408 = ~STATE2_REG_2_ | ~new_U5397;
  assign new_U5409 = ~new_U5408 | ~new_U5407;
  assign new_U5410 = ~new_U5394 | ~new_U2415;
  assign new_U5411 = ~new_U2516 | ~new_U2413;
  assign new_U5412 = ~new_U5393 | ~new_U2412;
  assign new_U5413 = ~new_U2397 | ~new_U5409;
  assign new_U5414 = ~INSTQUEUE_REG_0__7_ | ~new_U5404;
  assign new_U5415 = ~new_U5394 | ~new_U2416;
  assign new_U5416 = ~new_U2516 | ~new_U2411;
  assign new_U5417 = ~new_U5393 | ~new_U2410;
  assign new_U5418 = ~new_U2396 | ~new_U5409;
  assign new_U5419 = ~INSTQUEUE_REG_0__6_ | ~new_U5404;
  assign new_U5420 = ~new_U5394 | ~new_U2420;
  assign new_U5421 = ~new_U2516 | ~new_U2409;
  assign new_U5422 = ~new_U5393 | ~new_U2408;
  assign new_U5423 = ~new_U2395 | ~new_U5409;
  assign new_U5424 = ~INSTQUEUE_REG_0__5_ | ~new_U5404;
  assign new_U5425 = ~new_U5394 | ~new_U2419;
  assign new_U5426 = ~new_U2516 | ~new_U2407;
  assign new_U5427 = ~new_U5393 | ~new_U2406;
  assign new_U5428 = ~new_U2394 | ~new_U5409;
  assign new_U5429 = ~new_U5394 | ~new_U2418;
  assign new_U5430 = ~new_U2516 | ~new_U2405;
  assign new_U5431 = ~new_U5393 | ~new_U2404;
  assign new_U5432 = ~new_U2393 | ~new_U5409;
  assign new_U5433 = ~INSTQUEUE_REG_0__3_ | ~new_U5404;
  assign new_U5434 = ~new_U5394 | ~new_U2421;
  assign new_U5435 = ~new_U2516 | ~new_U2403;
  assign new_U5436 = ~new_U5393 | ~new_U2402;
  assign new_U5437 = ~new_U2392 | ~new_U5409;
  assign new_U5438 = ~INSTQUEUE_REG_0__2_ | ~new_U5404;
  assign new_U5439 = ~new_U5394 | ~new_U2414;
  assign new_U5440 = ~new_U2516 | ~new_U2401;
  assign new_U5441 = ~new_U5393 | ~new_U2400;
  assign new_U5442 = ~new_U2391 | ~new_U5409;
  assign new_U5443 = ~INSTQUEUE_REG_0__1_ | ~new_U5404;
  assign new_U5444 = ~new_U5394 | ~new_U2417;
  assign new_U5445 = ~new_U2516 | ~new_U2399;
  assign new_U5446 = ~new_U5393 | ~new_U2398;
  assign new_U5447 = ~new_U2390 | ~new_U5409;
  assign new_U5448 = ~INSTQUEUE_REG_0__0_ | ~new_U5404;
  assign new_U5449 = ~new_U3410;
  assign new_U5450 = ~new_U4491 | ~new_U3378 | ~new_U3381;
  assign new_U5451 = ~new_U4448 | ~new_U4388 | ~new_U4161;
  assign new_U5452 = ~new_U3231;
  assign new_U5453 = ~new_U4482 | ~new_U3276;
  assign new_U5454 = ~new_U5452 | ~new_U5453 | ~new_U3270;
  assign new_U5455 = ~new_U3720 | ~new_U2452;
  assign new_U5456 = ~new_U4196 | ~new_U5450;
  assign new_U5457 = ~new_U3721 | ~new_U7597;
  assign new_U5458 = ~new_GTE_485_U6 | ~new_U4203 | ~new_U3244;
  assign new_U5459 = ~new_U2449 | ~new_U7482;
  assign new_U5460 = ~new_U4245 | ~new_U4491;
  assign new_U5461 = ~new_U4170;
  assign new_U5462 = ~new_U2368 | ~new_U4170;
  assign new_U5463 = ~STATE2_REG_3_ | ~new_U3281;
  assign new_U5464 = ~new_U4160;
  assign new_U5465 = ~INSTQUEUERD_ADDR_REG_1_ | ~INSTQUEUERD_ADDR_REG_2_;
  assign new_U5466 = ~INSTQUEUERD_ADDR_REG_3_ | ~new_U5465;
  assign new_U5467 = ~new_U4369 | ~INSTQUEUERD_ADDR_REG_1_;
  assign new_U5468 = ~new_U3429;
  assign new_U5469 = ~new_U3486 | ~INSTQUEUERD_ADDR_REG_2_;
  assign new_U5470 = ~INSTQUEUERD_ADDR_REG_3_ | ~new_U5469;
  assign new_U5471 = ~new_U3425;
  assign new_U5472 = ~new_U3262 | ~new_U3251;
  assign new_U5473 = ~INSTQUEUERD_ADDR_REG_3_ | ~new_U5472;
  assign new_U5474 = ~new_U2469 | ~new_U3262;
  assign new_U5475 = ~new_U4482 | ~new_U3277;
  assign new_U5476 = ~new_U4388 | ~new_U2605;
  assign new_U5477 = ~new_U7482 | ~new_U7692 | ~new_U7691;
  assign new_U5478 = ~new_U4437 | ~new_U5476;
  assign new_U5479 = ~new_U3396 | ~new_U4388 | ~new_U3381;
  assign new_U5480 = ~new_U5479 | ~new_U4159;
  assign new_U5481 = ~new_U7617 | ~new_U5480;
  assign new_U5482 = ~new_U4448 | ~new_U4159;
  assign new_U5483 = ~new_U3382 | ~new_U5482;
  assign new_U5484 = ~new_U4196 | ~new_U5450;
  assign new_U5485 = ~new_U4245 | ~new_U4491;
  assign new_U5486 = ~new_U5483 | ~new_U3258;
  assign new_U5487 = ~new_U4482 | ~new_U7695;
  assign new_U5488 = ~new_U4178 | ~new_U3231;
  assign new_U5489 = ~new_U3279 | ~new_U4205;
  assign new_U5490 = ~new_U3728 | ~new_U5489;
  assign new_U5491 = ~new_R2182_U25 | ~new_U7497;
  assign new_U5492 = ~new_U4206 | ~new_U3425;
  assign new_U5493 = ~new_U4202 | ~new_U3429;
  assign new_U5494 = ~new_U5491 | ~new_U3735;
  assign new_U5495 = ~new_U4240 | ~new_U3425;
  assign new_U5496 = ~new_U2427 | ~new_U5494;
  assign new_U5497 = ~new_U5496 | ~new_U5495;
  assign new_U5498 = ~INSTQUEUERD_ADDR_REG_2_ | ~new_U3262;
  assign new_U5499 = ~new_U3388;
  assign new_U5500 = ~new_R2182_U42 | ~new_U7497;
  assign new_U5501 = ~new_U4202 | ~new_U3443;
  assign new_U5502 = ~new_U3737 | ~new_U5500;
  assign new_U5503 = ~new_U2446 | ~new_U3457;
  assign new_U5504 = ~new_U4240 | ~new_U3388;
  assign new_U5505 = ~new_U2427 | ~new_U5502;
  assign new_U5506 = ~new_U5504 | ~new_U5505 | ~new_U5503;
  assign new_U5507 = ~new_U3389;
  assign new_U5508 = ~new_U2431 | ~new_U4237;
  assign new_U5509 = ~new_U3279 | ~new_U5508;
  assign new_U5510 = ~new_U5507 | ~new_U5509;
  assign new_U5511 = ~new_R2182_U33 | ~new_U7497;
  assign new_U5512 = ~new_U4202 | ~new_U3252;
  assign new_U5513 = ~new_U3738 | ~new_U5511;
  assign new_U5514 = ~new_U7700 | ~new_U2446;
  assign new_U5515 = ~new_U5507 | ~new_U4240;
  assign new_U5516 = ~new_U2427 | ~new_U5513;
  assign new_U5517 = ~new_U5515 | ~new_U5516 | ~new_U5514;
  assign new_U5518 = ~new_R2182_U34 | ~new_U7497;
  assign new_U5519 = ~new_U4163 | ~new_U5518;
  assign new_U5520 = ~new_U4240 | ~new_U3253;
  assign new_U5521 = ~new_U2427 | ~new_U5519;
  assign new_U5522 = ~new_U7703 | ~STATE2_REG_1_;
  assign new_U5523 = ~new_U5520 | ~new_U5521 | ~new_U5522;
  assign new_U5524 = ~new_LT_589_U6 | ~new_U2428 | ~STATE2_REG_0_;
  assign new_U5525 = ~new_U3391;
  assign new_U5526 = ~STATE2_REG_1_ | ~new_U3283;
  assign new_U5527 = ~new_U4515 | ~new_U3441;
  assign new_U5528 = ~new_U3345 | ~new_U5527;
  assign new_U5529 = ~new_U3346 | ~new_U5528;
  assign new_U5530 = ~new_U2388 | ~new_U5529;
  assign new_U5531 = ~new_R2182_U25 | ~new_U5526;
  assign new_U5532 = ~new_U4214 | ~new_R2144_U8;
  assign new_U5533 = ~new_U3739 | ~new_U5530;
  assign new_U5534 = ~new_U2388 | ~new_U7721;
  assign new_U5535 = ~new_R2182_U42 | ~new_U5526;
  assign new_U5536 = ~new_U4214 | ~new_R2144_U49;
  assign new_U5537 = ~new_U3740 | ~new_U5534;
  assign new_U5538 = ~new_U3313 | ~new_U3320;
  assign new_U5539 = ~new_U2388 | ~new_U5538;
  assign new_U5540 = ~new_R2182_U33 | ~new_U5526;
  assign new_U5541 = ~new_U4214 | ~new_R2144_U50;
  assign new_U5542 = ~new_U3741 | ~new_U5539;
  assign new_U5543 = ~new_R2182_U34 | ~new_U5526;
  assign new_U5544 = ~new_R2144_U43 | ~new_U4197;
  assign new_U5545 = ~new_U4233 | ~new_U5543 | ~new_U5544;
  assign new_U5546 = ~new_U4465 | ~new_U3259;
  assign new_U5547 = ~new_U4248 | ~new_U2431;
  assign new_U5548 = ~new_U7730 | ~new_U7731 | ~new_U2518 | ~new_U5547;
  assign new_U5549 = ~new_U4180 | ~new_U4223 | ~new_U4491;
  assign new_U5550 = ~new_U2368 | ~new_U5548;
  assign new_U5551 = ~new_U4191 | ~new_U3250;
  assign new_U5552 = ~new_U3401;
  assign new_U5553 = ~new_U4250 | ~new_U4196;
  assign new_U5554 = ~new_U4244 | ~new_U2389;
  assign new_U5555 = ~new_U4254 | ~new_U4238;
  assign new_U5556 = ~new_U4252 | ~new_U4482;
  assign new_U5557 = ~new_U3746 | ~new_U2519;
  assign new_U5558 = ~new_R2099_U86 | ~new_U2380;
  assign new_U5559 = ~new_R2027_U5 | ~new_U2378;
  assign new_U5560 = ~new_R2278_U17 | ~new_U2377;
  assign new_U5561 = ~new_ADD_405_U4 | ~new_U2375;
  assign new_U5562 = ~INSTADDRPOINTER_REG_0_ | ~new_U2374;
  assign new_U5563 = ~REIP_REG_0_ | ~new_U2370;
  assign new_U5564 = ~new_U5552 | ~INSTADDRPOINTER_REG_0_;
  assign new_U5565 = ~new_R2099_U87 | ~new_U2380;
  assign new_U5566 = ~new_R2027_U71 | ~new_U2378;
  assign new_U5567 = ~new_R2278_U42 | ~new_U2377;
  assign new_U5568 = ~new_ADD_405_U81 | ~new_U2375;
  assign new_U5569 = ~new_ADD_515_U4 | ~new_U2374;
  assign new_U5570 = ~new_U2370 | ~REIP_REG_1_;
  assign new_U5571 = ~new_U5552 | ~INSTADDRPOINTER_REG_1_;
  assign new_U5572 = ~new_R2099_U138 | ~new_U2380;
  assign new_U5573 = ~new_R2027_U60 | ~new_U2378;
  assign new_U5574 = ~new_R2278_U101 | ~new_U2377;
  assign new_U5575 = ~new_ADD_405_U5 | ~new_U2375;
  assign new_U5576 = ~new_ADD_515_U71 | ~new_U2374;
  assign new_U5577 = ~new_U2370 | ~REIP_REG_2_;
  assign new_U5578 = ~INSTADDRPOINTER_REG_2_ | ~new_U5552;
  assign new_U5579 = ~new_R2099_U42 | ~new_U2380;
  assign new_U5580 = ~new_R2027_U57 | ~new_U2378;
  assign new_U5581 = ~new_R2278_U92 | ~new_U2377;
  assign new_U5582 = ~new_ADD_405_U93 | ~new_U2375;
  assign new_U5583 = ~new_ADD_515_U68 | ~new_U2374;
  assign new_U5584 = ~new_U2370 | ~REIP_REG_3_;
  assign new_U5585 = ~INSTADDRPOINTER_REG_3_ | ~new_U5552;
  assign new_U5586 = ~new_R2099_U41 | ~new_U2380;
  assign new_U5587 = ~new_R2027_U56 | ~new_U2378;
  assign new_U5588 = ~new_R2278_U89 | ~new_U2377;
  assign new_U5589 = ~new_ADD_405_U68 | ~new_U2375;
  assign new_U5590 = ~new_ADD_515_U67 | ~new_U2374;
  assign new_U5591 = ~new_U2370 | ~REIP_REG_4_;
  assign new_U5592 = ~INSTADDRPOINTER_REG_4_ | ~new_U5552;
  assign new_U5593 = ~new_R2099_U40 | ~new_U2380;
  assign new_U5594 = ~new_R2027_U55 | ~new_U2378;
  assign new_U5595 = ~new_R2278_U86 | ~new_U2377;
  assign new_U5596 = ~new_ADD_405_U67 | ~new_U2375;
  assign new_U5597 = ~new_ADD_515_U66 | ~new_U2374;
  assign new_U5598 = ~new_U2370 | ~REIP_REG_5_;
  assign new_U5599 = ~INSTADDRPOINTER_REG_5_ | ~new_U5552;
  assign new_U5600 = ~new_R2099_U39 | ~new_U2380;
  assign new_U5601 = ~new_R2027_U54 | ~new_U2378;
  assign new_U5602 = ~new_R2278_U83 | ~new_U2377;
  assign new_U5603 = ~new_ADD_405_U66 | ~new_U2375;
  assign new_U5604 = ~new_ADD_515_U65 | ~new_U2374;
  assign new_U5605 = ~new_U2370 | ~REIP_REG_6_;
  assign new_U5606 = ~INSTADDRPOINTER_REG_6_ | ~new_U5552;
  assign new_U5607 = ~new_R2099_U38 | ~new_U2380;
  assign new_U5608 = ~new_R2027_U53 | ~new_U2378;
  assign new_U5609 = ~new_R2278_U80 | ~new_U2377;
  assign new_U5610 = ~new_ADD_405_U65 | ~new_U2375;
  assign new_U5611 = ~new_ADD_515_U64 | ~new_U2374;
  assign new_U5612 = ~new_U2370 | ~REIP_REG_7_;
  assign new_U5613 = ~INSTADDRPOINTER_REG_7_ | ~new_U5552;
  assign new_U5614 = ~new_R2099_U37 | ~new_U2380;
  assign new_U5615 = ~new_R2027_U52 | ~new_U2378;
  assign new_U5616 = ~new_R2278_U77 | ~new_U2377;
  assign new_U5617 = ~new_ADD_405_U64 | ~new_U2375;
  assign new_U5618 = ~new_ADD_515_U63 | ~new_U2374;
  assign new_U5619 = ~new_U2370 | ~REIP_REG_8_;
  assign new_U5620 = ~INSTADDRPOINTER_REG_8_ | ~new_U5552;
  assign new_U5621 = ~new_R2099_U36 | ~new_U2380;
  assign new_U5622 = ~new_R2027_U51 | ~new_U2378;
  assign new_U5623 = ~new_R2278_U74 | ~new_U2377;
  assign new_U5624 = ~new_ADD_405_U63 | ~new_U2375;
  assign new_U5625 = ~new_ADD_515_U62 | ~new_U2374;
  assign new_U5626 = ~new_U2370 | ~REIP_REG_9_;
  assign new_U5627 = ~INSTADDRPOINTER_REG_9_ | ~new_U5552;
  assign new_U5628 = ~new_R2099_U85 | ~new_U2380;
  assign new_U5629 = ~new_R2027_U81 | ~new_U2378;
  assign new_U5630 = ~new_R2278_U160 | ~new_U2377;
  assign new_U5631 = ~new_ADD_405_U91 | ~new_U2375;
  assign new_U5632 = ~new_ADD_515_U91 | ~new_U2374;
  assign new_U5633 = ~new_U2370 | ~REIP_REG_10_;
  assign new_U5634 = ~INSTADDRPOINTER_REG_10_ | ~new_U5552;
  assign new_U5635 = ~new_R2099_U84 | ~new_U2380;
  assign new_U5636 = ~new_R2027_U80 | ~new_U2378;
  assign new_U5637 = ~new_R2278_U157 | ~new_U2377;
  assign new_U5638 = ~new_ADD_405_U90 | ~new_U2375;
  assign new_U5639 = ~new_ADD_515_U90 | ~new_U2374;
  assign new_U5640 = ~new_U2370 | ~REIP_REG_11_;
  assign new_U5641 = ~INSTADDRPOINTER_REG_11_ | ~new_U5552;
  assign new_U5642 = ~new_R2099_U83 | ~new_U2380;
  assign new_U5643 = ~new_R2027_U79 | ~new_U2378;
  assign new_U5644 = ~new_R2278_U154 | ~new_U2377;
  assign new_U5645 = ~new_ADD_405_U89 | ~new_U2375;
  assign new_U5646 = ~new_ADD_515_U89 | ~new_U2374;
  assign new_U5647 = ~new_U2370 | ~REIP_REG_12_;
  assign new_U5648 = ~INSTADDRPOINTER_REG_12_ | ~new_U5552;
  assign new_U5649 = ~new_R2099_U82 | ~new_U2380;
  assign new_U5650 = ~new_R2027_U78 | ~new_U2378;
  assign new_U5651 = ~new_R2278_U151 | ~new_U2377;
  assign new_U5652 = ~new_ADD_405_U88 | ~new_U2375;
  assign new_U5653 = ~new_ADD_515_U88 | ~new_U2374;
  assign new_U5654 = ~new_U2370 | ~REIP_REG_13_;
  assign new_U5655 = ~INSTADDRPOINTER_REG_13_ | ~new_U5552;
  assign new_U5656 = ~new_R2099_U81 | ~new_U2380;
  assign new_U5657 = ~new_R2027_U77 | ~new_U2378;
  assign new_U5658 = ~new_R2278_U148 | ~new_U2377;
  assign new_U5659 = ~new_ADD_405_U87 | ~new_U2375;
  assign new_U5660 = ~new_ADD_515_U87 | ~new_U2374;
  assign new_U5661 = ~new_U2370 | ~REIP_REG_14_;
  assign new_U5662 = ~INSTADDRPOINTER_REG_14_ | ~new_U5552;
  assign new_U5663 = ~new_R2099_U80 | ~new_U2380;
  assign new_U5664 = ~new_R2027_U76 | ~new_U2378;
  assign new_U5665 = ~new_R2278_U145 | ~new_U2377;
  assign new_U5666 = ~new_ADD_405_U86 | ~new_U2375;
  assign new_U5667 = ~new_ADD_515_U86 | ~new_U2374;
  assign new_U5668 = ~new_U2370 | ~REIP_REG_15_;
  assign new_U5669 = ~INSTADDRPOINTER_REG_15_ | ~new_U5552;
  assign new_U5670 = ~new_R2099_U79 | ~new_U2380;
  assign new_U5671 = ~new_R2027_U75 | ~new_U2378;
  assign new_U5672 = ~new_R2278_U142 | ~new_U2377;
  assign new_U5673 = ~new_ADD_405_U85 | ~new_U2375;
  assign new_U5674 = ~new_ADD_515_U85 | ~new_U2374;
  assign new_U5675 = ~new_U2370 | ~REIP_REG_16_;
  assign new_U5676 = ~INSTADDRPOINTER_REG_16_ | ~new_U5552;
  assign new_U5677 = ~new_R2099_U78 | ~new_U2380;
  assign new_U5678 = ~new_R2027_U74 | ~new_U2378;
  assign new_U5679 = ~new_R2278_U139 | ~new_U2377;
  assign new_U5680 = ~new_ADD_405_U84 | ~new_U2375;
  assign new_U5681 = ~new_ADD_515_U84 | ~new_U2374;
  assign new_U5682 = ~new_U2370 | ~REIP_REG_17_;
  assign new_U5683 = ~INSTADDRPOINTER_REG_17_ | ~new_U5552;
  assign new_U5684 = ~new_R2099_U77 | ~new_U2380;
  assign new_U5685 = ~new_R2027_U73 | ~new_U2378;
  assign new_U5686 = ~new_R2278_U136 | ~new_U2377;
  assign new_U5687 = ~new_ADD_405_U83 | ~new_U2375;
  assign new_U5688 = ~new_ADD_515_U83 | ~new_U2374;
  assign new_U5689 = ~new_U2370 | ~REIP_REG_18_;
  assign new_U5690 = ~INSTADDRPOINTER_REG_18_ | ~new_U5552;
  assign new_U5691 = ~new_R2099_U76 | ~new_U2380;
  assign new_U5692 = ~new_R2027_U72 | ~new_U2378;
  assign new_U5693 = ~new_R2278_U133 | ~new_U2377;
  assign new_U5694 = ~new_ADD_405_U82 | ~new_U2375;
  assign new_U5695 = ~new_ADD_515_U82 | ~new_U2374;
  assign new_U5696 = ~new_U2370 | ~REIP_REG_19_;
  assign new_U5697 = ~INSTADDRPOINTER_REG_19_ | ~new_U5552;
  assign new_U5698 = ~new_R2099_U75 | ~new_U2380;
  assign new_U5699 = ~new_R2027_U70 | ~new_U2378;
  assign new_U5700 = ~new_R2278_U129 | ~new_U2377;
  assign new_U5701 = ~new_ADD_405_U80 | ~new_U2375;
  assign new_U5702 = ~new_ADD_515_U81 | ~new_U2374;
  assign new_U5703 = ~new_U2370 | ~REIP_REG_20_;
  assign new_U5704 = ~INSTADDRPOINTER_REG_20_ | ~new_U5552;
  assign new_U5705 = ~new_R2099_U74 | ~new_U2380;
  assign new_U5706 = ~new_R2027_U69 | ~new_U2378;
  assign new_U5707 = ~new_R2278_U126 | ~new_U2377;
  assign new_U5708 = ~new_ADD_405_U79 | ~new_U2375;
  assign new_U5709 = ~new_ADD_515_U80 | ~new_U2374;
  assign new_U5710 = ~new_U2370 | ~REIP_REG_21_;
  assign new_U5711 = ~INSTADDRPOINTER_REG_21_ | ~new_U5552;
  assign new_U5712 = ~new_R2099_U73 | ~new_U2380;
  assign new_U5713 = ~new_R2027_U68 | ~new_U2378;
  assign new_U5714 = ~new_R2278_U123 | ~new_U2377;
  assign new_U5715 = ~new_ADD_405_U78 | ~new_U2375;
  assign new_U5716 = ~new_ADD_515_U79 | ~new_U2374;
  assign new_U5717 = ~new_U2370 | ~REIP_REG_22_;
  assign new_U5718 = ~INSTADDRPOINTER_REG_22_ | ~new_U5552;
  assign new_U5719 = ~new_R2099_U72 | ~new_U2380;
  assign new_U5720 = ~new_R2027_U67 | ~new_U2378;
  assign new_U5721 = ~new_R2278_U120 | ~new_U2377;
  assign new_U5722 = ~new_ADD_405_U77 | ~new_U2375;
  assign new_U5723 = ~new_ADD_515_U78 | ~new_U2374;
  assign new_U5724 = ~new_U2370 | ~REIP_REG_23_;
  assign new_U5725 = ~INSTADDRPOINTER_REG_23_ | ~new_U5552;
  assign new_U5726 = ~new_R2099_U71 | ~new_U2380;
  assign new_U5727 = ~new_R2027_U66 | ~new_U2378;
  assign new_U5728 = ~new_R2278_U117 | ~new_U2377;
  assign new_U5729 = ~new_ADD_405_U76 | ~new_U2375;
  assign new_U5730 = ~new_ADD_515_U77 | ~new_U2374;
  assign new_U5731 = ~new_U2370 | ~REIP_REG_24_;
  assign new_U5732 = ~INSTADDRPOINTER_REG_24_ | ~new_U5552;
  assign new_U5733 = ~new_R2099_U70 | ~new_U2380;
  assign new_U5734 = ~new_R2027_U65 | ~new_U2378;
  assign new_U5735 = ~new_R2278_U114 | ~new_U2377;
  assign new_U5736 = ~new_ADD_405_U75 | ~new_U2375;
  assign new_U5737 = ~new_ADD_515_U76 | ~new_U2374;
  assign new_U5738 = ~new_U2370 | ~REIP_REG_25_;
  assign new_U5739 = ~INSTADDRPOINTER_REG_25_ | ~new_U5552;
  assign new_U5740 = ~new_R2099_U69 | ~new_U2380;
  assign new_U5741 = ~new_R2027_U64 | ~new_U2378;
  assign new_U5742 = ~new_R2278_U111 | ~new_U2377;
  assign new_U5743 = ~new_ADD_405_U74 | ~new_U2375;
  assign new_U5744 = ~new_ADD_515_U75 | ~new_U2374;
  assign new_U5745 = ~new_U2370 | ~REIP_REG_26_;
  assign new_U5746 = ~INSTADDRPOINTER_REG_26_ | ~new_U5552;
  assign new_U5747 = ~new_R2099_U68 | ~new_U2380;
  assign new_U5748 = ~new_R2027_U63 | ~new_U2378;
  assign new_U5749 = ~new_R2278_U108 | ~new_U2377;
  assign new_U5750 = ~new_ADD_405_U73 | ~new_U2375;
  assign new_U5751 = ~new_ADD_515_U74 | ~new_U2374;
  assign new_U5752 = ~new_U2370 | ~REIP_REG_27_;
  assign new_U5753 = ~INSTADDRPOINTER_REG_27_ | ~new_U5552;
  assign new_U5754 = ~new_R2099_U67 | ~new_U2380;
  assign new_U5755 = ~new_R2027_U62 | ~new_U2378;
  assign new_U5756 = ~new_R2278_U105 | ~new_U2377;
  assign new_U5757 = ~new_ADD_405_U72 | ~new_U2375;
  assign new_U5758 = ~new_ADD_515_U73 | ~new_U2374;
  assign new_U5759 = ~new_U2370 | ~REIP_REG_28_;
  assign new_U5760 = ~INSTADDRPOINTER_REG_28_ | ~new_U5552;
  assign new_U5761 = ~new_R2099_U66 | ~new_U2380;
  assign new_U5762 = ~new_R2027_U61 | ~new_U2378;
  assign new_U5763 = ~new_R2278_U103 | ~new_U2377;
  assign new_U5764 = ~new_ADD_405_U71 | ~new_U2375;
  assign new_U5765 = ~new_ADD_515_U72 | ~new_U2374;
  assign new_U5766 = ~new_U2370 | ~REIP_REG_29_;
  assign new_U5767 = ~INSTADDRPOINTER_REG_29_ | ~new_U5552;
  assign new_U5768 = ~new_R2099_U65 | ~new_U2380;
  assign new_U5769 = ~new_R2027_U59 | ~new_U2378;
  assign new_U5770 = ~new_R2278_U98 | ~new_U2377;
  assign new_U5771 = ~new_ADD_405_U70 | ~new_U2375;
  assign new_U5772 = ~new_ADD_515_U70 | ~new_U2374;
  assign new_U5773 = ~new_U2370 | ~REIP_REG_30_;
  assign new_U5774 = ~INSTADDRPOINTER_REG_30_ | ~new_U5552;
  assign new_U5775 = ~new_R2099_U64 | ~new_U2380;
  assign new_U5776 = ~new_R2027_U58 | ~new_U2378;
  assign new_U5777 = ~new_R2278_U96 | ~new_U2377;
  assign new_U5778 = ~new_ADD_405_U69 | ~new_U2375;
  assign new_U5779 = ~new_ADD_515_U69 | ~new_U2374;
  assign new_U5780 = ~new_U2370 | ~REIP_REG_31_;
  assign new_U5781 = ~INSTADDRPOINTER_REG_31_ | ~new_U5552;
  assign new_U5782 = ~new_U4197 | ~new_U3281;
  assign new_U5783 = ~new_U3403;
  assign new_U5784 = ~STATE2_REG_2_ | ~new_U3281;
  assign new_U5785 = ~STATE2_REG_1_ | ~new_U3295;
  assign new_U5786 = ~new_U5785 | ~new_U5784;
  assign new_U5787 = ~PHYADDRPOINTER_REG_0_ | ~new_U2376;
  assign new_U5788 = ~new_U2372 | ~new_R2278_U17;
  assign new_U5789 = ~new_U2365 | ~REIP_REG_0_;
  assign new_U5790 = ~new_R2358_U82 | ~new_U2364;
  assign new_U5791 = ~PHYADDRPOINTER_REG_0_ | ~new_U5783;
  assign new_U5792 = ~new_R2337_U5 | ~new_U2376;
  assign new_U5793 = ~new_U2372 | ~new_R2278_U42;
  assign new_U5794 = ~new_U2365 | ~REIP_REG_1_;
  assign new_U5795 = ~new_R2358_U112 | ~new_U2364;
  assign new_U5796 = ~PHYADDRPOINTER_REG_1_ | ~new_U5783;
  assign new_U5797 = ~new_R2337_U60 | ~new_U2376;
  assign new_U5798 = ~new_U2372 | ~new_R2278_U101;
  assign new_U5799 = ~new_U2365 | ~REIP_REG_2_;
  assign new_U5800 = ~new_R2358_U19 | ~new_U2364;
  assign new_U5801 = ~PHYADDRPOINTER_REG_2_ | ~new_U5783;
  assign new_U5802 = ~new_R2337_U57 | ~new_U2376;
  assign new_U5803 = ~new_U2372 | ~new_R2278_U92;
  assign new_U5804 = ~new_U2365 | ~REIP_REG_3_;
  assign new_U5805 = ~new_R2358_U20 | ~new_U2364;
  assign new_U5806 = ~PHYADDRPOINTER_REG_3_ | ~new_U5783;
  assign new_U5807 = ~new_R2337_U56 | ~new_U2376;
  assign new_U5808 = ~new_U2372 | ~new_R2278_U89;
  assign new_U5809 = ~new_U2365 | ~REIP_REG_4_;
  assign new_U5810 = ~new_R2358_U90 | ~new_U2364;
  assign new_U5811 = ~PHYADDRPOINTER_REG_4_ | ~new_U5783;
  assign new_U5812 = ~new_R2337_U55 | ~new_U2376;
  assign new_U5813 = ~new_U2372 | ~new_R2278_U86;
  assign new_U5814 = ~new_U2365 | ~REIP_REG_5_;
  assign new_U5815 = ~new_R2358_U88 | ~new_U2364;
  assign new_U5816 = ~PHYADDRPOINTER_REG_5_ | ~new_U5783;
  assign new_U5817 = ~new_R2337_U54 | ~new_U2376;
  assign new_U5818 = ~new_U2372 | ~new_R2278_U83;
  assign new_U5819 = ~new_U2365 | ~REIP_REG_6_;
  assign new_U5820 = ~new_R2358_U86 | ~new_U2364;
  assign new_U5821 = ~PHYADDRPOINTER_REG_6_ | ~new_U5783;
  assign new_U5822 = ~new_R2337_U53 | ~new_U2376;
  assign new_U5823 = ~new_U2372 | ~new_R2278_U80;
  assign new_U5824 = ~new_U2365 | ~REIP_REG_7_;
  assign new_U5825 = ~new_R2358_U21 | ~new_U2364;
  assign new_U5826 = ~PHYADDRPOINTER_REG_7_ | ~new_U5783;
  assign new_U5827 = ~new_R2337_U52 | ~new_U2376;
  assign new_U5828 = ~new_U2372 | ~new_R2278_U77;
  assign new_U5829 = ~new_U2365 | ~REIP_REG_8_;
  assign new_U5830 = ~new_R2358_U85 | ~new_U2364;
  assign new_U5831 = ~PHYADDRPOINTER_REG_8_ | ~new_U5783;
  assign new_U5832 = ~new_R2337_U51 | ~new_U2376;
  assign new_U5833 = ~new_U2372 | ~new_R2278_U74;
  assign new_U5834 = ~new_U2365 | ~REIP_REG_9_;
  assign new_U5835 = ~new_R2358_U83 | ~new_U2364;
  assign new_U5836 = ~PHYADDRPOINTER_REG_9_ | ~new_U5783;
  assign new_U5837 = ~new_R2337_U80 | ~new_U2376;
  assign new_U5838 = ~new_U2372 | ~new_R2278_U160;
  assign new_U5839 = ~new_U2365 | ~REIP_REG_10_;
  assign new_U5840 = ~new_R2358_U14 | ~new_U2364;
  assign new_U5841 = ~PHYADDRPOINTER_REG_10_ | ~new_U5783;
  assign new_U5842 = ~new_R2337_U79 | ~new_U2376;
  assign new_U5843 = ~new_U2372 | ~new_R2278_U157;
  assign new_U5844 = ~new_U2365 | ~REIP_REG_11_;
  assign new_U5845 = ~new_R2358_U15 | ~new_U2364;
  assign new_U5846 = ~PHYADDRPOINTER_REG_11_ | ~new_U5783;
  assign new_U5847 = ~new_R2337_U78 | ~new_U2376;
  assign new_U5848 = ~new_U2372 | ~new_R2278_U154;
  assign new_U5849 = ~new_U2365 | ~REIP_REG_12_;
  assign new_U5850 = ~new_R2358_U122 | ~new_U2364;
  assign new_U5851 = ~PHYADDRPOINTER_REG_12_ | ~new_U5783;
  assign new_U5852 = ~new_R2337_U77 | ~new_U2376;
  assign new_U5853 = ~new_U2372 | ~new_R2278_U151;
  assign new_U5854 = ~new_U2365 | ~REIP_REG_13_;
  assign new_U5855 = ~new_R2358_U120 | ~new_U2364;
  assign new_U5856 = ~PHYADDRPOINTER_REG_13_ | ~new_U5783;
  assign new_U5857 = ~new_R2337_U76 | ~new_U2376;
  assign new_U5858 = ~new_U2372 | ~new_R2278_U148;
  assign new_U5859 = ~new_U2365 | ~REIP_REG_14_;
  assign new_U5860 = ~new_R2358_U119 | ~new_U2364;
  assign new_U5861 = ~PHYADDRPOINTER_REG_14_ | ~new_U5783;
  assign new_U5862 = ~new_R2337_U75 | ~new_U2376;
  assign new_U5863 = ~new_U2372 | ~new_R2278_U145;
  assign new_U5864 = ~new_U2365 | ~REIP_REG_15_;
  assign new_U5865 = ~new_R2358_U16 | ~new_U2364;
  assign new_U5866 = ~PHYADDRPOINTER_REG_15_ | ~new_U5783;
  assign new_U5867 = ~new_R2337_U74 | ~new_U2376;
  assign new_U5868 = ~new_U2372 | ~new_R2278_U142;
  assign new_U5869 = ~new_U2365 | ~REIP_REG_16_;
  assign new_U5870 = ~new_R2358_U17 | ~new_U2364;
  assign new_U5871 = ~PHYADDRPOINTER_REG_16_ | ~new_U5783;
  assign new_U5872 = ~new_R2337_U73 | ~new_U2376;
  assign new_U5873 = ~new_U2372 | ~new_R2278_U139;
  assign new_U5874 = ~new_U2365 | ~REIP_REG_17_;
  assign new_U5875 = ~new_R2358_U118 | ~new_U2364;
  assign new_U5876 = ~PHYADDRPOINTER_REG_17_ | ~new_U5783;
  assign new_U5877 = ~new_R2337_U72 | ~new_U2376;
  assign new_U5878 = ~new_U2372 | ~new_R2278_U136;
  assign new_U5879 = ~new_U2365 | ~REIP_REG_18_;
  assign new_U5880 = ~new_R2358_U116 | ~new_U2364;
  assign new_U5881 = ~PHYADDRPOINTER_REG_18_ | ~new_U5783;
  assign new_U5882 = ~new_R2337_U71 | ~new_U2376;
  assign new_U5883 = ~new_U2372 | ~new_R2278_U133;
  assign new_U5884 = ~new_U2365 | ~REIP_REG_19_;
  assign new_U5885 = ~new_R2358_U114 | ~new_U2364;
  assign new_U5886 = ~PHYADDRPOINTER_REG_19_ | ~new_U5783;
  assign new_U5887 = ~new_R2337_U70 | ~new_U2376;
  assign new_U5888 = ~new_U2372 | ~new_R2278_U129;
  assign new_U5889 = ~new_U2365 | ~REIP_REG_20_;
  assign new_U5890 = ~new_R2358_U110 | ~new_U2364;
  assign new_U5891 = ~PHYADDRPOINTER_REG_20_ | ~new_U5783;
  assign new_U5892 = ~new_R2337_U69 | ~new_U2376;
  assign new_U5893 = ~new_U2372 | ~new_R2278_U126;
  assign new_U5894 = ~new_U2365 | ~REIP_REG_21_;
  assign new_U5895 = ~new_R2358_U18 | ~new_U2364;
  assign new_U5896 = ~PHYADDRPOINTER_REG_21_ | ~new_U5783;
  assign new_U5897 = ~new_R2337_U68 | ~new_U2376;
  assign new_U5898 = ~new_U2372 | ~new_R2278_U123;
  assign new_U5899 = ~new_U2365 | ~REIP_REG_22_;
  assign new_U5900 = ~new_R2358_U109 | ~new_U2364;
  assign new_U5901 = ~PHYADDRPOINTER_REG_22_ | ~new_U5783;
  assign new_U5902 = ~new_R2337_U67 | ~new_U2376;
  assign new_U5903 = ~new_U2372 | ~new_R2278_U120;
  assign new_U5904 = ~new_U2365 | ~REIP_REG_23_;
  assign new_U5905 = ~new_R2358_U107 | ~new_U2364;
  assign new_U5906 = ~PHYADDRPOINTER_REG_23_ | ~new_U5783;
  assign new_U5907 = ~new_R2337_U66 | ~new_U2376;
  assign new_U5908 = ~new_U2372 | ~new_R2278_U117;
  assign new_U5909 = ~new_U2365 | ~REIP_REG_24_;
  assign new_U5910 = ~new_R2358_U105 | ~new_U2364;
  assign new_U5911 = ~PHYADDRPOINTER_REG_24_ | ~new_U5783;
  assign new_U5912 = ~new_R2337_U65 | ~new_U2376;
  assign new_U5913 = ~new_U2372 | ~new_R2278_U114;
  assign new_U5914 = ~new_U2365 | ~REIP_REG_25_;
  assign new_U5915 = ~new_R2358_U103 | ~new_U2364;
  assign new_U5916 = ~PHYADDRPOINTER_REG_25_ | ~new_U5783;
  assign new_U5917 = ~new_R2337_U64 | ~new_U2376;
  assign new_U5918 = ~new_U2372 | ~new_R2278_U111;
  assign new_U5919 = ~new_U2365 | ~REIP_REG_26_;
  assign new_U5920 = ~new_R2358_U101 | ~new_U2364;
  assign new_U5921 = ~PHYADDRPOINTER_REG_26_ | ~new_U5783;
  assign new_U5922 = ~new_R2337_U63 | ~new_U2376;
  assign new_U5923 = ~new_U2372 | ~new_R2278_U108;
  assign new_U5924 = ~new_U2365 | ~REIP_REG_27_;
  assign new_U5925 = ~new_R2358_U99 | ~new_U2364;
  assign new_U5926 = ~PHYADDRPOINTER_REG_27_ | ~new_U5783;
  assign new_U5927 = ~new_R2337_U62 | ~new_U2376;
  assign new_U5928 = ~new_U2372 | ~new_R2278_U105;
  assign new_U5929 = ~new_U2365 | ~REIP_REG_28_;
  assign new_U5930 = ~new_R2358_U97 | ~new_U2364;
  assign new_U5931 = ~PHYADDRPOINTER_REG_28_ | ~new_U5783;
  assign new_U5932 = ~new_R2337_U61 | ~new_U2376;
  assign new_U5933 = ~new_U2372 | ~new_R2278_U103;
  assign new_U5934 = ~new_U2365 | ~REIP_REG_29_;
  assign new_U5935 = ~new_R2358_U95 | ~new_U2364;
  assign new_U5936 = ~PHYADDRPOINTER_REG_29_ | ~new_U5783;
  assign new_U5937 = ~new_R2337_U59 | ~new_U2376;
  assign new_U5938 = ~new_U2372 | ~new_R2278_U98;
  assign new_U5939 = ~new_U2365 | ~REIP_REG_30_;
  assign new_U5940 = ~new_R2358_U93 | ~new_U2364;
  assign new_U5941 = ~PHYADDRPOINTER_REG_30_ | ~new_U5783;
  assign new_U5942 = ~new_R2337_U58 | ~new_U2376;
  assign new_U5943 = ~new_U2372 | ~new_R2278_U96;
  assign new_U5944 = ~new_U2365 | ~REIP_REG_31_;
  assign new_U5945 = ~new_R2358_U91 | ~new_U2364;
  assign new_U5946 = ~PHYADDRPOINTER_REG_31_ | ~new_U5783;
  assign new_U5947 = ~READY_N | ~new_U3269;
  assign new_U5948 = ~EAX_REG_15_ | ~new_U2382;
  assign new_U5949 = ~DATAI_15_ | ~new_U2381;
  assign new_U5950 = ~new_U5949 | ~new_U5948;
  assign new_U5951 = ~EAX_REG_14_ | ~new_U2382;
  assign new_U5952 = ~DATAI_14_ | ~new_U2381;
  assign new_U5953 = ~new_U5952 | ~new_U5951;
  assign new_U5954 = ~EAX_REG_13_ | ~new_U2382;
  assign new_U5955 = ~DATAI_13_ | ~new_U2381;
  assign new_U5956 = ~new_U5955 | ~new_U5954;
  assign new_U5957 = ~EAX_REG_12_ | ~new_U2382;
  assign new_U5958 = ~DATAI_12_ | ~new_U2381;
  assign new_U5959 = ~new_U5958 | ~new_U5957;
  assign new_U5960 = ~EAX_REG_11_ | ~new_U2382;
  assign new_U5961 = ~DATAI_11_ | ~new_U2381;
  assign new_U5962 = ~new_U5961 | ~new_U5960;
  assign new_U5963 = ~EAX_REG_10_ | ~new_U2382;
  assign new_U5964 = ~DATAI_10_ | ~new_U2381;
  assign new_U5965 = ~new_U5964 | ~new_U5963;
  assign new_U5966 = ~EAX_REG_9_ | ~new_U2382;
  assign new_U5967 = ~DATAI_9_ | ~new_U2381;
  assign new_U5968 = ~new_U5967 | ~new_U5966;
  assign new_U5969 = ~EAX_REG_8_ | ~new_U2382;
  assign new_U5970 = ~DATAI_8_ | ~new_U2381;
  assign new_U5971 = ~new_U5970 | ~new_U5969;
  assign new_U5972 = ~EAX_REG_7_ | ~new_U2382;
  assign new_U5973 = ~new_U2381 | ~DATAI_7_;
  assign new_U5974 = ~new_U5973 | ~new_U5972;
  assign new_U5975 = ~EAX_REG_6_ | ~new_U2382;
  assign new_U5976 = ~new_U2381 | ~DATAI_6_;
  assign new_U5977 = ~new_U5976 | ~new_U5975;
  assign new_U5978 = ~EAX_REG_5_ | ~new_U2382;
  assign new_U5979 = ~new_U2381 | ~DATAI_5_;
  assign new_U5980 = ~new_U5979 | ~new_U5978;
  assign new_U5981 = ~EAX_REG_4_ | ~new_U2382;
  assign new_U5982 = ~new_U2381 | ~DATAI_4_;
  assign new_U5983 = ~new_U5982 | ~new_U5981;
  assign new_U5984 = ~EAX_REG_3_ | ~new_U2382;
  assign new_U5985 = ~new_U2381 | ~DATAI_3_;
  assign new_U5986 = ~new_U5985 | ~new_U5984;
  assign new_U5987 = ~EAX_REG_2_ | ~new_U2382;
  assign new_U5988 = ~new_U2381 | ~DATAI_2_;
  assign new_U5989 = ~new_U5988 | ~new_U5987;
  assign new_U5990 = ~EAX_REG_1_ | ~new_U2382;
  assign new_U5991 = ~new_U2381 | ~DATAI_1_;
  assign new_U5992 = ~new_U5991 | ~new_U5990;
  assign new_U5993 = ~EAX_REG_0_ | ~new_U2382;
  assign new_U5994 = ~new_U2381 | ~DATAI_0_;
  assign new_U5995 = ~new_U5994 | ~new_U5993;
  assign new_U5996 = ~EAX_REG_30_ | ~new_U2382;
  assign new_U5997 = ~DATAI_14_ | ~new_U2381;
  assign new_U5998 = ~new_U5997 | ~new_U5996;
  assign new_U5999 = ~EAX_REG_29_ | ~new_U2382;
  assign new_U6000 = ~DATAI_13_ | ~new_U2381;
  assign new_U6001 = ~new_U6000 | ~new_U5999;
  assign new_U6002 = ~EAX_REG_28_ | ~new_U2382;
  assign new_U6003 = ~DATAI_12_ | ~new_U2381;
  assign new_U6004 = ~new_U6003 | ~new_U6002;
  assign new_U6005 = ~EAX_REG_27_ | ~new_U2382;
  assign new_U6006 = ~DATAI_11_ | ~new_U2381;
  assign new_U6007 = ~new_U6006 | ~new_U6005;
  assign new_U6008 = ~EAX_REG_26_ | ~new_U2382;
  assign new_U6009 = ~DATAI_10_ | ~new_U2381;
  assign new_U6010 = ~new_U6009 | ~new_U6008;
  assign new_U6011 = ~EAX_REG_25_ | ~new_U2382;
  assign new_U6012 = ~DATAI_9_ | ~new_U2381;
  assign new_U6013 = ~new_U6012 | ~new_U6011;
  assign new_U6014 = ~EAX_REG_24_ | ~new_U2382;
  assign new_U6015 = ~DATAI_8_ | ~new_U2381;
  assign new_U6016 = ~new_U6015 | ~new_U6014;
  assign new_U6017 = ~EAX_REG_23_ | ~new_U2382;
  assign new_U6018 = ~new_U2381 | ~DATAI_7_;
  assign new_U6019 = ~new_U6018 | ~new_U6017;
  assign new_U6020 = ~EAX_REG_22_ | ~new_U2382;
  assign new_U6021 = ~new_U2381 | ~DATAI_6_;
  assign new_U6022 = ~new_U6021 | ~new_U6020;
  assign new_U6023 = ~EAX_REG_21_ | ~new_U2382;
  assign new_U6024 = ~new_U2381 | ~DATAI_5_;
  assign new_U6025 = ~new_U6024 | ~new_U6023;
  assign new_U6026 = ~EAX_REG_20_ | ~new_U2382;
  assign new_U6027 = ~new_U2381 | ~DATAI_4_;
  assign new_U6028 = ~new_U6027 | ~new_U6026;
  assign new_U6029 = ~EAX_REG_19_ | ~new_U2382;
  assign new_U6030 = ~new_U2381 | ~DATAI_3_;
  assign new_U6031 = ~new_U6030 | ~new_U6029;
  assign new_U6032 = ~EAX_REG_18_ | ~new_U2382;
  assign new_U6033 = ~new_U2381 | ~DATAI_2_;
  assign new_U6034 = ~new_U6033 | ~new_U6032;
  assign new_U6035 = ~EAX_REG_17_ | ~new_U2382;
  assign new_U6036 = ~new_U2381 | ~DATAI_1_;
  assign new_U6037 = ~new_U6036 | ~new_U6035;
  assign new_U6038 = ~EAX_REG_16_ | ~new_U2382;
  assign new_U6039 = ~new_U2381 | ~DATAI_0_;
  assign new_U6040 = ~new_U6039 | ~new_U6038;
  assign new_U6041 = ~new_U4247 | ~new_U4223 | ~new_U7594;
  assign new_U6042 = ~new_U2428 | ~new_U3281;
  assign new_U6043 = ~new_U3404;
  assign new_U6044 = ~new_U2385 | ~LWORD_REG_0_;
  assign new_U6045 = ~new_U2384 | ~EAX_REG_0_;
  assign new_U6046 = ~DATAO_REG_0_ | ~new_U6043;
  assign new_U6047 = ~new_U2385 | ~LWORD_REG_1_;
  assign new_U6048 = ~new_U2384 | ~EAX_REG_1_;
  assign new_U6049 = ~DATAO_REG_1_ | ~new_U6043;
  assign new_U6050 = ~new_U2385 | ~LWORD_REG_2_;
  assign new_U6051 = ~new_U2384 | ~EAX_REG_2_;
  assign new_U6052 = ~DATAO_REG_2_ | ~new_U6043;
  assign new_U6053 = ~new_U2385 | ~LWORD_REG_3_;
  assign new_U6054 = ~new_U2384 | ~EAX_REG_3_;
  assign new_U6055 = ~DATAO_REG_3_ | ~new_U6043;
  assign new_U6056 = ~new_U2385 | ~LWORD_REG_4_;
  assign new_U6057 = ~new_U2384 | ~EAX_REG_4_;
  assign new_U6058 = ~DATAO_REG_4_ | ~new_U6043;
  assign new_U6059 = ~new_U2385 | ~LWORD_REG_5_;
  assign new_U6060 = ~new_U2384 | ~EAX_REG_5_;
  assign new_U6061 = ~DATAO_REG_5_ | ~new_U6043;
  assign new_U6062 = ~new_U2385 | ~LWORD_REG_6_;
  assign new_U6063 = ~new_U2384 | ~EAX_REG_6_;
  assign new_U6064 = ~DATAO_REG_6_ | ~new_U6043;
  assign new_U6065 = ~new_U2385 | ~LWORD_REG_7_;
  assign new_U6066 = ~new_U2384 | ~EAX_REG_7_;
  assign new_U6067 = ~DATAO_REG_7_ | ~new_U6043;
  assign new_U6068 = ~new_U2385 | ~LWORD_REG_8_;
  assign new_U6069 = ~new_U2384 | ~EAX_REG_8_;
  assign new_U6070 = ~DATAO_REG_8_ | ~new_U6043;
  assign new_U6071 = ~new_U2385 | ~LWORD_REG_9_;
  assign new_U6072 = ~new_U2384 | ~EAX_REG_9_;
  assign new_U6073 = ~DATAO_REG_9_ | ~new_U6043;
  assign new_U6074 = ~new_U2385 | ~LWORD_REG_10_;
  assign new_U6075 = ~new_U2384 | ~EAX_REG_10_;
  assign new_U6076 = ~DATAO_REG_10_ | ~new_U6043;
  assign new_U6077 = ~new_U2385 | ~LWORD_REG_11_;
  assign new_U6078 = ~new_U2384 | ~EAX_REG_11_;
  assign new_U6079 = ~DATAO_REG_11_ | ~new_U6043;
  assign new_U6080 = ~new_U2385 | ~LWORD_REG_12_;
  assign new_U6081 = ~new_U2384 | ~EAX_REG_12_;
  assign new_U6082 = ~DATAO_REG_12_ | ~new_U6043;
  assign new_U6083 = ~new_U2385 | ~LWORD_REG_13_;
  assign new_U6084 = ~new_U2384 | ~EAX_REG_13_;
  assign new_U6085 = ~DATAO_REG_13_ | ~new_U6043;
  assign new_U6086 = ~new_U2385 | ~LWORD_REG_14_;
  assign new_U6087 = ~new_U2384 | ~EAX_REG_14_;
  assign new_U6088 = ~DATAO_REG_14_ | ~new_U6043;
  assign new_U6089 = ~new_U2385 | ~LWORD_REG_15_;
  assign new_U6090 = ~new_U2384 | ~EAX_REG_15_;
  assign new_U6091 = ~DATAO_REG_15_ | ~new_U6043;
  assign new_U6092 = ~new_U2424 | ~EAX_REG_16_;
  assign new_U6093 = ~new_U2385 | ~UWORD_REG_0_;
  assign new_U6094 = ~DATAO_REG_16_ | ~new_U6043;
  assign new_U6095 = ~new_U2424 | ~EAX_REG_17_;
  assign new_U6096 = ~new_U2385 | ~UWORD_REG_1_;
  assign new_U6097 = ~DATAO_REG_17_ | ~new_U6043;
  assign new_U6098 = ~new_U2424 | ~EAX_REG_18_;
  assign new_U6099 = ~new_U2385 | ~UWORD_REG_2_;
  assign new_U6100 = ~DATAO_REG_18_ | ~new_U6043;
  assign new_U6101 = ~new_U2424 | ~EAX_REG_19_;
  assign new_U6102 = ~new_U2385 | ~UWORD_REG_3_;
  assign new_U6103 = ~DATAO_REG_19_ | ~new_U6043;
  assign new_U6104 = ~new_U2424 | ~EAX_REG_20_;
  assign new_U6105 = ~new_U2385 | ~UWORD_REG_4_;
  assign new_U6106 = ~DATAO_REG_20_ | ~new_U6043;
  assign new_U6107 = ~new_U2424 | ~EAX_REG_21_;
  assign new_U6108 = ~new_U2385 | ~UWORD_REG_5_;
  assign new_U6109 = ~DATAO_REG_21_ | ~new_U6043;
  assign new_U6110 = ~new_U2424 | ~EAX_REG_22_;
  assign new_U6111 = ~new_U2385 | ~UWORD_REG_6_;
  assign new_U6112 = ~DATAO_REG_22_ | ~new_U6043;
  assign new_U6113 = ~new_U2424 | ~EAX_REG_23_;
  assign new_U6114 = ~new_U2385 | ~UWORD_REG_7_;
  assign new_U6115 = ~DATAO_REG_23_ | ~new_U6043;
  assign new_U6116 = ~new_U2424 | ~EAX_REG_24_;
  assign new_U6117 = ~new_U2385 | ~UWORD_REG_8_;
  assign new_U6118 = ~DATAO_REG_24_ | ~new_U6043;
  assign new_U6119 = ~new_U2424 | ~EAX_REG_25_;
  assign new_U6120 = ~new_U2385 | ~UWORD_REG_9_;
  assign new_U6121 = ~DATAO_REG_25_ | ~new_U6043;
  assign new_U6122 = ~new_U2424 | ~EAX_REG_26_;
  assign new_U6123 = ~new_U2385 | ~UWORD_REG_10_;
  assign new_U6124 = ~DATAO_REG_26_ | ~new_U6043;
  assign new_U6125 = ~new_U2424 | ~EAX_REG_27_;
  assign new_U6126 = ~new_U2385 | ~UWORD_REG_11_;
  assign new_U6127 = ~DATAO_REG_27_ | ~new_U6043;
  assign new_U6128 = ~new_U2424 | ~EAX_REG_28_;
  assign new_U6129 = ~new_U2385 | ~UWORD_REG_12_;
  assign new_U6130 = ~DATAO_REG_28_ | ~new_U6043;
  assign new_U6131 = ~new_U2424 | ~EAX_REG_29_;
  assign new_U6132 = ~new_U2385 | ~UWORD_REG_13_;
  assign new_U6133 = ~DATAO_REG_29_ | ~new_U6043;
  assign new_U6134 = ~new_U2424 | ~EAX_REG_30_;
  assign new_U6135 = ~new_U2385 | ~UWORD_REG_14_;
  assign new_U6136 = ~DATAO_REG_30_ | ~new_U6043;
  assign new_U6137 = ~new_GTE_485_U6 | ~new_U4182 | ~new_U2447;
  assign new_U6138 = ~new_U4182 | ~new_U4242 | ~new_U4185;
  assign new_U6139 = ~new_R2167_U17 | ~new_U4188 | ~new_U3270;
  assign new_U6140 = ~new_U7491 | ~new_U3244;
  assign new_U6141 = ~new_U3871 | ~new_U6140;
  assign new_U6142 = ~new_U2422 | ~DATAI_0_;
  assign new_U6143 = ~new_U2386 | ~new_R2358_U82;
  assign new_U6144 = ~EAX_REG_0_ | ~new_U3411;
  assign new_U6145 = ~new_U2422 | ~DATAI_1_;
  assign new_U6146 = ~new_U2386 | ~new_R2358_U112;
  assign new_U6147 = ~EAX_REG_1_ | ~new_U3411;
  assign new_U6148 = ~new_U2422 | ~DATAI_2_;
  assign new_U6149 = ~new_U2386 | ~new_R2358_U19;
  assign new_U6150 = ~EAX_REG_2_ | ~new_U3411;
  assign new_U6151 = ~new_U2422 | ~DATAI_3_;
  assign new_U6152 = ~new_U2386 | ~new_R2358_U20;
  assign new_U6153 = ~EAX_REG_3_ | ~new_U3411;
  assign new_U6154 = ~new_U2422 | ~DATAI_4_;
  assign new_U6155 = ~new_U2386 | ~new_R2358_U90;
  assign new_U6156 = ~EAX_REG_4_ | ~new_U3411;
  assign new_U6157 = ~new_U2422 | ~DATAI_5_;
  assign new_U6158 = ~new_U2386 | ~new_R2358_U88;
  assign new_U6159 = ~EAX_REG_5_ | ~new_U3411;
  assign new_U6160 = ~new_U2422 | ~DATAI_6_;
  assign new_U6161 = ~new_U2386 | ~new_R2358_U86;
  assign new_U6162 = ~EAX_REG_6_ | ~new_U3411;
  assign new_U6163 = ~new_U2422 | ~DATAI_7_;
  assign new_U6164 = ~new_U2386 | ~new_R2358_U21;
  assign new_U6165 = ~EAX_REG_7_ | ~new_U3411;
  assign new_U6166 = ~new_U2422 | ~DATAI_8_;
  assign new_U6167 = ~new_U2386 | ~new_R2358_U85;
  assign new_U6168 = ~EAX_REG_8_ | ~new_U3411;
  assign new_U6169 = ~new_U2422 | ~DATAI_9_;
  assign new_U6170 = ~new_U2386 | ~new_R2358_U83;
  assign new_U6171 = ~EAX_REG_9_ | ~new_U3411;
  assign new_U6172 = ~new_U2422 | ~DATAI_10_;
  assign new_U6173 = ~new_U2386 | ~new_R2358_U14;
  assign new_U6174 = ~EAX_REG_10_ | ~new_U3411;
  assign new_U6175 = ~new_U2422 | ~DATAI_11_;
  assign new_U6176 = ~new_U2386 | ~new_R2358_U15;
  assign new_U6177 = ~EAX_REG_11_ | ~new_U3411;
  assign new_U6178 = ~new_U2422 | ~DATAI_12_;
  assign new_U6179 = ~new_U2386 | ~new_R2358_U122;
  assign new_U6180 = ~EAX_REG_12_ | ~new_U3411;
  assign new_U6181 = ~new_U2422 | ~DATAI_13_;
  assign new_U6182 = ~new_U2386 | ~new_R2358_U120;
  assign new_U6183 = ~EAX_REG_13_ | ~new_U3411;
  assign new_U6184 = ~new_U2422 | ~DATAI_14_;
  assign new_U6185 = ~new_U2386 | ~new_R2358_U119;
  assign new_U6186 = ~EAX_REG_14_ | ~new_U3411;
  assign new_U6187 = ~new_U2422 | ~DATAI_15_;
  assign new_U6188 = ~new_U2386 | ~new_R2358_U16;
  assign new_U6189 = ~EAX_REG_15_ | ~new_U3411;
  assign new_U6190 = ~new_U2423 | ~DATAI_16_;
  assign new_U6191 = ~new_U2387 | ~DATAI_0_;
  assign new_U6192 = ~new_U2386 | ~new_R2358_U17;
  assign new_U6193 = ~EAX_REG_16_ | ~new_U3411;
  assign new_U6194 = ~new_U2423 | ~DATAI_17_;
  assign new_U6195 = ~new_U2387 | ~DATAI_1_;
  assign new_U6196 = ~new_U2386 | ~new_R2358_U118;
  assign new_U6197 = ~EAX_REG_17_ | ~new_U3411;
  assign new_U6198 = ~new_U2423 | ~DATAI_18_;
  assign new_U6199 = ~new_U2387 | ~DATAI_2_;
  assign new_U6200 = ~new_U2386 | ~new_R2358_U116;
  assign new_U6201 = ~EAX_REG_18_ | ~new_U3411;
  assign new_U6202 = ~new_U2423 | ~DATAI_19_;
  assign new_U6203 = ~new_U2387 | ~DATAI_3_;
  assign new_U6204 = ~new_U2386 | ~new_R2358_U114;
  assign new_U6205 = ~EAX_REG_19_ | ~new_U3411;
  assign new_U6206 = ~new_U2423 | ~DATAI_20_;
  assign new_U6207 = ~new_U2387 | ~DATAI_4_;
  assign new_U6208 = ~new_U2386 | ~new_R2358_U110;
  assign new_U6209 = ~EAX_REG_20_ | ~new_U3411;
  assign new_U6210 = ~new_U2423 | ~DATAI_21_;
  assign new_U6211 = ~new_U2387 | ~DATAI_5_;
  assign new_U6212 = ~new_U2386 | ~new_R2358_U18;
  assign new_U6213 = ~EAX_REG_21_ | ~new_U3411;
  assign new_U6214 = ~new_U2423 | ~DATAI_22_;
  assign new_U6215 = ~new_U2387 | ~DATAI_6_;
  assign new_U6216 = ~new_U2386 | ~new_R2358_U109;
  assign new_U6217 = ~EAX_REG_22_ | ~new_U3411;
  assign new_U6218 = ~new_U2423 | ~DATAI_23_;
  assign new_U6219 = ~new_U2387 | ~DATAI_7_;
  assign new_U6220 = ~new_U2386 | ~new_R2358_U107;
  assign new_U6221 = ~EAX_REG_23_ | ~new_U3411;
  assign new_U6222 = ~new_U2423 | ~DATAI_24_;
  assign new_U6223 = ~new_U2387 | ~DATAI_8_;
  assign new_U6224 = ~new_U2386 | ~new_R2358_U105;
  assign new_U6225 = ~EAX_REG_24_ | ~new_U3411;
  assign new_U6226 = ~new_U2423 | ~DATAI_25_;
  assign new_U6227 = ~new_U2387 | ~DATAI_9_;
  assign new_U6228 = ~new_U2386 | ~new_R2358_U103;
  assign new_U6229 = ~EAX_REG_25_ | ~new_U3411;
  assign new_U6230 = ~new_U2423 | ~DATAI_26_;
  assign new_U6231 = ~new_U2387 | ~DATAI_10_;
  assign new_U6232 = ~new_U2386 | ~new_R2358_U101;
  assign new_U6233 = ~EAX_REG_26_ | ~new_U3411;
  assign new_U6234 = ~new_U2423 | ~DATAI_27_;
  assign new_U6235 = ~new_U2387 | ~DATAI_11_;
  assign new_U6236 = ~new_U2386 | ~new_R2358_U99;
  assign new_U6237 = ~EAX_REG_27_ | ~new_U3411;
  assign new_U6238 = ~new_U2423 | ~DATAI_28_;
  assign new_U6239 = ~new_U2387 | ~DATAI_12_;
  assign new_U6240 = ~new_U2386 | ~new_R2358_U97;
  assign new_U6241 = ~EAX_REG_28_ | ~new_U3411;
  assign new_U6242 = ~new_U2423 | ~DATAI_29_;
  assign new_U6243 = ~new_U2387 | ~DATAI_13_;
  assign new_U6244 = ~new_U2386 | ~new_R2358_U95;
  assign new_U6245 = ~EAX_REG_29_ | ~new_U3411;
  assign new_U6246 = ~new_U2423 | ~DATAI_30_;
  assign new_U6247 = ~new_U2387 | ~DATAI_14_;
  assign new_U6248 = ~new_U2386 | ~new_R2358_U93;
  assign new_U6249 = ~EAX_REG_30_ | ~new_U3411;
  assign new_U6250 = ~new_U2423 | ~DATAI_31_;
  assign new_U6251 = ~new_U4186 | ~new_U3260;
  assign new_U6252 = ~new_U4193 | ~new_U6251;
  assign new_U6253 = ~new_U2383 | ~new_R2358_U82;
  assign new_U6254 = ~new_U2371 | ~new_R2099_U86;
  assign new_U6255 = ~EBX_REG_0_ | ~new_U3413;
  assign new_U6256 = ~new_U2383 | ~new_R2358_U112;
  assign new_U6257 = ~new_U2371 | ~new_R2099_U87;
  assign new_U6258 = ~EBX_REG_1_ | ~new_U3413;
  assign new_U6259 = ~new_U2383 | ~new_R2358_U19;
  assign new_U6260 = ~new_U2371 | ~new_R2099_U138;
  assign new_U6261 = ~EBX_REG_2_ | ~new_U3413;
  assign new_U6262 = ~new_U2383 | ~new_R2358_U20;
  assign new_U6263 = ~new_U2371 | ~new_R2099_U42;
  assign new_U6264 = ~EBX_REG_3_ | ~new_U3413;
  assign new_U6265 = ~new_U2383 | ~new_R2358_U90;
  assign new_U6266 = ~new_U2371 | ~new_R2099_U41;
  assign new_U6267 = ~EBX_REG_4_ | ~new_U3413;
  assign new_U6268 = ~new_U2383 | ~new_R2358_U88;
  assign new_U6269 = ~new_U2371 | ~new_R2099_U40;
  assign new_U6270 = ~EBX_REG_5_ | ~new_U3413;
  assign new_U6271 = ~new_U2383 | ~new_R2358_U86;
  assign new_U6272 = ~new_U2371 | ~new_R2099_U39;
  assign new_U6273 = ~EBX_REG_6_ | ~new_U3413;
  assign new_U6274 = ~new_U2383 | ~new_R2358_U21;
  assign new_U6275 = ~new_U2371 | ~new_R2099_U38;
  assign new_U6276 = ~EBX_REG_7_ | ~new_U3413;
  assign new_U6277 = ~new_U2383 | ~new_R2358_U85;
  assign new_U6278 = ~new_U2371 | ~new_R2099_U37;
  assign new_U6279 = ~EBX_REG_8_ | ~new_U3413;
  assign new_U6280 = ~new_U2383 | ~new_R2358_U83;
  assign new_U6281 = ~new_U2371 | ~new_R2099_U36;
  assign new_U6282 = ~EBX_REG_9_ | ~new_U3413;
  assign new_U6283 = ~new_U2383 | ~new_R2358_U14;
  assign new_U6284 = ~new_U2371 | ~new_R2099_U85;
  assign new_U6285 = ~EBX_REG_10_ | ~new_U3413;
  assign new_U6286 = ~new_U2383 | ~new_R2358_U15;
  assign new_U6287 = ~new_U2371 | ~new_R2099_U84;
  assign new_U6288 = ~EBX_REG_11_ | ~new_U3413;
  assign new_U6289 = ~new_U2383 | ~new_R2358_U122;
  assign new_U6290 = ~new_U2371 | ~new_R2099_U83;
  assign new_U6291 = ~EBX_REG_12_ | ~new_U3413;
  assign new_U6292 = ~new_U2383 | ~new_R2358_U120;
  assign new_U6293 = ~new_U2371 | ~new_R2099_U82;
  assign new_U6294 = ~EBX_REG_13_ | ~new_U3413;
  assign new_U6295 = ~new_U2383 | ~new_R2358_U119;
  assign new_U6296 = ~new_U2371 | ~new_R2099_U81;
  assign new_U6297 = ~EBX_REG_14_ | ~new_U3413;
  assign new_U6298 = ~new_U2383 | ~new_R2358_U16;
  assign new_U6299 = ~new_U2371 | ~new_R2099_U80;
  assign new_U6300 = ~EBX_REG_15_ | ~new_U3413;
  assign new_U6301 = ~new_U2383 | ~new_R2358_U17;
  assign new_U6302 = ~new_U2371 | ~new_R2099_U79;
  assign new_U6303 = ~EBX_REG_16_ | ~new_U3413;
  assign new_U6304 = ~new_U2383 | ~new_R2358_U118;
  assign new_U6305 = ~new_U2371 | ~new_R2099_U78;
  assign new_U6306 = ~EBX_REG_17_ | ~new_U3413;
  assign new_U6307 = ~new_U2383 | ~new_R2358_U116;
  assign new_U6308 = ~new_U2371 | ~new_R2099_U77;
  assign new_U6309 = ~EBX_REG_18_ | ~new_U3413;
  assign new_U6310 = ~new_U2383 | ~new_R2358_U114;
  assign new_U6311 = ~new_U2371 | ~new_R2099_U76;
  assign new_U6312 = ~EBX_REG_19_ | ~new_U3413;
  assign new_U6313 = ~new_U2383 | ~new_R2358_U110;
  assign new_U6314 = ~new_U2371 | ~new_R2099_U75;
  assign new_U6315 = ~EBX_REG_20_ | ~new_U3413;
  assign new_U6316 = ~new_U2383 | ~new_R2358_U18;
  assign new_U6317 = ~new_U2371 | ~new_R2099_U74;
  assign new_U6318 = ~EBX_REG_21_ | ~new_U3413;
  assign new_U6319 = ~new_U2383 | ~new_R2358_U109;
  assign new_U6320 = ~new_U2371 | ~new_R2099_U73;
  assign new_U6321 = ~EBX_REG_22_ | ~new_U3413;
  assign new_U6322 = ~new_U2383 | ~new_R2358_U107;
  assign new_U6323 = ~new_U2371 | ~new_R2099_U72;
  assign new_U6324 = ~EBX_REG_23_ | ~new_U3413;
  assign new_U6325 = ~new_U2383 | ~new_R2358_U105;
  assign new_U6326 = ~new_U2371 | ~new_R2099_U71;
  assign new_U6327 = ~EBX_REG_24_ | ~new_U3413;
  assign new_U6328 = ~new_U2383 | ~new_R2358_U103;
  assign new_U6329 = ~new_U2371 | ~new_R2099_U70;
  assign new_U6330 = ~EBX_REG_25_ | ~new_U3413;
  assign new_U6331 = ~new_U2383 | ~new_R2358_U101;
  assign new_U6332 = ~new_U2371 | ~new_R2099_U69;
  assign new_U6333 = ~EBX_REG_26_ | ~new_U3413;
  assign new_U6334 = ~new_U2383 | ~new_R2358_U99;
  assign new_U6335 = ~new_U2371 | ~new_R2099_U68;
  assign new_U6336 = ~EBX_REG_27_ | ~new_U3413;
  assign new_U6337 = ~new_U2383 | ~new_R2358_U97;
  assign new_U6338 = ~new_U2371 | ~new_R2099_U67;
  assign new_U6339 = ~EBX_REG_28_ | ~new_U3413;
  assign new_U6340 = ~new_U2383 | ~new_R2358_U95;
  assign new_U6341 = ~new_U2371 | ~new_R2099_U66;
  assign new_U6342 = ~EBX_REG_29_ | ~new_U3413;
  assign new_U6343 = ~new_U2383 | ~new_R2358_U93;
  assign new_U6344 = ~new_U2371 | ~new_R2099_U65;
  assign new_U6345 = ~EBX_REG_30_ | ~new_U3413;
  assign new_U6346 = ~new_U2371 | ~new_R2099_U64;
  assign new_U6347 = ~EBX_REG_31_ | ~new_U3413;
  assign new_U6348 = ~new_U4192 | ~new_GTE_485_U6;
  assign new_U6349 = ~new_U4190 | ~new_R2167_U17;
  assign new_U6350 = ~new_U4191 | ~new_U3250;
  assign new_U6351 = ~new_U3418;
  assign new_U6352 = ~new_U4237 | ~STATE2_REG_2_;
  assign new_U6353 = ~new_R2337_U58 | ~STATE2_REG_1_;
  assign new_U6354 = ~new_U6353 | ~new_U6352;
  assign new_U6355 = STATEBS16_REG | READY_N;
  assign new_U6356 = ~new_U2604 | ~new_R2099_U86;
  assign new_U6357 = ~REIP_REG_0_ | ~new_U7473;
  assign new_U6358 = ~EBX_REG_0_ | ~new_U7472;
  assign new_U6359 = ~new_U2429 | ~new_R2358_U82;
  assign new_U6360 = ~new_U2426 | ~new_R2182_U34;
  assign new_U6361 = ~new_U2373 | ~PHYADDRPOINTER_REG_0_;
  assign new_U6362 = ~new_U2366 | ~PHYADDRPOINTER_REG_0_;
  assign new_U6363 = ~new_U6351 | ~REIP_REG_0_;
  assign new_U6364 = ~new_U2604 | ~new_R2099_U87;
  assign new_U6365 = ~new_R2096_U4 | ~new_U7473;
  assign new_U6366 = ~EBX_REG_1_ | ~new_U7472;
  assign new_U6367 = ~new_U2429 | ~new_R2358_U112;
  assign new_U6368 = ~new_U2426 | ~new_R2182_U33;
  assign new_U6369 = ~new_U2373 | ~PHYADDRPOINTER_REG_1_;
  assign new_U6370 = ~new_U2366 | ~new_R2337_U5;
  assign new_U6371 = ~new_U6351 | ~REIP_REG_1_;
  assign new_U6372 = ~new_U2604 | ~new_R2099_U138;
  assign new_U6373 = ~new_R2096_U71 | ~new_U7473;
  assign new_U6374 = ~EBX_REG_2_ | ~new_U7472;
  assign new_U6375 = ~new_U2429 | ~new_R2358_U19;
  assign new_U6376 = ~new_U2426 | ~new_R2182_U42;
  assign new_U6377 = ~new_U2373 | ~PHYADDRPOINTER_REG_2_;
  assign new_U6378 = ~new_U2366 | ~new_R2337_U60;
  assign new_U6379 = ~new_U6351 | ~REIP_REG_2_;
  assign new_U6380 = ~new_U2604 | ~new_R2099_U42;
  assign new_U6381 = ~new_R2096_U68 | ~new_U7473;
  assign new_U6382 = ~EBX_REG_3_ | ~new_U7472;
  assign new_U6383 = ~new_U2429 | ~new_R2358_U20;
  assign new_U6384 = ~new_U2426 | ~new_R2182_U25;
  assign new_U6385 = ~new_U2373 | ~PHYADDRPOINTER_REG_3_;
  assign new_U6386 = ~new_U2366 | ~new_R2337_U57;
  assign new_U6387 = ~new_U6351 | ~REIP_REG_3_;
  assign new_U6388 = ~new_U2604 | ~new_R2099_U41;
  assign new_U6389 = ~new_R2096_U67 | ~new_U7473;
  assign new_U6390 = ~EBX_REG_4_ | ~new_U7472;
  assign new_U6391 = ~new_U2429 | ~new_R2358_U90;
  assign new_U6392 = ~new_U2426 | ~new_R2182_U24;
  assign new_U6393 = ~new_U2373 | ~PHYADDRPOINTER_REG_4_;
  assign new_U6394 = ~new_U2366 | ~new_R2337_U56;
  assign new_U6395 = ~new_U6351 | ~REIP_REG_4_;
  assign new_U6396 = ~new_U2604 | ~new_R2099_U40;
  assign new_U6397 = ~new_R2096_U66 | ~new_U7473;
  assign new_U6398 = ~EBX_REG_5_ | ~new_U7472;
  assign new_U6399 = ~new_U2429 | ~new_R2358_U88;
  assign new_U6400 = ~new_R2182_U5 | ~new_U2426;
  assign new_U6401 = ~new_U2373 | ~PHYADDRPOINTER_REG_5_;
  assign new_U6402 = ~new_U2366 | ~new_R2337_U55;
  assign new_U6403 = ~new_U6351 | ~REIP_REG_5_;
  assign new_U6404 = ~new_U2604 | ~new_R2099_U39;
  assign new_U6405 = ~new_R2096_U65 | ~new_U7473;
  assign new_U6406 = ~EBX_REG_6_ | ~new_U7472;
  assign new_U6407 = ~new_U2373 | ~PHYADDRPOINTER_REG_6_;
  assign new_U6408 = ~new_U2367 | ~new_R2358_U86;
  assign new_U6409 = ~new_U2366 | ~new_R2337_U54;
  assign new_U6410 = ~new_U6351 | ~REIP_REG_6_;
  assign new_U6411 = ~new_U2604 | ~new_R2099_U38;
  assign new_U6412 = ~new_R2096_U64 | ~new_U7473;
  assign new_U6413 = ~EBX_REG_7_ | ~new_U7472;
  assign new_U6414 = ~new_U2373 | ~PHYADDRPOINTER_REG_7_;
  assign new_U6415 = ~new_U2367 | ~new_R2358_U21;
  assign new_U6416 = ~new_U2366 | ~new_R2337_U53;
  assign new_U6417 = ~new_U6351 | ~REIP_REG_7_;
  assign new_U6418 = ~new_U2604 | ~new_R2099_U37;
  assign new_U6419 = ~new_R2096_U63 | ~new_U7473;
  assign new_U6420 = ~EBX_REG_8_ | ~new_U7472;
  assign new_U6421 = ~new_U2373 | ~PHYADDRPOINTER_REG_8_;
  assign new_U6422 = ~new_U2367 | ~new_R2358_U85;
  assign new_U6423 = ~new_U2366 | ~new_R2337_U52;
  assign new_U6424 = ~new_U6351 | ~REIP_REG_8_;
  assign new_U6425 = ~new_U2604 | ~new_R2099_U36;
  assign new_U6426 = ~new_R2096_U62 | ~new_U7473;
  assign new_U6427 = ~EBX_REG_9_ | ~new_U7472;
  assign new_U6428 = ~new_U2373 | ~PHYADDRPOINTER_REG_9_;
  assign new_U6429 = ~new_U2367 | ~new_R2358_U83;
  assign new_U6430 = ~new_U2366 | ~new_R2337_U51;
  assign new_U6431 = ~new_U6351 | ~REIP_REG_9_;
  assign new_U6432 = ~new_U2604 | ~new_R2099_U85;
  assign new_U6433 = ~new_R2096_U91 | ~new_U7473;
  assign new_U6434 = ~EBX_REG_10_ | ~new_U7472;
  assign new_U6435 = ~new_U2373 | ~PHYADDRPOINTER_REG_10_;
  assign new_U6436 = ~new_U2367 | ~new_R2358_U14;
  assign new_U6437 = ~new_U2366 | ~new_R2337_U80;
  assign new_U6438 = ~new_U6351 | ~REIP_REG_10_;
  assign new_U6439 = ~new_U2604 | ~new_R2099_U84;
  assign new_U6440 = ~new_R2096_U90 | ~new_U7473;
  assign new_U6441 = ~EBX_REG_11_ | ~new_U7472;
  assign new_U6442 = ~new_U2373 | ~PHYADDRPOINTER_REG_11_;
  assign new_U6443 = ~new_U2367 | ~new_R2358_U15;
  assign new_U6444 = ~new_U2366 | ~new_R2337_U79;
  assign new_U6445 = ~new_U6351 | ~REIP_REG_11_;
  assign new_U6446 = ~new_U2604 | ~new_R2099_U83;
  assign new_U6447 = ~new_R2096_U89 | ~new_U7473;
  assign new_U6448 = ~EBX_REG_12_ | ~new_U7472;
  assign new_U6449 = ~new_U2373 | ~PHYADDRPOINTER_REG_12_;
  assign new_U6450 = ~new_U2367 | ~new_R2358_U122;
  assign new_U6451 = ~new_U2366 | ~new_R2337_U78;
  assign new_U6452 = ~new_U6351 | ~REIP_REG_12_;
  assign new_U6453 = ~new_U2604 | ~new_R2099_U82;
  assign new_U6454 = ~new_R2096_U88 | ~new_U7473;
  assign new_U6455 = ~EBX_REG_13_ | ~new_U7472;
  assign new_U6456 = ~new_U2373 | ~PHYADDRPOINTER_REG_13_;
  assign new_U6457 = ~new_U2367 | ~new_R2358_U120;
  assign new_U6458 = ~new_U2366 | ~new_R2337_U77;
  assign new_U6459 = ~new_U6351 | ~REIP_REG_13_;
  assign new_U6460 = ~new_U2604 | ~new_R2099_U81;
  assign new_U6461 = ~new_R2096_U87 | ~new_U7473;
  assign new_U6462 = ~EBX_REG_14_ | ~new_U7472;
  assign new_U6463 = ~new_U2373 | ~PHYADDRPOINTER_REG_14_;
  assign new_U6464 = ~new_U2367 | ~new_R2358_U119;
  assign new_U6465 = ~new_U2366 | ~new_R2337_U76;
  assign new_U6466 = ~new_U6351 | ~REIP_REG_14_;
  assign new_U6467 = ~new_U2604 | ~new_R2099_U80;
  assign new_U6468 = ~new_R2096_U86 | ~new_U7473;
  assign new_U6469 = ~EBX_REG_15_ | ~new_U7472;
  assign new_U6470 = ~new_U2373 | ~PHYADDRPOINTER_REG_15_;
  assign new_U6471 = ~new_U2367 | ~new_R2358_U16;
  assign new_U6472 = ~new_U2366 | ~new_R2337_U75;
  assign new_U6473 = ~new_U6351 | ~REIP_REG_15_;
  assign new_U6474 = ~new_U2604 | ~new_R2099_U79;
  assign new_U6475 = ~new_R2096_U85 | ~new_U7473;
  assign new_U6476 = ~EBX_REG_16_ | ~new_U7472;
  assign new_U6477 = ~new_U2373 | ~PHYADDRPOINTER_REG_16_;
  assign new_U6478 = ~new_U2367 | ~new_R2358_U17;
  assign new_U6479 = ~new_U2366 | ~new_R2337_U74;
  assign new_U6480 = ~new_U6351 | ~REIP_REG_16_;
  assign new_U6481 = ~new_U2604 | ~new_R2099_U78;
  assign new_U6482 = ~new_R2096_U84 | ~new_U7473;
  assign new_U6483 = ~EBX_REG_17_ | ~new_U7472;
  assign new_U6484 = ~new_U2373 | ~PHYADDRPOINTER_REG_17_;
  assign new_U6485 = ~new_U2367 | ~new_R2358_U118;
  assign new_U6486 = ~new_U2366 | ~new_R2337_U73;
  assign new_U6487 = ~new_U6351 | ~REIP_REG_17_;
  assign new_U6488 = ~new_U2604 | ~new_R2099_U77;
  assign new_U6489 = ~new_R2096_U83 | ~new_U7473;
  assign new_U6490 = ~EBX_REG_18_ | ~new_U7472;
  assign new_U6491 = ~new_U2373 | ~PHYADDRPOINTER_REG_18_;
  assign new_U6492 = ~new_U2367 | ~new_R2358_U116;
  assign new_U6493 = ~new_U2366 | ~new_R2337_U72;
  assign new_U6494 = ~new_U6351 | ~REIP_REG_18_;
  assign new_U6495 = ~new_U2604 | ~new_R2099_U76;
  assign new_U6496 = ~new_R2096_U82 | ~new_U7473;
  assign new_U6497 = ~EBX_REG_19_ | ~new_U7472;
  assign new_U6498 = ~new_U2373 | ~PHYADDRPOINTER_REG_19_;
  assign new_U6499 = ~new_U2367 | ~new_R2358_U114;
  assign new_U6500 = ~new_U2366 | ~new_R2337_U71;
  assign new_U6501 = ~new_U6351 | ~REIP_REG_19_;
  assign new_U6502 = ~new_U2604 | ~new_R2099_U75;
  assign new_U6503 = ~new_R2096_U81 | ~new_U7473;
  assign new_U6504 = ~EBX_REG_20_ | ~new_U7472;
  assign new_U6505 = ~new_U2373 | ~PHYADDRPOINTER_REG_20_;
  assign new_U6506 = ~new_U2367 | ~new_R2358_U110;
  assign new_U6507 = ~new_U2366 | ~new_R2337_U70;
  assign new_U6508 = ~new_U6351 | ~REIP_REG_20_;
  assign new_U6509 = ~new_U2604 | ~new_R2099_U74;
  assign new_U6510 = ~new_R2096_U80 | ~new_U7473;
  assign new_U6511 = ~EBX_REG_21_ | ~new_U7472;
  assign new_U6512 = ~new_U2373 | ~PHYADDRPOINTER_REG_21_;
  assign new_U6513 = ~new_U2367 | ~new_R2358_U18;
  assign new_U6514 = ~new_U2366 | ~new_R2337_U69;
  assign new_U6515 = ~new_U6351 | ~REIP_REG_21_;
  assign new_U6516 = ~new_U2604 | ~new_R2099_U73;
  assign new_U6517 = ~new_R2096_U79 | ~new_U7473;
  assign new_U6518 = ~EBX_REG_22_ | ~new_U7472;
  assign new_U6519 = ~new_U2373 | ~PHYADDRPOINTER_REG_22_;
  assign new_U6520 = ~new_U2367 | ~new_R2358_U109;
  assign new_U6521 = ~new_U2366 | ~new_R2337_U68;
  assign new_U6522 = ~new_U6351 | ~REIP_REG_22_;
  assign new_U6523 = ~new_U2604 | ~new_R2099_U72;
  assign new_U6524 = ~new_R2096_U78 | ~new_U7473;
  assign new_U6525 = ~EBX_REG_23_ | ~new_U7472;
  assign new_U6526 = ~new_U2373 | ~PHYADDRPOINTER_REG_23_;
  assign new_U6527 = ~new_U2367 | ~new_R2358_U107;
  assign new_U6528 = ~new_U2366 | ~new_R2337_U67;
  assign new_U6529 = ~new_U6351 | ~REIP_REG_23_;
  assign new_U6530 = ~new_U2604 | ~new_R2099_U71;
  assign new_U6531 = ~new_R2096_U77 | ~new_U7473;
  assign new_U6532 = ~EBX_REG_24_ | ~new_U7472;
  assign new_U6533 = ~new_U2373 | ~PHYADDRPOINTER_REG_24_;
  assign new_U6534 = ~new_U2367 | ~new_R2358_U105;
  assign new_U6535 = ~new_U2366 | ~new_R2337_U66;
  assign new_U6536 = ~new_U6351 | ~REIP_REG_24_;
  assign new_U6537 = ~new_U2604 | ~new_R2099_U70;
  assign new_U6538 = ~new_R2096_U76 | ~new_U7473;
  assign new_U6539 = ~EBX_REG_25_ | ~new_U7472;
  assign new_U6540 = ~new_U2373 | ~PHYADDRPOINTER_REG_25_;
  assign new_U6541 = ~new_U2367 | ~new_R2358_U103;
  assign new_U6542 = ~new_U2366 | ~new_R2337_U65;
  assign new_U6543 = ~new_U6351 | ~REIP_REG_25_;
  assign new_U6544 = ~new_U2604 | ~new_R2099_U69;
  assign new_U6545 = ~new_R2096_U75 | ~new_U7473;
  assign new_U6546 = ~EBX_REG_26_ | ~new_U7472;
  assign new_U6547 = ~new_U2373 | ~PHYADDRPOINTER_REG_26_;
  assign new_U6548 = ~new_U2367 | ~new_R2358_U101;
  assign new_U6549 = ~new_U2366 | ~new_R2337_U64;
  assign new_U6550 = ~new_U6351 | ~REIP_REG_26_;
  assign new_U6551 = ~new_U2604 | ~new_R2099_U68;
  assign new_U6552 = ~new_R2096_U74 | ~new_U7473;
  assign new_U6553 = ~EBX_REG_27_ | ~new_U7472;
  assign new_U6554 = ~new_U2373 | ~PHYADDRPOINTER_REG_27_;
  assign new_U6555 = ~new_U2367 | ~new_R2358_U99;
  assign new_U6556 = ~new_U2366 | ~new_R2337_U63;
  assign new_U6557 = ~new_U6351 | ~REIP_REG_27_;
  assign new_U6558 = ~new_U2604 | ~new_R2099_U67;
  assign new_U6559 = ~new_R2096_U73 | ~new_U7473;
  assign new_U6560 = ~EBX_REG_28_ | ~new_U7472;
  assign new_U6561 = ~new_U2373 | ~PHYADDRPOINTER_REG_28_;
  assign new_U6562 = ~new_U2367 | ~new_R2358_U97;
  assign new_U6563 = ~new_U2366 | ~new_R2337_U62;
  assign new_U6564 = ~new_U6351 | ~REIP_REG_28_;
  assign new_U6565 = ~new_U2604 | ~new_R2099_U66;
  assign new_U6566 = ~new_R2096_U72 | ~new_U7473;
  assign new_U6567 = ~EBX_REG_29_ | ~new_U7472;
  assign new_U6568 = ~new_U2373 | ~PHYADDRPOINTER_REG_29_;
  assign new_U6569 = ~new_U2367 | ~new_R2358_U95;
  assign new_U6570 = ~new_U2366 | ~new_R2337_U61;
  assign new_U6571 = ~new_U6351 | ~REIP_REG_29_;
  assign new_U6572 = ~new_U2604 | ~new_R2099_U65;
  assign new_U6573 = ~new_R2096_U70 | ~new_U7473;
  assign new_U6574 = ~EBX_REG_30_ | ~new_U7472;
  assign new_U6575 = ~new_U2373 | ~PHYADDRPOINTER_REG_30_;
  assign new_U6576 = ~new_U2367 | ~new_R2358_U93;
  assign new_U6577 = ~new_U2366 | ~new_R2337_U59;
  assign new_U6578 = ~new_U6351 | ~REIP_REG_30_;
  assign new_U6579 = ~new_U2604 | ~new_R2099_U64;
  assign new_U6580 = ~new_R2096_U69 | ~new_U7473;
  assign new_U6581 = ~EBX_REG_31_ | ~new_U7472;
  assign new_U6582 = ~new_U2373 | ~PHYADDRPOINTER_REG_31_;
  assign new_U6583 = ~new_U2367 | ~new_R2358_U91;
  assign new_U6584 = ~new_U2366 | ~new_R2337_U58;
  assign new_U6585 = ~new_U6351 | ~REIP_REG_31_;
  assign new_U6586 = ~DATAWIDTH_REG_1_ | ~DATAWIDTH_REG_0_;
  assign new_U6587 = REIP_REG_1_ | REIP_REG_0_;
  assign new_U6588 = ~new_U4165;
  assign new_U6589 = ~FLUSH_REG | ~new_U4165;
  assign new_U6590 = ~new_U3954 | ~new_U2428;
  assign new_U6591 = ~new_U4168;
  assign new_U6592 = ~STATEBS16_REG | ~new_U4485;
  assign new_U6593 = ~new_U4196 | ~new_U6592;
  assign new_U6594 = ~new_U3952 | ~new_U6593;
  assign new_U6595 = ~STATE2_REG_0_ | ~new_U6594;
  assign new_U6596 = ~new_U4181 | ~new_U3259;
  assign new_U6597 = ~new_U3953 | ~new_U6595;
  assign new_U6598 = ~new_U2368 | ~new_U2473;
  assign new_U6599 = ~CODEFETCH_REG | ~new_U6598;
  assign new_U6600 = ~new_U4243 | ~STATE2_REG_0_;
  assign new_U6601 = ~ADS_N_REG | ~STATE_REG_0_;
  assign new_U6602 = ~new_U4169;
  assign new_U6603 = ~new_U3956 | ~new_U3278;
  assign new_U6604 = ~new_U3393 | ~new_U4487 | ~new_U3957;
  assign new_U6605 = ~MEMORYFETCH_REG | ~new_U6604;
  assign new_U6606 = ~new_U2544 | ~INSTQUEUE_REG_15__7_;
  assign new_U6607 = ~new_U2543 | ~INSTQUEUE_REG_14__7_;
  assign new_U6608 = ~new_U2542 | ~INSTQUEUE_REG_13__7_;
  assign new_U6609 = ~new_U2541 | ~INSTQUEUE_REG_12__7_;
  assign new_U6610 = ~new_U2539 | ~INSTQUEUE_REG_11__7_;
  assign new_U6611 = ~new_U2538 | ~INSTQUEUE_REG_10__7_;
  assign new_U6612 = ~new_U2537 | ~INSTQUEUE_REG_9__7_;
  assign new_U6613 = ~new_U2536 | ~INSTQUEUE_REG_8__7_;
  assign new_U6614 = ~new_U2534 | ~INSTQUEUE_REG_7__7_;
  assign new_U6615 = ~new_U2533 | ~INSTQUEUE_REG_6__7_;
  assign new_U6616 = ~new_U2532 | ~INSTQUEUE_REG_5__7_;
  assign new_U6617 = ~new_U2531 | ~INSTQUEUE_REG_4__7_;
  assign new_U6618 = ~new_U2529 | ~INSTQUEUE_REG_3__7_;
  assign new_U6619 = ~new_U2527 | ~INSTQUEUE_REG_2__7_;
  assign new_U6620 = ~new_U2525 | ~INSTQUEUE_REG_1__7_;
  assign new_U6621 = ~new_U2523 | ~INSTQUEUE_REG_0__7_;
  assign new_U6622 = ~new_U2544 | ~INSTQUEUE_REG_15__6_;
  assign new_U6623 = ~new_U2543 | ~INSTQUEUE_REG_14__6_;
  assign new_U6624 = ~new_U2542 | ~INSTQUEUE_REG_13__6_;
  assign new_U6625 = ~new_U2541 | ~INSTQUEUE_REG_12__6_;
  assign new_U6626 = ~new_U2539 | ~INSTQUEUE_REG_11__6_;
  assign new_U6627 = ~new_U2538 | ~INSTQUEUE_REG_10__6_;
  assign new_U6628 = ~new_U2537 | ~INSTQUEUE_REG_9__6_;
  assign new_U6629 = ~new_U2536 | ~INSTQUEUE_REG_8__6_;
  assign new_U6630 = ~new_U2534 | ~INSTQUEUE_REG_7__6_;
  assign new_U6631 = ~new_U2533 | ~INSTQUEUE_REG_6__6_;
  assign new_U6632 = ~new_U2532 | ~INSTQUEUE_REG_5__6_;
  assign new_U6633 = ~new_U2531 | ~INSTQUEUE_REG_4__6_;
  assign new_U6634 = ~new_U2529 | ~INSTQUEUE_REG_3__6_;
  assign new_U6635 = ~new_U2527 | ~INSTQUEUE_REG_2__6_;
  assign new_U6636 = ~new_U2525 | ~INSTQUEUE_REG_1__6_;
  assign new_U6637 = ~new_U2523 | ~INSTQUEUE_REG_0__6_;
  assign new_U6638 = ~new_U2544 | ~INSTQUEUE_REG_15__5_;
  assign new_U6639 = ~new_U2543 | ~INSTQUEUE_REG_14__5_;
  assign new_U6640 = ~new_U2542 | ~INSTQUEUE_REG_13__5_;
  assign new_U6641 = ~new_U2541 | ~INSTQUEUE_REG_12__5_;
  assign new_U6642 = ~new_U2539 | ~INSTQUEUE_REG_11__5_;
  assign new_U6643 = ~new_U2538 | ~INSTQUEUE_REG_10__5_;
  assign new_U6644 = ~new_U2537 | ~INSTQUEUE_REG_9__5_;
  assign new_U6645 = ~new_U2536 | ~INSTQUEUE_REG_8__5_;
  assign new_U6646 = ~new_U2534 | ~INSTQUEUE_REG_7__5_;
  assign new_U6647 = ~new_U2533 | ~INSTQUEUE_REG_6__5_;
  assign new_U6648 = ~new_U2532 | ~INSTQUEUE_REG_5__5_;
  assign new_U6649 = ~new_U2531 | ~INSTQUEUE_REG_4__5_;
  assign new_U6650 = ~new_U2529 | ~INSTQUEUE_REG_3__5_;
  assign new_U6651 = ~new_U2527 | ~INSTQUEUE_REG_2__5_;
  assign new_U6652 = ~new_U2525 | ~INSTQUEUE_REG_1__5_;
  assign new_U6653 = ~new_U2523 | ~INSTQUEUE_REG_0__5_;
  assign new_U6654 = ~new_U2544 | ~INSTQUEUE_REG_15__4_;
  assign new_U6655 = ~new_U2543 | ~INSTQUEUE_REG_14__4_;
  assign new_U6656 = ~new_U2542 | ~INSTQUEUE_REG_13__4_;
  assign new_U6657 = ~new_U2541 | ~INSTQUEUE_REG_12__4_;
  assign new_U6658 = ~new_U2539 | ~INSTQUEUE_REG_11__4_;
  assign new_U6659 = ~new_U2538 | ~INSTQUEUE_REG_10__4_;
  assign new_U6660 = ~new_U2537 | ~INSTQUEUE_REG_9__4_;
  assign new_U6661 = ~new_U2536 | ~INSTQUEUE_REG_8__4_;
  assign new_U6662 = ~new_U2534 | ~INSTQUEUE_REG_7__4_;
  assign new_U6663 = ~new_U2533 | ~INSTQUEUE_REG_6__4_;
  assign new_U6664 = ~new_U2532 | ~INSTQUEUE_REG_5__4_;
  assign new_U6665 = ~new_U2531 | ~INSTQUEUE_REG_4__4_;
  assign new_U6666 = ~new_U2529 | ~INSTQUEUE_REG_3__4_;
  assign new_U6667 = ~new_U2527 | ~INSTQUEUE_REG_2__4_;
  assign new_U6668 = ~new_U2525 | ~INSTQUEUE_REG_1__4_;
  assign new_U6669 = ~new_U2544 | ~INSTQUEUE_REG_15__3_;
  assign new_U6670 = ~new_U2543 | ~INSTQUEUE_REG_14__3_;
  assign new_U6671 = ~new_U2542 | ~INSTQUEUE_REG_13__3_;
  assign new_U6672 = ~new_U2541 | ~INSTQUEUE_REG_12__3_;
  assign new_U6673 = ~new_U2539 | ~INSTQUEUE_REG_11__3_;
  assign new_U6674 = ~new_U2538 | ~INSTQUEUE_REG_10__3_;
  assign new_U6675 = ~new_U2537 | ~INSTQUEUE_REG_9__3_;
  assign new_U6676 = ~new_U2536 | ~INSTQUEUE_REG_8__3_;
  assign new_U6677 = ~new_U2534 | ~INSTQUEUE_REG_7__3_;
  assign new_U6678 = ~new_U2533 | ~INSTQUEUE_REG_6__3_;
  assign new_U6679 = ~new_U2532 | ~INSTQUEUE_REG_5__3_;
  assign new_U6680 = ~new_U2531 | ~INSTQUEUE_REG_4__3_;
  assign new_U6681 = ~new_U2529 | ~INSTQUEUE_REG_3__3_;
  assign new_U6682 = ~new_U2527 | ~INSTQUEUE_REG_2__3_;
  assign new_U6683 = ~new_U2525 | ~INSTQUEUE_REG_1__3_;
  assign new_U6684 = ~new_U2523 | ~INSTQUEUE_REG_0__3_;
  assign new_U6685 = ~new_U2544 | ~INSTQUEUE_REG_15__2_;
  assign new_U6686 = ~new_U2543 | ~INSTQUEUE_REG_14__2_;
  assign new_U6687 = ~new_U2542 | ~INSTQUEUE_REG_13__2_;
  assign new_U6688 = ~new_U2541 | ~INSTQUEUE_REG_12__2_;
  assign new_U6689 = ~new_U2539 | ~INSTQUEUE_REG_11__2_;
  assign new_U6690 = ~new_U2538 | ~INSTQUEUE_REG_10__2_;
  assign new_U6691 = ~new_U2537 | ~INSTQUEUE_REG_9__2_;
  assign new_U6692 = ~new_U2536 | ~INSTQUEUE_REG_8__2_;
  assign new_U6693 = ~new_U2534 | ~INSTQUEUE_REG_7__2_;
  assign new_U6694 = ~new_U2533 | ~INSTQUEUE_REG_6__2_;
  assign new_U6695 = ~new_U2532 | ~INSTQUEUE_REG_5__2_;
  assign new_U6696 = ~new_U2531 | ~INSTQUEUE_REG_4__2_;
  assign new_U6697 = ~new_U2529 | ~INSTQUEUE_REG_3__2_;
  assign new_U6698 = ~new_U2527 | ~INSTQUEUE_REG_2__2_;
  assign new_U6699 = ~new_U2525 | ~INSTQUEUE_REG_1__2_;
  assign new_U6700 = ~new_U2523 | ~INSTQUEUE_REG_0__2_;
  assign new_U6701 = ~new_U2544 | ~INSTQUEUE_REG_15__1_;
  assign new_U6702 = ~new_U2543 | ~INSTQUEUE_REG_14__1_;
  assign new_U6703 = ~new_U2542 | ~INSTQUEUE_REG_13__1_;
  assign new_U6704 = ~new_U2541 | ~INSTQUEUE_REG_12__1_;
  assign new_U6705 = ~new_U2539 | ~INSTQUEUE_REG_11__1_;
  assign new_U6706 = ~new_U2538 | ~INSTQUEUE_REG_10__1_;
  assign new_U6707 = ~new_U2537 | ~INSTQUEUE_REG_9__1_;
  assign new_U6708 = ~new_U2536 | ~INSTQUEUE_REG_8__1_;
  assign new_U6709 = ~new_U2534 | ~INSTQUEUE_REG_7__1_;
  assign new_U6710 = ~new_U2533 | ~INSTQUEUE_REG_6__1_;
  assign new_U6711 = ~new_U2532 | ~INSTQUEUE_REG_5__1_;
  assign new_U6712 = ~new_U2531 | ~INSTQUEUE_REG_4__1_;
  assign new_U6713 = ~new_U2529 | ~INSTQUEUE_REG_3__1_;
  assign new_U6714 = ~new_U2527 | ~INSTQUEUE_REG_2__1_;
  assign new_U6715 = ~new_U2525 | ~INSTQUEUE_REG_1__1_;
  assign new_U6716 = ~new_U2523 | ~INSTQUEUE_REG_0__1_;
  assign new_U6717 = ~new_U2544 | ~INSTQUEUE_REG_15__0_;
  assign new_U6718 = ~new_U2543 | ~INSTQUEUE_REG_14__0_;
  assign new_U6719 = ~new_U2542 | ~INSTQUEUE_REG_13__0_;
  assign new_U6720 = ~new_U2541 | ~INSTQUEUE_REG_12__0_;
  assign new_U6721 = ~new_U2539 | ~INSTQUEUE_REG_11__0_;
  assign new_U6722 = ~new_U2538 | ~INSTQUEUE_REG_10__0_;
  assign new_U6723 = ~new_U2537 | ~INSTQUEUE_REG_9__0_;
  assign new_U6724 = ~new_U2536 | ~INSTQUEUE_REG_8__0_;
  assign new_U6725 = ~new_U2534 | ~INSTQUEUE_REG_7__0_;
  assign new_U6726 = ~new_U2533 | ~INSTQUEUE_REG_6__0_;
  assign new_U6727 = ~new_U2532 | ~INSTQUEUE_REG_5__0_;
  assign new_U6728 = ~new_U2531 | ~INSTQUEUE_REG_4__0_;
  assign new_U6729 = ~new_U2529 | ~INSTQUEUE_REG_3__0_;
  assign new_U6730 = ~new_U2527 | ~INSTQUEUE_REG_2__0_;
  assign new_U6731 = ~new_U2525 | ~INSTQUEUE_REG_1__0_;
  assign new_U6732 = ~new_U2523 | ~INSTQUEUE_REG_0__0_;
  assign new_U6733 = ~new_U4448 | ~STATE2_REG_2_;
  assign new_U6734 = ~new_U3399 | ~new_U6733;
  assign new_U6735 = ~new_U4176 | ~EAX_REG_9_;
  assign new_U6736 = ~new_U4175 | ~PHYADDRPOINTER_REG_9_;
  assign new_U6737 = ~new_R2337_U51 | ~new_U2352;
  assign new_U6738 = ~new_U4176 | ~EAX_REG_8_;
  assign new_U6739 = ~new_U4175 | ~PHYADDRPOINTER_REG_8_;
  assign new_U6740 = ~new_R2337_U52 | ~new_U2352;
  assign new_U6741 = ~new_U4176 | ~EAX_REG_7_;
  assign new_U6742 = ~new_U4175 | ~PHYADDRPOINTER_REG_7_;
  assign new_U6743 = ~new_R2337_U53 | ~new_U2352;
  assign new_U6744 = ~new_U4176 | ~EAX_REG_6_;
  assign new_U6745 = ~new_U4175 | ~PHYADDRPOINTER_REG_6_;
  assign new_U6746 = ~new_R2337_U54 | ~new_U2352;
  assign new_U6747 = ~new_R2182_U5 | ~new_U6734;
  assign new_U6748 = ~new_U4176 | ~EAX_REG_5_;
  assign new_U6749 = ~new_U4175 | ~PHYADDRPOINTER_REG_5_;
  assign new_U6750 = ~new_R2337_U55 | ~new_U2352;
  assign new_U6751 = ~new_R2182_U24 | ~new_U6734;
  assign new_U6752 = ~new_U4176 | ~EAX_REG_4_;
  assign new_U6753 = ~new_U4175 | ~PHYADDRPOINTER_REG_4_;
  assign new_U6754 = ~new_R2337_U56 | ~new_U2352;
  assign new_U6755 = ~new_U2353 | ~INSTQUEUERD_ADDR_REG_4_;
  assign new_U6756 = ~new_U4176 | ~EAX_REG_31_;
  assign new_U6757 = ~new_U4175 | ~PHYADDRPOINTER_REG_31_;
  assign new_U6758 = ~new_R2337_U58 | ~new_U2352;
  assign new_U6759 = ~new_R2182_U26 | ~new_U6734;
  assign new_U6760 = ~new_U4176 | ~EAX_REG_30_;
  assign new_U6761 = ~new_U4175 | ~PHYADDRPOINTER_REG_30_;
  assign new_U6762 = ~new_R2337_U59 | ~new_U2352;
  assign new_U6763 = ~new_R2182_U25 | ~new_U6734;
  assign new_U6764 = ~new_U4176 | ~EAX_REG_3_;
  assign new_U6765 = ~new_U4175 | ~PHYADDRPOINTER_REG_3_;
  assign new_U6766 = ~new_R2337_U57 | ~new_U2352;
  assign new_U6767 = ~new_U2353 | ~INSTQUEUERD_ADDR_REG_3_;
  assign new_U6768 = ~new_R2182_U27 | ~new_U6734;
  assign new_U6769 = ~new_U4176 | ~EAX_REG_29_;
  assign new_U6770 = ~new_U4175 | ~PHYADDRPOINTER_REG_29_;
  assign new_U6771 = ~new_R2337_U61 | ~new_U2352;
  assign new_U6772 = ~new_R2182_U28 | ~new_U6734;
  assign new_U6773 = ~new_U4176 | ~EAX_REG_28_;
  assign new_U6774 = ~new_U4175 | ~PHYADDRPOINTER_REG_28_;
  assign new_U6775 = ~new_R2337_U62 | ~new_U2352;
  assign new_U6776 = ~new_R2182_U29 | ~new_U6734;
  assign new_U6777 = ~new_U4176 | ~EAX_REG_27_;
  assign new_U6778 = ~new_U4175 | ~PHYADDRPOINTER_REG_27_;
  assign new_U6779 = ~new_R2337_U63 | ~new_U2352;
  assign new_U6780 = ~new_R2182_U30 | ~new_U6734;
  assign new_U6781 = ~new_U4176 | ~EAX_REG_26_;
  assign new_U6782 = ~new_U4175 | ~PHYADDRPOINTER_REG_26_;
  assign new_U6783 = ~new_R2337_U64 | ~new_U2352;
  assign new_U6784 = ~new_R2182_U31 | ~new_U6734;
  assign new_U6785 = ~new_U4176 | ~EAX_REG_25_;
  assign new_U6786 = ~new_U4175 | ~PHYADDRPOINTER_REG_25_;
  assign new_U6787 = ~new_R2337_U65 | ~new_U2352;
  assign new_U6788 = ~new_R2182_U32 | ~new_U6734;
  assign new_U6789 = ~new_U4176 | ~EAX_REG_24_;
  assign new_U6790 = ~new_U4175 | ~PHYADDRPOINTER_REG_24_;
  assign new_U6791 = ~new_R2337_U66 | ~new_U2352;
  assign new_U6792 = ~new_R2182_U6 | ~new_U6734;
  assign new_U6793 = ~new_U4176 | ~EAX_REG_23_;
  assign new_U6794 = ~new_U4175 | ~PHYADDRPOINTER_REG_23_;
  assign new_U6795 = ~new_R2337_U67 | ~new_U2352;
  assign new_U6796 = ~new_U2724 | ~new_U6734;
  assign new_U6797 = ~new_U4176 | ~EAX_REG_22_;
  assign new_U6798 = ~new_U4175 | ~PHYADDRPOINTER_REG_22_;
  assign new_U6799 = ~new_R2337_U68 | ~new_U2352;
  assign new_U6800 = ~new_U2725 | ~new_U6734;
  assign new_U6801 = ~new_U4176 | ~EAX_REG_21_;
  assign new_U6802 = ~new_U4175 | ~PHYADDRPOINTER_REG_21_;
  assign new_U6803 = ~new_R2337_U69 | ~new_U2352;
  assign new_U6804 = ~new_U2726 | ~new_U6734;
  assign new_U6805 = ~new_U4176 | ~EAX_REG_20_;
  assign new_U6806 = ~new_U4175 | ~PHYADDRPOINTER_REG_20_;
  assign new_U6807 = ~new_R2337_U70 | ~new_U2352;
  assign new_U6808 = ~new_R2182_U42 | ~new_U6734;
  assign new_U6809 = ~new_U4176 | ~EAX_REG_2_;
  assign new_U6810 = ~new_U4175 | ~PHYADDRPOINTER_REG_2_;
  assign new_U6811 = ~new_R2337_U60 | ~new_U2352;
  assign new_U6812 = ~new_U2353 | ~INSTQUEUERD_ADDR_REG_2_;
  assign new_U6813 = ~new_U2727 | ~new_U6734;
  assign new_U6814 = ~new_U4176 | ~EAX_REG_19_;
  assign new_U6815 = ~new_U4175 | ~PHYADDRPOINTER_REG_19_;
  assign new_U6816 = ~new_R2337_U71 | ~new_U2352;
  assign new_U6817 = ~new_U2728 | ~new_U6734;
  assign new_U6818 = ~new_U4176 | ~EAX_REG_18_;
  assign new_U6819 = ~new_U4175 | ~PHYADDRPOINTER_REG_18_;
  assign new_U6820 = ~new_R2337_U72 | ~new_U2352;
  assign new_U6821 = ~new_U2729 | ~new_U6734;
  assign new_U6822 = ~new_U4176 | ~EAX_REG_17_;
  assign new_U6823 = ~new_U4175 | ~PHYADDRPOINTER_REG_17_;
  assign new_U6824 = ~new_R2337_U73 | ~new_U2352;
  assign new_U6825 = ~new_U2730 | ~new_U6734;
  assign new_U6826 = ~new_U4176 | ~EAX_REG_16_;
  assign new_U6827 = ~new_U4175 | ~PHYADDRPOINTER_REG_16_;
  assign new_U6828 = ~new_R2337_U74 | ~new_U2352;
  assign new_U6829 = ~new_U4176 | ~EAX_REG_15_;
  assign new_U6830 = ~new_U4175 | ~PHYADDRPOINTER_REG_15_;
  assign new_U6831 = ~new_R2337_U75 | ~new_U2352;
  assign new_U6832 = ~new_U4176 | ~EAX_REG_14_;
  assign new_U6833 = ~new_U4175 | ~PHYADDRPOINTER_REG_14_;
  assign new_U6834 = ~new_R2337_U76 | ~new_U2352;
  assign new_U6835 = ~new_U4176 | ~EAX_REG_13_;
  assign new_U6836 = ~new_U4175 | ~PHYADDRPOINTER_REG_13_;
  assign new_U6837 = ~new_R2337_U77 | ~new_U2352;
  assign new_U6838 = ~new_U4176 | ~EAX_REG_12_;
  assign new_U6839 = ~new_U4175 | ~PHYADDRPOINTER_REG_12_;
  assign new_U6840 = ~new_R2337_U78 | ~new_U2352;
  assign new_U6841 = ~new_U4176 | ~EAX_REG_11_;
  assign new_U6842 = ~new_U4175 | ~PHYADDRPOINTER_REG_11_;
  assign new_U6843 = ~new_R2337_U79 | ~new_U2352;
  assign new_U6844 = ~new_U4176 | ~EAX_REG_10_;
  assign new_U6845 = ~new_U4175 | ~PHYADDRPOINTER_REG_10_;
  assign new_U6846 = ~new_R2337_U80 | ~new_U2352;
  assign new_U6847 = ~new_R2182_U33 | ~new_U6734;
  assign new_U6848 = ~new_U4176 | ~EAX_REG_1_;
  assign new_U6849 = ~new_U4175 | ~PHYADDRPOINTER_REG_1_;
  assign new_U6850 = ~new_R2337_U5 | ~new_U2352;
  assign new_U6851 = ~new_U2353 | ~INSTQUEUERD_ADDR_REG_1_;
  assign new_U6852 = ~new_R2182_U34 | ~new_U6734;
  assign new_U6853 = ~new_U4176 | ~EAX_REG_0_;
  assign new_U6854 = ~new_U4175 | ~PHYADDRPOINTER_REG_0_;
  assign new_U6855 = ~PHYADDRPOINTER_REG_0_ | ~new_U2352;
  assign new_U6856 = ~new_U2353 | ~INSTQUEUERD_ADDR_REG_0_;
  assign new_U6857 = ~new_R2144_U49 | ~new_U6734;
  assign new_U6858 = ~new_U3296 | ~new_U3426 | ~new_U4448;
  assign new_U6859 = ~new_U4147 | ~new_R2144_U80;
  assign new_U6860 = ~new_ADD_371_U6 | ~new_U4196;
  assign new_U6861 = ~new_U4147 | ~new_R2144_U10;
  assign new_U6862 = ~new_ADD_371_U17 | ~new_U4196;
  assign new_U6863 = ~new_U4147 | ~new_R2144_U9;
  assign new_U6864 = ~new_ADD_371_U18 | ~new_U4196;
  assign new_U6865 = ~new_U4147 | ~new_R2144_U45;
  assign new_U6866 = ~new_ADD_371_U19 | ~new_U4196;
  assign new_U6867 = ~new_U4147 | ~new_R2144_U47;
  assign new_U6868 = ~new_ADD_371_U20 | ~new_U4196;
  assign new_U6869 = ~new_U4147 | ~new_R2144_U8;
  assign new_U6870 = ~new_ADD_371_U25 | ~new_U4196;
  assign new_U6871 = ~new_U4147 | ~new_R2144_U49;
  assign new_U6872 = ~new_ADD_371_U5 | ~new_U4196;
  assign new_U6873 = ~new_U4482 | ~new_U3270;
  assign new_U6874 = ~new_U4147 | ~new_R2144_U50;
  assign new_U6875 = ~new_ADD_371_U21 | ~new_U4196;
  assign new_U6876 = ~new_U2605 | ~new_U3271;
  assign new_U6877 = ~new_U4147 | ~new_R2144_U43;
  assign new_U6878 = ~new_ADD_371_U4 | ~new_U4196;
  assign new_U6879 = ~new_U4482 | ~new_U3270;
  assign new_U6880 = ~new_U2564 | ~INSTQUEUE_REG_15__1_;
  assign new_U6881 = ~new_U2563 | ~INSTQUEUE_REG_14__1_;
  assign new_U6882 = ~new_U2562 | ~INSTQUEUE_REG_13__1_;
  assign new_U6883 = ~new_U2561 | ~INSTQUEUE_REG_12__1_;
  assign new_U6884 = ~new_U2559 | ~INSTQUEUE_REG_11__1_;
  assign new_U6885 = ~new_U2558 | ~INSTQUEUE_REG_10__1_;
  assign new_U6886 = ~new_U2557 | ~INSTQUEUE_REG_9__1_;
  assign new_U6887 = ~new_U2556 | ~INSTQUEUE_REG_8__1_;
  assign new_U6888 = ~new_U2554 | ~INSTQUEUE_REG_7__1_;
  assign new_U6889 = ~new_U2553 | ~INSTQUEUE_REG_6__1_;
  assign new_U6890 = ~new_U2552 | ~INSTQUEUE_REG_5__1_;
  assign new_U6891 = ~new_U2551 | ~INSTQUEUE_REG_4__1_;
  assign new_U6892 = ~new_U2549 | ~INSTQUEUE_REG_3__1_;
  assign new_U6893 = ~new_U2548 | ~INSTQUEUE_REG_2__1_;
  assign new_U6894 = ~new_U2547 | ~INSTQUEUE_REG_1__1_;
  assign new_U6895 = ~new_U2546 | ~INSTQUEUE_REG_0__1_;
  assign new_U6896 = ~new_U4017 | ~new_U4018 | ~new_U4020 | ~new_U4019;
  assign new_U6897 = ~new_U3392 | ~new_U3405;
  assign new_U6898 = ~new_U2564 | ~INSTQUEUE_REG_15__0_;
  assign new_U6899 = ~new_U2563 | ~INSTQUEUE_REG_14__0_;
  assign new_U6900 = ~new_U2562 | ~INSTQUEUE_REG_13__0_;
  assign new_U6901 = ~new_U2561 | ~INSTQUEUE_REG_12__0_;
  assign new_U6902 = ~new_U2559 | ~INSTQUEUE_REG_11__0_;
  assign new_U6903 = ~new_U2558 | ~INSTQUEUE_REG_10__0_;
  assign new_U6904 = ~new_U2557 | ~INSTQUEUE_REG_9__0_;
  assign new_U6905 = ~new_U2556 | ~INSTQUEUE_REG_8__0_;
  assign new_U6906 = ~new_U2554 | ~INSTQUEUE_REG_7__0_;
  assign new_U6907 = ~new_U2553 | ~INSTQUEUE_REG_6__0_;
  assign new_U6908 = ~new_U2552 | ~INSTQUEUE_REG_5__0_;
  assign new_U6909 = ~new_U2551 | ~INSTQUEUE_REG_4__0_;
  assign new_U6910 = ~new_U2549 | ~INSTQUEUE_REG_3__0_;
  assign new_U6911 = ~new_U2548 | ~INSTQUEUE_REG_2__0_;
  assign new_U6912 = ~new_U2547 | ~INSTQUEUE_REG_1__0_;
  assign new_U6913 = ~new_U2546 | ~INSTQUEUE_REG_0__0_;
  assign new_U6914 = ~new_U4021 | ~new_U4022 | ~new_U4024 | ~new_U4023;
  assign new_U6915 = ~new_U4195 | ~new_U3221;
  assign new_U6916 = ~new_U2355 | ~new_SUB_357_U8;
  assign new_U6917 = ~new_U4195 | ~new_U3220;
  assign new_U6918 = ~new_SUB_357_U6 | ~new_U2355;
  assign new_U6919 = ~new_U4195 | ~new_U3219;
  assign new_U6920 = ~new_SUB_357_U9 | ~new_U2355;
  assign new_U6921 = ~new_U4195 | ~new_U3218;
  assign new_U6922 = ~new_SUB_357_U13 | ~new_U2355;
  assign new_U6923 = ~new_U4195 | ~new_U3217;
  assign new_U6924 = ~new_SUB_357_U11 | ~new_U2355;
  assign new_U6925 = ~new_R2182_U25 | ~new_U3281;
  assign new_U6926 = ~new_U4195 | ~new_U3216;
  assign new_U6927 = ~new_SUB_357_U12 | ~new_U2355;
  assign new_U6928 = ~new_R2182_U42 | ~new_U3281;
  assign new_U6929 = ~new_U2564 | ~INSTQUEUE_REG_15__7_;
  assign new_U6930 = ~new_U2563 | ~INSTQUEUE_REG_14__7_;
  assign new_U6931 = ~new_U2562 | ~INSTQUEUE_REG_13__7_;
  assign new_U6932 = ~new_U2561 | ~INSTQUEUE_REG_12__7_;
  assign new_U6933 = ~new_U2559 | ~INSTQUEUE_REG_11__7_;
  assign new_U6934 = ~new_U2558 | ~INSTQUEUE_REG_10__7_;
  assign new_U6935 = ~new_U2557 | ~INSTQUEUE_REG_9__7_;
  assign new_U6936 = ~new_U2556 | ~INSTQUEUE_REG_8__7_;
  assign new_U6937 = ~new_U2554 | ~INSTQUEUE_REG_7__7_;
  assign new_U6938 = ~new_U2553 | ~INSTQUEUE_REG_6__7_;
  assign new_U6939 = ~new_U2552 | ~INSTQUEUE_REG_5__7_;
  assign new_U6940 = ~new_U2551 | ~INSTQUEUE_REG_4__7_;
  assign new_U6941 = ~new_U2549 | ~INSTQUEUE_REG_3__7_;
  assign new_U6942 = ~new_U2548 | ~INSTQUEUE_REG_2__7_;
  assign new_U6943 = ~new_U2547 | ~INSTQUEUE_REG_1__7_;
  assign new_U6944 = ~new_U2546 | ~INSTQUEUE_REG_0__7_;
  assign new_U6945 = ~new_U4025 | ~new_U4026 | ~new_U4028 | ~new_U4027;
  assign new_U6946 = ~new_U2564 | ~INSTQUEUE_REG_15__6_;
  assign new_U6947 = ~new_U2563 | ~INSTQUEUE_REG_14__6_;
  assign new_U6948 = ~new_U2562 | ~INSTQUEUE_REG_13__6_;
  assign new_U6949 = ~new_U2561 | ~INSTQUEUE_REG_12__6_;
  assign new_U6950 = ~new_U2559 | ~INSTQUEUE_REG_11__6_;
  assign new_U6951 = ~new_U2558 | ~INSTQUEUE_REG_10__6_;
  assign new_U6952 = ~new_U2557 | ~INSTQUEUE_REG_9__6_;
  assign new_U6953 = ~new_U2556 | ~INSTQUEUE_REG_8__6_;
  assign new_U6954 = ~new_U2554 | ~INSTQUEUE_REG_7__6_;
  assign new_U6955 = ~new_U2553 | ~INSTQUEUE_REG_6__6_;
  assign new_U6956 = ~new_U2552 | ~INSTQUEUE_REG_5__6_;
  assign new_U6957 = ~new_U2551 | ~INSTQUEUE_REG_4__6_;
  assign new_U6958 = ~new_U2549 | ~INSTQUEUE_REG_3__6_;
  assign new_U6959 = ~new_U2548 | ~INSTQUEUE_REG_2__6_;
  assign new_U6960 = ~new_U2547 | ~INSTQUEUE_REG_1__6_;
  assign new_U6961 = ~new_U2546 | ~INSTQUEUE_REG_0__6_;
  assign new_U6962 = ~new_U4029 | ~new_U4030 | ~new_U4032 | ~new_U4031;
  assign new_U6963 = ~new_U2564 | ~INSTQUEUE_REG_15__5_;
  assign new_U6964 = ~new_U2563 | ~INSTQUEUE_REG_14__5_;
  assign new_U6965 = ~new_U2562 | ~INSTQUEUE_REG_13__5_;
  assign new_U6966 = ~new_U2561 | ~INSTQUEUE_REG_12__5_;
  assign new_U6967 = ~new_U2559 | ~INSTQUEUE_REG_11__5_;
  assign new_U6968 = ~new_U2558 | ~INSTQUEUE_REG_10__5_;
  assign new_U6969 = ~new_U2557 | ~INSTQUEUE_REG_9__5_;
  assign new_U6970 = ~new_U2556 | ~INSTQUEUE_REG_8__5_;
  assign new_U6971 = ~new_U2554 | ~INSTQUEUE_REG_7__5_;
  assign new_U6972 = ~new_U2553 | ~INSTQUEUE_REG_6__5_;
  assign new_U6973 = ~new_U2552 | ~INSTQUEUE_REG_5__5_;
  assign new_U6974 = ~new_U2551 | ~INSTQUEUE_REG_4__5_;
  assign new_U6975 = ~new_U2549 | ~INSTQUEUE_REG_3__5_;
  assign new_U6976 = ~new_U2548 | ~INSTQUEUE_REG_2__5_;
  assign new_U6977 = ~new_U2547 | ~INSTQUEUE_REG_1__5_;
  assign new_U6978 = ~new_U2546 | ~INSTQUEUE_REG_0__5_;
  assign new_U6979 = ~new_U4033 | ~new_U4034 | ~new_U4036 | ~new_U4035;
  assign new_U6980 = ~new_U2564 | ~INSTQUEUE_REG_15__4_;
  assign new_U6981 = ~new_U2563 | ~INSTQUEUE_REG_14__4_;
  assign new_U6982 = ~new_U2562 | ~INSTQUEUE_REG_13__4_;
  assign new_U6983 = ~new_U2561 | ~INSTQUEUE_REG_12__4_;
  assign new_U6984 = ~new_U2559 | ~INSTQUEUE_REG_11__4_;
  assign new_U6985 = ~new_U2558 | ~INSTQUEUE_REG_10__4_;
  assign new_U6986 = ~new_U2557 | ~INSTQUEUE_REG_9__4_;
  assign new_U6987 = ~new_U2556 | ~INSTQUEUE_REG_8__4_;
  assign new_U6988 = ~new_U2554 | ~INSTQUEUE_REG_7__4_;
  assign new_U6989 = ~new_U2553 | ~INSTQUEUE_REG_6__4_;
  assign new_U6990 = ~new_U2552 | ~INSTQUEUE_REG_5__4_;
  assign new_U6991 = ~new_U2551 | ~INSTQUEUE_REG_4__4_;
  assign new_U6992 = ~new_U2549 | ~INSTQUEUE_REG_3__4_;
  assign new_U6993 = ~new_U2548 | ~INSTQUEUE_REG_2__4_;
  assign new_U6994 = ~new_U2547 | ~INSTQUEUE_REG_1__4_;
  assign new_U6995 = ~new_U2564 | ~INSTQUEUE_REG_15__3_;
  assign new_U6996 = ~new_U2563 | ~INSTQUEUE_REG_14__3_;
  assign new_U6997 = ~new_U2562 | ~INSTQUEUE_REG_13__3_;
  assign new_U6998 = ~new_U2561 | ~INSTQUEUE_REG_12__3_;
  assign new_U6999 = ~new_U2559 | ~INSTQUEUE_REG_11__3_;
  assign new_U7000 = ~new_U2558 | ~INSTQUEUE_REG_10__3_;
  assign new_U7001 = ~new_U2557 | ~INSTQUEUE_REG_9__3_;
  assign new_U7002 = ~new_U2556 | ~INSTQUEUE_REG_8__3_;
  assign new_U7003 = ~new_U2554 | ~INSTQUEUE_REG_7__3_;
  assign new_U7004 = ~new_U2553 | ~INSTQUEUE_REG_6__3_;
  assign new_U7005 = ~new_U2552 | ~INSTQUEUE_REG_5__3_;
  assign new_U7006 = ~new_U2551 | ~INSTQUEUE_REG_4__3_;
  assign new_U7007 = ~new_U2549 | ~INSTQUEUE_REG_3__3_;
  assign new_U7008 = ~new_U2548 | ~INSTQUEUE_REG_2__3_;
  assign new_U7009 = ~new_U2547 | ~INSTQUEUE_REG_1__3_;
  assign new_U7010 = ~new_U2546 | ~INSTQUEUE_REG_0__3_;
  assign new_U7011 = ~new_U4041 | ~new_U4042 | ~new_U4044 | ~new_U4043;
  assign new_U7012 = ~new_U2564 | ~INSTQUEUE_REG_15__2_;
  assign new_U7013 = ~new_U2563 | ~INSTQUEUE_REG_14__2_;
  assign new_U7014 = ~new_U2562 | ~INSTQUEUE_REG_13__2_;
  assign new_U7015 = ~new_U2561 | ~INSTQUEUE_REG_12__2_;
  assign new_U7016 = ~new_U2559 | ~INSTQUEUE_REG_11__2_;
  assign new_U7017 = ~new_U2558 | ~INSTQUEUE_REG_10__2_;
  assign new_U7018 = ~new_U2557 | ~INSTQUEUE_REG_9__2_;
  assign new_U7019 = ~new_U2556 | ~INSTQUEUE_REG_8__2_;
  assign new_U7020 = ~new_U2554 | ~INSTQUEUE_REG_7__2_;
  assign new_U7021 = ~new_U2553 | ~INSTQUEUE_REG_6__2_;
  assign new_U7022 = ~new_U2552 | ~INSTQUEUE_REG_5__2_;
  assign new_U7023 = ~new_U2551 | ~INSTQUEUE_REG_4__2_;
  assign new_U7024 = ~new_U2549 | ~INSTQUEUE_REG_3__2_;
  assign new_U7025 = ~new_U2548 | ~INSTQUEUE_REG_2__2_;
  assign new_U7026 = ~new_U2547 | ~INSTQUEUE_REG_1__2_;
  assign new_U7027 = ~new_U2546 | ~INSTQUEUE_REG_0__2_;
  assign new_U7028 = ~new_U4045 | ~new_U4046 | ~new_U4048 | ~new_U4047;
  assign new_U7029 = ~new_U4195 | ~new_U3215;
  assign new_U7030 = ~new_SUB_357_U7 | ~new_U2355;
  assign new_U7031 = ~new_R2182_U33 | ~new_U3281;
  assign new_U7032 = ~new_U4195 | ~new_U3214;
  assign new_U7033 = ~new_SUB_357_U10 | ~new_U2355;
  assign new_U7034 = ~new_R2182_U34 | ~new_U3281;
  assign new_U7035 = ~new_U4194 | ~new_U3221;
  assign new_U7036 = ~new_U4180 | ~INSTQUEUE_REG_0__7_;
  assign new_U7037 = ~new_U4194 | ~new_U3220;
  assign new_U7038 = ~new_U4180 | ~INSTQUEUE_REG_0__6_;
  assign new_U7039 = ~new_U4194 | ~new_U3219;
  assign new_U7040 = ~new_U4180 | ~INSTQUEUE_REG_0__5_;
  assign new_U7041 = ~new_U4194 | ~new_U3218;
  assign new_U7042 = ~new_U4194 | ~new_U3217;
  assign new_U7043 = ~new_U4180 | ~INSTQUEUE_REG_0__3_;
  assign new_U7044 = ~new_U4194 | ~new_U3216;
  assign new_U7045 = ~new_U4180 | ~INSTQUEUE_REG_0__2_;
  assign new_U7046 = ~new_U4194 | ~new_U3215;
  assign new_U7047 = ~new_U4180 | ~INSTQUEUE_REG_0__1_;
  assign new_U7048 = ~new_U4194 | ~new_U3214;
  assign new_U7049 = ~new_U3221 | ~new_U4388;
  assign new_U7050 = ~new_U4180 | ~INSTQUEUE_REG_0__0_;
  assign new_U7051 = ~new_U3415 | ~new_U3414;
  assign new_U7052 = ~INSTQUEUERD_ADDR_REG_3_ | ~new_U3251;
  assign new_U7053 = ~new_U3432;
  assign new_U7054 = ~new_U2582 | ~INSTQUEUE_REG_8__7_;
  assign new_U7055 = ~new_U2581 | ~INSTQUEUE_REG_9__7_;
  assign new_U7056 = ~new_U2580 | ~INSTQUEUE_REG_10__7_;
  assign new_U7057 = ~new_U2579 | ~INSTQUEUE_REG_11__7_;
  assign new_U7058 = ~new_U2577 | ~INSTQUEUE_REG_12__7_;
  assign new_U7059 = ~new_U2576 | ~INSTQUEUE_REG_13__7_;
  assign new_U7060 = ~new_U2575 | ~INSTQUEUE_REG_14__7_;
  assign new_U7061 = ~new_U2574 | ~INSTQUEUE_REG_15__7_;
  assign new_U7062 = ~new_U2573 | ~INSTQUEUE_REG_0__7_;
  assign new_U7063 = ~new_U2572 | ~INSTQUEUE_REG_1__7_;
  assign new_U7064 = ~new_U2571 | ~INSTQUEUE_REG_2__7_;
  assign new_U7065 = ~new_U2570 | ~INSTQUEUE_REG_3__7_;
  assign new_U7066 = ~new_U2568 | ~INSTQUEUE_REG_4__7_;
  assign new_U7067 = ~new_U2567 | ~INSTQUEUE_REG_5__7_;
  assign new_U7068 = ~new_U2566 | ~INSTQUEUE_REG_6__7_;
  assign new_U7069 = ~new_U2565 | ~INSTQUEUE_REG_7__7_;
  assign new_U7070 = ~new_U4051 | ~new_U4052 | ~new_U4054 | ~new_U4053;
  assign new_U7071 = ~new_U3412 | ~new_U3408;
  assign new_U7072 = ~new_U4061 | ~new_U4179;
  assign new_U7073 = ~new_U7072 | ~new_U3409;
  assign new_U7074 = ~new_U4491 | ~new_U3265;
  assign new_U7075 = ~new_U3232;
  assign new_U7076 = ~new_U3381 | ~new_U4142 | ~new_U4388 | ~new_U4491;
  assign new_U7077 = ~new_U4177 | ~STATE2_REG_0_;
  assign new_U7078 = ~new_U4055 | ~new_U3232;
  assign new_U7079 = ~new_U3438;
  assign new_U7080 = ~new_U7617 | ~new_U3438 | ~new_U5480;
  assign new_U7081 = ~new_U4182 | ~new_U7080;
  assign new_U7082 = ~new_U3437;
  assign new_U7083 = ~INSTQUEUEWR_ADDR_REG_3_ | ~new_U3284;
  assign new_U7084 = ~INSTQUEUERD_ADDR_REG_3_ | ~new_U3437;
  assign new_U7085 = ~new_U4191 | ~new_U3347;
  assign new_U7086 = ~new_U2582 | ~INSTQUEUE_REG_8__6_;
  assign new_U7087 = ~new_U2581 | ~INSTQUEUE_REG_9__6_;
  assign new_U7088 = ~new_U2580 | ~INSTQUEUE_REG_10__6_;
  assign new_U7089 = ~new_U2579 | ~INSTQUEUE_REG_11__6_;
  assign new_U7090 = ~new_U2577 | ~INSTQUEUE_REG_12__6_;
  assign new_U7091 = ~new_U2576 | ~INSTQUEUE_REG_13__6_;
  assign new_U7092 = ~new_U2575 | ~INSTQUEUE_REG_14__6_;
  assign new_U7093 = ~new_U2574 | ~INSTQUEUE_REG_15__6_;
  assign new_U7094 = ~new_U2573 | ~INSTQUEUE_REG_0__6_;
  assign new_U7095 = ~new_U2572 | ~INSTQUEUE_REG_1__6_;
  assign new_U7096 = ~new_U2571 | ~INSTQUEUE_REG_2__6_;
  assign new_U7097 = ~new_U2570 | ~INSTQUEUE_REG_3__6_;
  assign new_U7098 = ~new_U2568 | ~INSTQUEUE_REG_4__6_;
  assign new_U7099 = ~new_U2567 | ~INSTQUEUE_REG_5__6_;
  assign new_U7100 = ~new_U2566 | ~INSTQUEUE_REG_6__6_;
  assign new_U7101 = ~new_U2565 | ~INSTQUEUE_REG_7__6_;
  assign new_U7102 = ~new_U4067 | ~new_U4068 | ~new_U4070 | ~new_U4069;
  assign new_U7103 = ~new_U2582 | ~INSTQUEUE_REG_8__5_;
  assign new_U7104 = ~new_U2581 | ~INSTQUEUE_REG_9__5_;
  assign new_U7105 = ~new_U2580 | ~INSTQUEUE_REG_10__5_;
  assign new_U7106 = ~new_U2579 | ~INSTQUEUE_REG_11__5_;
  assign new_U7107 = ~new_U2577 | ~INSTQUEUE_REG_12__5_;
  assign new_U7108 = ~new_U2576 | ~INSTQUEUE_REG_13__5_;
  assign new_U7109 = ~new_U2575 | ~INSTQUEUE_REG_14__5_;
  assign new_U7110 = ~new_U2574 | ~INSTQUEUE_REG_15__5_;
  assign new_U7111 = ~new_U2573 | ~INSTQUEUE_REG_0__5_;
  assign new_U7112 = ~new_U2572 | ~INSTQUEUE_REG_1__5_;
  assign new_U7113 = ~new_U2571 | ~INSTQUEUE_REG_2__5_;
  assign new_U7114 = ~new_U2570 | ~INSTQUEUE_REG_3__5_;
  assign new_U7115 = ~new_U2568 | ~INSTQUEUE_REG_4__5_;
  assign new_U7116 = ~new_U2567 | ~INSTQUEUE_REG_5__5_;
  assign new_U7117 = ~new_U2566 | ~INSTQUEUE_REG_6__5_;
  assign new_U7118 = ~new_U2565 | ~INSTQUEUE_REG_7__5_;
  assign new_U7119 = ~new_U4071 | ~new_U4072 | ~new_U4074 | ~new_U4073;
  assign new_U7120 = ~new_U2582 | ~INSTQUEUE_REG_8__4_;
  assign new_U7121 = ~new_U2581 | ~INSTQUEUE_REG_9__4_;
  assign new_U7122 = ~new_U2580 | ~INSTQUEUE_REG_10__4_;
  assign new_U7123 = ~new_U2579 | ~INSTQUEUE_REG_11__4_;
  assign new_U7124 = ~new_U2577 | ~INSTQUEUE_REG_12__4_;
  assign new_U7125 = ~new_U2576 | ~INSTQUEUE_REG_13__4_;
  assign new_U7126 = ~new_U2575 | ~INSTQUEUE_REG_14__4_;
  assign new_U7127 = ~new_U2574 | ~INSTQUEUE_REG_15__4_;
  assign new_U7128 = ~new_U2572 | ~INSTQUEUE_REG_1__4_;
  assign new_U7129 = ~new_U2571 | ~INSTQUEUE_REG_2__4_;
  assign new_U7130 = ~new_U2570 | ~INSTQUEUE_REG_3__4_;
  assign new_U7131 = ~new_U2568 | ~INSTQUEUE_REG_4__4_;
  assign new_U7132 = ~new_U2567 | ~INSTQUEUE_REG_5__4_;
  assign new_U7133 = ~new_U2566 | ~INSTQUEUE_REG_6__4_;
  assign new_U7134 = ~new_U2565 | ~INSTQUEUE_REG_7__4_;
  assign new_U7135 = ~new_U2582 | ~INSTQUEUE_REG_8__3_;
  assign new_U7136 = ~new_U2581 | ~INSTQUEUE_REG_9__3_;
  assign new_U7137 = ~new_U2580 | ~INSTQUEUE_REG_10__3_;
  assign new_U7138 = ~new_U2579 | ~INSTQUEUE_REG_11__3_;
  assign new_U7139 = ~new_U2577 | ~INSTQUEUE_REG_12__3_;
  assign new_U7140 = ~new_U2576 | ~INSTQUEUE_REG_13__3_;
  assign new_U7141 = ~new_U2575 | ~INSTQUEUE_REG_14__3_;
  assign new_U7142 = ~new_U2574 | ~INSTQUEUE_REG_15__3_;
  assign new_U7143 = ~new_U2573 | ~INSTQUEUE_REG_0__3_;
  assign new_U7144 = ~new_U2572 | ~INSTQUEUE_REG_1__3_;
  assign new_U7145 = ~new_U2571 | ~INSTQUEUE_REG_2__3_;
  assign new_U7146 = ~new_U2570 | ~INSTQUEUE_REG_3__3_;
  assign new_U7147 = ~new_U2568 | ~INSTQUEUE_REG_4__3_;
  assign new_U7148 = ~new_U2567 | ~INSTQUEUE_REG_5__3_;
  assign new_U7149 = ~new_U2566 | ~INSTQUEUE_REG_6__3_;
  assign new_U7150 = ~new_U2565 | ~INSTQUEUE_REG_7__3_;
  assign new_U7151 = ~new_U4080 | ~new_U4081 | ~new_U4083 | ~new_U4082;
  assign new_U7152 = ~new_U2582 | ~INSTQUEUE_REG_8__2_;
  assign new_U7153 = ~new_U2581 | ~INSTQUEUE_REG_9__2_;
  assign new_U7154 = ~new_U2580 | ~INSTQUEUE_REG_10__2_;
  assign new_U7155 = ~new_U2579 | ~INSTQUEUE_REG_11__2_;
  assign new_U7156 = ~new_U2577 | ~INSTQUEUE_REG_12__2_;
  assign new_U7157 = ~new_U2576 | ~INSTQUEUE_REG_13__2_;
  assign new_U7158 = ~new_U2575 | ~INSTQUEUE_REG_14__2_;
  assign new_U7159 = ~new_U2574 | ~INSTQUEUE_REG_15__2_;
  assign new_U7160 = ~new_U2573 | ~INSTQUEUE_REG_0__2_;
  assign new_U7161 = ~new_U2572 | ~INSTQUEUE_REG_1__2_;
  assign new_U7162 = ~new_U2571 | ~INSTQUEUE_REG_2__2_;
  assign new_U7163 = ~new_U2570 | ~INSTQUEUE_REG_3__2_;
  assign new_U7164 = ~new_U2568 | ~INSTQUEUE_REG_4__2_;
  assign new_U7165 = ~new_U2567 | ~INSTQUEUE_REG_5__2_;
  assign new_U7166 = ~new_U2566 | ~INSTQUEUE_REG_6__2_;
  assign new_U7167 = ~new_U2565 | ~INSTQUEUE_REG_7__2_;
  assign new_U7168 = ~new_U4084 | ~new_U4085 | ~new_U4087 | ~new_U4086;
  assign new_U7169 = ~new_U2582 | ~INSTQUEUE_REG_8__1_;
  assign new_U7170 = ~new_U2581 | ~INSTQUEUE_REG_9__1_;
  assign new_U7171 = ~new_U2580 | ~INSTQUEUE_REG_10__1_;
  assign new_U7172 = ~new_U2579 | ~INSTQUEUE_REG_11__1_;
  assign new_U7173 = ~new_U2577 | ~INSTQUEUE_REG_12__1_;
  assign new_U7174 = ~new_U2576 | ~INSTQUEUE_REG_13__1_;
  assign new_U7175 = ~new_U2575 | ~INSTQUEUE_REG_14__1_;
  assign new_U7176 = ~new_U2574 | ~INSTQUEUE_REG_15__1_;
  assign new_U7177 = ~new_U2573 | ~INSTQUEUE_REG_0__1_;
  assign new_U7178 = ~new_U2572 | ~INSTQUEUE_REG_1__1_;
  assign new_U7179 = ~new_U2571 | ~INSTQUEUE_REG_2__1_;
  assign new_U7180 = ~new_U2570 | ~INSTQUEUE_REG_3__1_;
  assign new_U7181 = ~new_U2568 | ~INSTQUEUE_REG_4__1_;
  assign new_U7182 = ~new_U2567 | ~INSTQUEUE_REG_5__1_;
  assign new_U7183 = ~new_U2566 | ~INSTQUEUE_REG_6__1_;
  assign new_U7184 = ~new_U2565 | ~INSTQUEUE_REG_7__1_;
  assign new_U7185 = ~new_U4088 | ~new_U4089 | ~new_U4091 | ~new_U4090;
  assign new_U7186 = ~new_U2582 | ~INSTQUEUE_REG_8__0_;
  assign new_U7187 = ~new_U2581 | ~INSTQUEUE_REG_9__0_;
  assign new_U7188 = ~new_U2580 | ~INSTQUEUE_REG_10__0_;
  assign new_U7189 = ~new_U2579 | ~INSTQUEUE_REG_11__0_;
  assign new_U7190 = ~new_U2577 | ~INSTQUEUE_REG_12__0_;
  assign new_U7191 = ~new_U2576 | ~INSTQUEUE_REG_13__0_;
  assign new_U7192 = ~new_U2575 | ~INSTQUEUE_REG_14__0_;
  assign new_U7193 = ~new_U2574 | ~INSTQUEUE_REG_15__0_;
  assign new_U7194 = ~new_U2573 | ~INSTQUEUE_REG_0__0_;
  assign new_U7195 = ~new_U2572 | ~INSTQUEUE_REG_1__0_;
  assign new_U7196 = ~new_U2571 | ~INSTQUEUE_REG_2__0_;
  assign new_U7197 = ~new_U2570 | ~INSTQUEUE_REG_3__0_;
  assign new_U7198 = ~new_U2568 | ~INSTQUEUE_REG_4__0_;
  assign new_U7199 = ~new_U2567 | ~INSTQUEUE_REG_5__0_;
  assign new_U7200 = ~new_U2566 | ~INSTQUEUE_REG_6__0_;
  assign new_U7201 = ~new_U2565 | ~INSTQUEUE_REG_7__0_;
  assign new_U7202 = ~new_U4092 | ~new_U4093 | ~new_U4095 | ~new_U4094;
  assign new_U7203 = ~INSTQUEUEWR_ADDR_REG_2_ | ~new_U3284;
  assign new_U7204 = ~new_U4191 | ~new_U3442;
  assign new_U7205 = ~INSTQUEUEWR_ADDR_REG_1_ | ~new_U3284;
  assign new_U7206 = ~new_U4191 | ~new_U3222;
  assign new_U7207 = ~new_U4171;
  assign new_U7208 = ~new_U2602 | ~INSTQUEUE_REG_8__7_;
  assign new_U7209 = ~new_U2601 | ~INSTQUEUE_REG_9__7_;
  assign new_U7210 = ~new_U2600 | ~INSTQUEUE_REG_10__7_;
  assign new_U7211 = ~new_U2599 | ~INSTQUEUE_REG_11__7_;
  assign new_U7212 = ~new_U2597 | ~INSTQUEUE_REG_12__7_;
  assign new_U7213 = ~new_U2596 | ~INSTQUEUE_REG_13__7_;
  assign new_U7214 = ~new_U2595 | ~INSTQUEUE_REG_14__7_;
  assign new_U7215 = ~new_U2594 | ~INSTQUEUE_REG_15__7_;
  assign new_U7216 = ~new_U2592 | ~INSTQUEUE_REG_0__7_;
  assign new_U7217 = ~new_U2591 | ~INSTQUEUE_REG_1__7_;
  assign new_U7218 = ~new_U2590 | ~INSTQUEUE_REG_2__7_;
  assign new_U7219 = ~new_U2589 | ~INSTQUEUE_REG_3__7_;
  assign new_U7220 = ~new_U2587 | ~INSTQUEUE_REG_4__7_;
  assign new_U7221 = ~new_U2586 | ~INSTQUEUE_REG_5__7_;
  assign new_U7222 = ~new_U2585 | ~INSTQUEUE_REG_6__7_;
  assign new_U7223 = ~new_U2584 | ~INSTQUEUE_REG_7__7_;
  assign new_U7224 = ~new_U4109 | ~new_U4110 | ~new_U4112 | ~new_U4111;
  assign new_U7225 = ~new_U2602 | ~INSTQUEUE_REG_8__6_;
  assign new_U7226 = ~new_U2601 | ~INSTQUEUE_REG_9__6_;
  assign new_U7227 = ~new_U2600 | ~INSTQUEUE_REG_10__6_;
  assign new_U7228 = ~new_U2599 | ~INSTQUEUE_REG_11__6_;
  assign new_U7229 = ~new_U2597 | ~INSTQUEUE_REG_12__6_;
  assign new_U7230 = ~new_U2596 | ~INSTQUEUE_REG_13__6_;
  assign new_U7231 = ~new_U2595 | ~INSTQUEUE_REG_14__6_;
  assign new_U7232 = ~new_U2594 | ~INSTQUEUE_REG_15__6_;
  assign new_U7233 = ~new_U2592 | ~INSTQUEUE_REG_0__6_;
  assign new_U7234 = ~new_U2591 | ~INSTQUEUE_REG_1__6_;
  assign new_U7235 = ~new_U2590 | ~INSTQUEUE_REG_2__6_;
  assign new_U7236 = ~new_U2589 | ~INSTQUEUE_REG_3__6_;
  assign new_U7237 = ~new_U2587 | ~INSTQUEUE_REG_4__6_;
  assign new_U7238 = ~new_U2586 | ~INSTQUEUE_REG_5__6_;
  assign new_U7239 = ~new_U2585 | ~INSTQUEUE_REG_6__6_;
  assign new_U7240 = ~new_U2584 | ~INSTQUEUE_REG_7__6_;
  assign new_U7241 = ~new_U4113 | ~new_U4114 | ~new_U4116 | ~new_U4115;
  assign new_U7242 = ~new_U2602 | ~INSTQUEUE_REG_8__5_;
  assign new_U7243 = ~new_U2601 | ~INSTQUEUE_REG_9__5_;
  assign new_U7244 = ~new_U2600 | ~INSTQUEUE_REG_10__5_;
  assign new_U7245 = ~new_U2599 | ~INSTQUEUE_REG_11__5_;
  assign new_U7246 = ~new_U2597 | ~INSTQUEUE_REG_12__5_;
  assign new_U7247 = ~new_U2596 | ~INSTQUEUE_REG_13__5_;
  assign new_U7248 = ~new_U2595 | ~INSTQUEUE_REG_14__5_;
  assign new_U7249 = ~new_U2594 | ~INSTQUEUE_REG_15__5_;
  assign new_U7250 = ~new_U2592 | ~INSTQUEUE_REG_0__5_;
  assign new_U7251 = ~new_U2591 | ~INSTQUEUE_REG_1__5_;
  assign new_U7252 = ~new_U2590 | ~INSTQUEUE_REG_2__5_;
  assign new_U7253 = ~new_U2589 | ~INSTQUEUE_REG_3__5_;
  assign new_U7254 = ~new_U2587 | ~INSTQUEUE_REG_4__5_;
  assign new_U7255 = ~new_U2586 | ~INSTQUEUE_REG_5__5_;
  assign new_U7256 = ~new_U2585 | ~INSTQUEUE_REG_6__5_;
  assign new_U7257 = ~new_U2584 | ~INSTQUEUE_REG_7__5_;
  assign new_U7258 = ~new_U4117 | ~new_U4118 | ~new_U4120 | ~new_U4119;
  assign new_U7259 = ~new_U2602 | ~INSTQUEUE_REG_8__4_;
  assign new_U7260 = ~new_U2601 | ~INSTQUEUE_REG_9__4_;
  assign new_U7261 = ~new_U2600 | ~INSTQUEUE_REG_10__4_;
  assign new_U7262 = ~new_U2599 | ~INSTQUEUE_REG_11__4_;
  assign new_U7263 = ~new_U2597 | ~INSTQUEUE_REG_12__4_;
  assign new_U7264 = ~new_U2596 | ~INSTQUEUE_REG_13__4_;
  assign new_U7265 = ~new_U2595 | ~INSTQUEUE_REG_14__4_;
  assign new_U7266 = ~new_U2594 | ~INSTQUEUE_REG_15__4_;
  assign new_U7267 = ~new_U2591 | ~INSTQUEUE_REG_1__4_;
  assign new_U7268 = ~new_U2590 | ~INSTQUEUE_REG_2__4_;
  assign new_U7269 = ~new_U2589 | ~INSTQUEUE_REG_3__4_;
  assign new_U7270 = ~new_U2587 | ~INSTQUEUE_REG_4__4_;
  assign new_U7271 = ~new_U2586 | ~INSTQUEUE_REG_5__4_;
  assign new_U7272 = ~new_U2585 | ~INSTQUEUE_REG_6__4_;
  assign new_U7273 = ~new_U2584 | ~INSTQUEUE_REG_7__4_;
  assign new_U7274 = ~new_U2602 | ~INSTQUEUE_REG_8__3_;
  assign new_U7275 = ~new_U2601 | ~INSTQUEUE_REG_9__3_;
  assign new_U7276 = ~new_U2600 | ~INSTQUEUE_REG_10__3_;
  assign new_U7277 = ~new_U2599 | ~INSTQUEUE_REG_11__3_;
  assign new_U7278 = ~new_U2597 | ~INSTQUEUE_REG_12__3_;
  assign new_U7279 = ~new_U2596 | ~INSTQUEUE_REG_13__3_;
  assign new_U7280 = ~new_U2595 | ~INSTQUEUE_REG_14__3_;
  assign new_U7281 = ~new_U2594 | ~INSTQUEUE_REG_15__3_;
  assign new_U7282 = ~new_U2592 | ~INSTQUEUE_REG_0__3_;
  assign new_U7283 = ~new_U2591 | ~INSTQUEUE_REG_1__3_;
  assign new_U7284 = ~new_U2590 | ~INSTQUEUE_REG_2__3_;
  assign new_U7285 = ~new_U2589 | ~INSTQUEUE_REG_3__3_;
  assign new_U7286 = ~new_U2587 | ~INSTQUEUE_REG_4__3_;
  assign new_U7287 = ~new_U2586 | ~INSTQUEUE_REG_5__3_;
  assign new_U7288 = ~new_U2585 | ~INSTQUEUE_REG_6__3_;
  assign new_U7289 = ~new_U2584 | ~INSTQUEUE_REG_7__3_;
  assign new_U7290 = ~new_U4125 | ~new_U4126 | ~new_U4128 | ~new_U4127;
  assign new_U7291 = ~new_U2602 | ~INSTQUEUE_REG_8__2_;
  assign new_U7292 = ~new_U2601 | ~INSTQUEUE_REG_9__2_;
  assign new_U7293 = ~new_U2600 | ~INSTQUEUE_REG_10__2_;
  assign new_U7294 = ~new_U2599 | ~INSTQUEUE_REG_11__2_;
  assign new_U7295 = ~new_U2597 | ~INSTQUEUE_REG_12__2_;
  assign new_U7296 = ~new_U2596 | ~INSTQUEUE_REG_13__2_;
  assign new_U7297 = ~new_U2595 | ~INSTQUEUE_REG_14__2_;
  assign new_U7298 = ~new_U2594 | ~INSTQUEUE_REG_15__2_;
  assign new_U7299 = ~new_U2592 | ~INSTQUEUE_REG_0__2_;
  assign new_U7300 = ~new_U2591 | ~INSTQUEUE_REG_1__2_;
  assign new_U7301 = ~new_U2590 | ~INSTQUEUE_REG_2__2_;
  assign new_U7302 = ~new_U2589 | ~INSTQUEUE_REG_3__2_;
  assign new_U7303 = ~new_U2587 | ~INSTQUEUE_REG_4__2_;
  assign new_U7304 = ~new_U2586 | ~INSTQUEUE_REG_5__2_;
  assign new_U7305 = ~new_U2585 | ~INSTQUEUE_REG_6__2_;
  assign new_U7306 = ~new_U2584 | ~INSTQUEUE_REG_7__2_;
  assign new_U7307 = ~new_U4129 | ~new_U4130 | ~new_U4132 | ~new_U4131;
  assign new_U7308 = ~new_U2602 | ~INSTQUEUE_REG_8__1_;
  assign new_U7309 = ~new_U2601 | ~INSTQUEUE_REG_9__1_;
  assign new_U7310 = ~new_U2600 | ~INSTQUEUE_REG_10__1_;
  assign new_U7311 = ~new_U2599 | ~INSTQUEUE_REG_11__1_;
  assign new_U7312 = ~new_U2597 | ~INSTQUEUE_REG_12__1_;
  assign new_U7313 = ~new_U2596 | ~INSTQUEUE_REG_13__1_;
  assign new_U7314 = ~new_U2595 | ~INSTQUEUE_REG_14__1_;
  assign new_U7315 = ~new_U2594 | ~INSTQUEUE_REG_15__1_;
  assign new_U7316 = ~new_U2592 | ~INSTQUEUE_REG_0__1_;
  assign new_U7317 = ~new_U2591 | ~INSTQUEUE_REG_1__1_;
  assign new_U7318 = ~new_U2590 | ~INSTQUEUE_REG_2__1_;
  assign new_U7319 = ~new_U2589 | ~INSTQUEUE_REG_3__1_;
  assign new_U7320 = ~new_U2587 | ~INSTQUEUE_REG_4__1_;
  assign new_U7321 = ~new_U2586 | ~INSTQUEUE_REG_5__1_;
  assign new_U7322 = ~new_U2585 | ~INSTQUEUE_REG_6__1_;
  assign new_U7323 = ~new_U2584 | ~INSTQUEUE_REG_7__1_;
  assign new_U7324 = ~new_U4133 | ~new_U4134 | ~new_U4136 | ~new_U4135;
  assign new_U7325 = ~new_U2602 | ~INSTQUEUE_REG_8__0_;
  assign new_U7326 = ~new_U2601 | ~INSTQUEUE_REG_9__0_;
  assign new_U7327 = ~new_U2600 | ~INSTQUEUE_REG_10__0_;
  assign new_U7328 = ~new_U2599 | ~INSTQUEUE_REG_11__0_;
  assign new_U7329 = ~new_U2597 | ~INSTQUEUE_REG_12__0_;
  assign new_U7330 = ~new_U2596 | ~INSTQUEUE_REG_13__0_;
  assign new_U7331 = ~new_U2595 | ~INSTQUEUE_REG_14__0_;
  assign new_U7332 = ~new_U2594 | ~INSTQUEUE_REG_15__0_;
  assign new_U7333 = ~new_U2592 | ~INSTQUEUE_REG_0__0_;
  assign new_U7334 = ~new_U2591 | ~INSTQUEUE_REG_1__0_;
  assign new_U7335 = ~new_U2590 | ~INSTQUEUE_REG_2__0_;
  assign new_U7336 = ~new_U2589 | ~INSTQUEUE_REG_3__0_;
  assign new_U7337 = ~new_U2587 | ~INSTQUEUE_REG_4__0_;
  assign new_U7338 = ~new_U2586 | ~INSTQUEUE_REG_5__0_;
  assign new_U7339 = ~new_U2585 | ~INSTQUEUE_REG_6__0_;
  assign new_U7340 = ~new_U2584 | ~INSTQUEUE_REG_7__0_;
  assign new_U7341 = ~new_U4137 | ~new_U4138 | ~new_U4140 | ~new_U4139;
  assign new_U7342 = ~new_U4222 | ~new_U4219 | ~new_U2354;
  assign new_U7343 = ~new_U4141 | ~new_U7075;
  assign new_U7344 = ~new_U3383 | ~new_U3397;
  assign new_U7345 = ~new_U4222 | ~new_U7344;
  assign new_U7346 = ~new_U4178 | ~new_U2452;
  assign new_U7347 = ~new_U7343 | ~new_U3258;
  assign new_U7348 = ~new_U4196 | ~new_U7076;
  assign new_U7349 = ~new_U4148 | ~new_U4196;
  assign new_U7350 = ~new_U2451 | ~new_U4198;
  assign new_U7351 = ~new_U7349 | ~new_U7350 | ~new_U4183 | ~new_U3407 | ~new_U3421;
  assign new_U7352 = ~new_R2238_U6 | ~new_U7351;
  assign new_U7353 = ~new_SUB_450_U6 | ~new_U2354;
  assign new_U7354 = ~new_R2238_U19 | ~new_U7351;
  assign new_U7355 = ~new_SUB_450_U19 | ~new_U2354;
  assign new_U7356 = ~new_R2238_U20 | ~new_U7351;
  assign new_U7357 = ~new_SUB_450_U20 | ~new_U2354;
  assign new_U7358 = ~new_R2238_U21 | ~new_U7351;
  assign new_U7359 = ~new_SUB_450_U21 | ~new_U2354;
  assign new_U7360 = ~new_R2238_U22 | ~new_U7351;
  assign new_U7361 = ~new_SUB_450_U22 | ~new_U2354;
  assign new_U7362 = ~new_R2238_U7 | ~new_U7351;
  assign new_U7363 = ~new_SUB_450_U7 | ~new_U2354;
  assign new_U7364 = ~new_R2238_U19 | ~new_U4180;
  assign new_U7365 = ~INSTQUEUERD_ADDR_REG_4_ | ~new_U3281;
  assign new_U7366 = ~new_R2238_U20 | ~new_U4180;
  assign new_U7367 = ~INSTQUEUERD_ADDR_REG_3_ | ~new_U3281;
  assign new_U7368 = ~STATE2_REG_0_ | ~new_U4161;
  assign new_U7369 = ~new_U3407 | ~new_U7368;
  assign new_U7370 = ~new_R2238_U21 | ~new_U4180;
  assign new_U7371 = ~INSTQUEUERD_ADDR_REG_2_ | ~new_U3281;
  assign new_U7372 = ~new_U2450 | ~new_U3258;
  assign new_U7373 = ~new_R2238_U22 | ~new_U4180;
  assign new_U7374 = ~INSTQUEUERD_ADDR_REG_1_ | ~new_U3281;
  assign new_U7375 = ~new_U2451 | ~new_U3271;
  assign new_U7376 = ~new_R2238_U7 | ~new_U4180;
  assign new_U7377 = ~INSTQUEUERD_ADDR_REG_0_ | ~new_U3281;
  assign new_U7378 = ~new_U3380 | ~new_U3277;
  assign new_U7379 = ~new_U3271 | ~new_U3436;
  assign new_U7380 = ~INSTADDRPOINTER_REG_9_ | ~new_U7379;
  assign new_U7381 = ~EBX_REG_9_ | ~new_U7378;
  assign new_U7382 = ~INSTADDRPOINTER_REG_8_ | ~new_U7379;
  assign new_U7383 = ~EBX_REG_8_ | ~new_U7378;
  assign new_U7384 = ~INSTADDRPOINTER_REG_7_ | ~new_U7379;
  assign new_U7385 = ~EBX_REG_7_ | ~new_U7378;
  assign new_U7386 = ~INSTADDRPOINTER_REG_6_ | ~new_U7379;
  assign new_U7387 = ~EBX_REG_6_ | ~new_U7378;
  assign new_U7388 = ~INSTADDRPOINTER_REG_5_ | ~new_U7379;
  assign new_U7389 = ~EBX_REG_5_ | ~new_U7378;
  assign new_U7390 = ~INSTADDRPOINTER_REG_4_ | ~new_U7379;
  assign new_U7391 = ~EBX_REG_4_ | ~new_U7378;
  assign new_U7392 = ~INSTADDRPOINTER_REG_31_ | ~new_U7379;
  assign new_U7393 = ~EBX_REG_31_ | ~new_U7378;
  assign new_U7394 = ~INSTADDRPOINTER_REG_30_ | ~new_U7379;
  assign new_U7395 = ~EBX_REG_30_ | ~new_U7378;
  assign new_U7396 = ~INSTADDRPOINTER_REG_3_ | ~new_U7379;
  assign new_U7397 = ~EBX_REG_3_ | ~new_U7378;
  assign new_U7398 = ~INSTADDRPOINTER_REG_29_ | ~new_U7379;
  assign new_U7399 = ~EBX_REG_29_ | ~new_U7378;
  assign new_U7400 = ~INSTADDRPOINTER_REG_28_ | ~new_U7379;
  assign new_U7401 = ~EBX_REG_28_ | ~new_U7378;
  assign new_U7402 = ~INSTADDRPOINTER_REG_27_ | ~new_U7379;
  assign new_U7403 = ~EBX_REG_27_ | ~new_U7378;
  assign new_U7404 = ~INSTADDRPOINTER_REG_26_ | ~new_U7379;
  assign new_U7405 = ~EBX_REG_26_ | ~new_U7378;
  assign new_U7406 = ~INSTADDRPOINTER_REG_25_ | ~new_U7379;
  assign new_U7407 = ~EBX_REG_25_ | ~new_U7378;
  assign new_U7408 = ~INSTADDRPOINTER_REG_24_ | ~new_U7379;
  assign new_U7409 = ~EBX_REG_24_ | ~new_U7378;
  assign new_U7410 = ~INSTADDRPOINTER_REG_23_ | ~new_U7379;
  assign new_U7411 = ~EBX_REG_23_ | ~new_U7378;
  assign new_U7412 = ~INSTADDRPOINTER_REG_22_ | ~new_U7379;
  assign new_U7413 = ~EBX_REG_22_ | ~new_U7378;
  assign new_U7414 = ~INSTADDRPOINTER_REG_21_ | ~new_U7379;
  assign new_U7415 = ~EBX_REG_21_ | ~new_U7378;
  assign new_U7416 = ~INSTADDRPOINTER_REG_20_ | ~new_U7379;
  assign new_U7417 = ~EBX_REG_20_ | ~new_U7378;
  assign new_U7418 = ~INSTADDRPOINTER_REG_2_ | ~new_U7379;
  assign new_U7419 = ~EBX_REG_2_ | ~new_U7378;
  assign new_U7420 = ~INSTADDRPOINTER_REG_19_ | ~new_U7379;
  assign new_U7421 = ~EBX_REG_19_ | ~new_U7378;
  assign new_U7422 = ~INSTADDRPOINTER_REG_18_ | ~new_U7379;
  assign new_U7423 = ~EBX_REG_18_ | ~new_U7378;
  assign new_U7424 = ~INSTADDRPOINTER_REG_17_ | ~new_U7379;
  assign new_U7425 = ~EBX_REG_17_ | ~new_U7378;
  assign new_U7426 = ~INSTADDRPOINTER_REG_16_ | ~new_U7379;
  assign new_U7427 = ~EBX_REG_16_ | ~new_U7378;
  assign new_U7428 = ~INSTADDRPOINTER_REG_15_ | ~new_U7379;
  assign new_U7429 = ~EBX_REG_15_ | ~new_U7378;
  assign new_U7430 = ~INSTADDRPOINTER_REG_14_ | ~new_U7379;
  assign new_U7431 = ~EBX_REG_14_ | ~new_U7378;
  assign new_U7432 = ~INSTADDRPOINTER_REG_13_ | ~new_U7379;
  assign new_U7433 = ~EBX_REG_13_ | ~new_U7378;
  assign new_U7434 = ~INSTADDRPOINTER_REG_12_ | ~new_U7379;
  assign new_U7435 = ~EBX_REG_12_ | ~new_U7378;
  assign new_U7436 = ~INSTADDRPOINTER_REG_11_ | ~new_U7379;
  assign new_U7437 = ~EBX_REG_11_ | ~new_U7378;
  assign new_U7438 = ~INSTADDRPOINTER_REG_10_ | ~new_U7379;
  assign new_U7439 = ~EBX_REG_10_ | ~new_U7378;
  assign new_U7440 = ~INSTADDRPOINTER_REG_1_ | ~new_U7379;
  assign new_U7441 = ~EBX_REG_1_ | ~new_U7378;
  assign new_U7442 = ~INSTADDRPOINTER_REG_0_ | ~new_U7379;
  assign new_U7443 = ~EBX_REG_0_ | ~new_U7378;
  assign new_U7444 = ~new_U4465 | ~new_U4484;
  assign new_U7445 = ~new_U2430 | ~INSTQUEUERD_ADDR_REG_4_;
  assign new_U7446 = ~new_U3476 | ~new_U3249;
  assign new_U7447 = ~new_U2430 | ~INSTQUEUERD_ADDR_REG_3_;
  assign new_U7448 = ~new_U3477 | ~new_U3249;
  assign new_U7449 = ~new_U3457 | ~FLUSH_REG | ~new_U2446;
  assign new_U7450 = ~new_U2430 | ~INSTQUEUERD_ADDR_REG_2_;
  assign new_U7451 = ~new_U3478 | ~new_U3249;
  assign new_U7452 = ~new_U7700 | ~new_U2446 | ~FLUSH_REG;
  assign new_U7453 = ~new_U2430 | ~INSTQUEUERD_ADDR_REG_1_;
  assign new_U7454 = ~new_U3479 | ~new_U3249;
  assign new_U7455 = ~new_U2430 | ~INSTQUEUERD_ADDR_REG_0_;
  assign new_U7456 = ~STATE_REG_0_ | ~new_U4173;
  assign new_U7457 = READY_N | STATE2_REG_2_;
  assign new_U7458 = ~new_U4098 | ~new_U7206;
  assign new_U7459 = ~new_U7072 | ~new_U3409;
  assign new_U7460 = ~new_U4199 | ~STATE2_REG_0_;
  assign new_U7461 = ~new_U4200 | ~STATE2_REG_0_;
  assign new_U7462 = ~new_U4201 | ~STATE2_REG_0_;
  assign new_U7463 = ~new_U4224 | ~STATE2_REG_0_;
  assign new_U7464 = ~new_U4252 | ~STATE2_REG_0_;
  assign new_U7465 = ~STATE2_REG_0_ | ~new_U7620;
  assign new_U7466 = ~new_U2608 | ~new_U3253;
  assign new_U7467 = ~new_U4108 | ~new_U4106 | ~new_U4105 | ~new_U7081;
  assign new_U7468 = ~STATE2_REG_0_ | ~new_U7620;
  assign new_U7469 = ~new_U2379 | ~new_U3416;
  assign new_U7470 = ~new_U2369 | ~new_U6355;
  assign new_U7471 = ~new_U3876 | ~new_U2369;
  assign new_U7472 = ~new_U7470 | ~new_U7469 | ~new_U4217;
  assign new_U7473 = ~new_U7471 | ~new_U4218;
  assign new_U7474 = ~new_U4182 | ~new_U5479 | ~new_U4159;
  assign new_U7475 = ~new_U7079 | ~new_U4182;
  assign new_U7476 = ~new_U4182 | ~new_U3379;
  assign new_U7477 = ~new_U4224 | ~STATE2_REG_0_;
  assign new_U7478 = ~new_U4060 | ~new_U7773 | ~new_U7772;
  assign new_U7479 = ~new_U4096 | ~new_U7204;
  assign new_U7480 = ~new_U4097 | ~new_U7082;
  assign new_U7481 = ~new_U3266;
  assign new_U7482 = ~new_U3263;
  assign new_U7483 = ~new_U4056 | ~new_U4057 | ~new_U4058 | ~new_U4059 | ~new_U2607;
  assign new_U7484 = ~new_U3722 | ~new_U7481;
  assign new_U7485 = ~new_U3723 | ~new_U5457;
  assign new_U7486 = ~new_U2425 | ~new_U7481;
  assign new_U7487 = ~new_U2425 | ~new_U7481;
  assign new_U7488 = ~new_U7487 | ~new_U6349 | ~new_U6348;
  assign new_U7489 = ~new_U7481 | ~new_R2167_U17;
  assign new_U7490 = ~new_R2167_U17 | ~new_U7481 | ~new_U4189;
  assign new_U7491 = ~new_U7490 | ~new_U6137;
  assign new_U7492 = ~new_U7481 | ~new_U7073;
  assign new_U7493 = ~new_U7481 | ~new_U7459;
  assign new_U7494 = ~new_U4102 | ~new_U4104 | ~new_U4103;
  assign new_U7495 = ~new_U3747 | ~new_U7481;
  assign new_U7496 = ~new_U3748 | ~new_U3749 | ~new_U5553;
  assign new_U7497 = ~new_U3734 | ~new_U2519;
  assign new_U7498 = ~new_U7481 | ~new_U5950;
  assign new_U7499 = ~new_U7481 | ~new_U5953;
  assign new_U7500 = ~new_U7481 | ~new_U5956;
  assign new_U7501 = ~new_U7481 | ~new_U5959;
  assign new_U7502 = ~new_U7481 | ~new_U5962;
  assign new_U7503 = ~new_U7481 | ~new_U5965;
  assign new_U7504 = ~new_U7481 | ~new_U5968;
  assign new_U7505 = ~new_U7481 | ~new_U5971;
  assign new_U7506 = ~new_U7481 | ~new_U5974;
  assign new_U7507 = ~new_U7481 | ~new_U5977;
  assign new_U7508 = ~new_U7481 | ~new_U5980;
  assign new_U7509 = ~new_U7481 | ~new_U5983;
  assign new_U7510 = ~new_U7481 | ~new_U5986;
  assign new_U7511 = ~new_U7481 | ~new_U5989;
  assign new_U7512 = ~new_U7481 | ~new_U5992;
  assign new_U7513 = ~new_U7481 | ~new_U5995;
  assign new_U7514 = ~new_U7481 | ~new_U5998;
  assign new_U7515 = ~new_U7481 | ~new_U6001;
  assign new_U7516 = ~new_U7481 | ~new_U6004;
  assign new_U7517 = ~new_U7481 | ~new_U6007;
  assign new_U7518 = ~new_U7481 | ~new_U6010;
  assign new_U7519 = ~new_U7481 | ~new_U6013;
  assign new_U7520 = ~new_U7481 | ~new_U6016;
  assign new_U7521 = ~new_U7481 | ~new_U6019;
  assign new_U7522 = ~new_U7481 | ~new_U6022;
  assign new_U7523 = ~new_U7481 | ~new_U6025;
  assign new_U7524 = ~new_U7481 | ~new_U6028;
  assign new_U7525 = ~new_U7481 | ~new_U6031;
  assign new_U7526 = ~new_U7481 | ~new_U6034;
  assign new_U7527 = ~new_U7481 | ~new_U6037;
  assign new_U7528 = ~new_U7481 | ~new_U6040;
  assign new_U7529 = ~new_U2357 | ~new_U7481;
  assign new_U7530 = ~UWORD_REG_0_ | ~new_U7529;
  assign new_U7531 = ~new_U2357 | ~new_U7481;
  assign new_U7532 = ~UWORD_REG_1_ | ~new_U7531;
  assign new_U7533 = ~new_U2357 | ~new_U7481;
  assign new_U7534 = ~UWORD_REG_2_ | ~new_U7533;
  assign new_U7535 = ~new_U2357 | ~new_U7481;
  assign new_U7536 = ~UWORD_REG_3_ | ~new_U7535;
  assign new_U7537 = ~new_U2357 | ~new_U7481;
  assign new_U7538 = ~UWORD_REG_4_ | ~new_U7537;
  assign new_U7539 = ~new_U2357 | ~new_U7481;
  assign new_U7540 = ~UWORD_REG_5_ | ~new_U7539;
  assign new_U7541 = ~new_U2357 | ~new_U7481;
  assign new_U7542 = ~UWORD_REG_6_ | ~new_U7541;
  assign new_U7543 = ~new_U2357 | ~new_U7481;
  assign new_U7544 = ~UWORD_REG_7_ | ~new_U7543;
  assign new_U7545 = ~new_U2357 | ~new_U7481;
  assign new_U7546 = ~UWORD_REG_8_ | ~new_U7545;
  assign new_U7547 = ~new_U2357 | ~new_U7481;
  assign new_U7548 = ~UWORD_REG_9_ | ~new_U7547;
  assign new_U7549 = ~new_U2357 | ~new_U7481;
  assign new_U7550 = ~UWORD_REG_10_ | ~new_U7549;
  assign new_U7551 = ~new_U2357 | ~new_U7481;
  assign new_U7552 = ~UWORD_REG_11_ | ~new_U7551;
  assign new_U7553 = ~new_U2357 | ~new_U7481;
  assign new_U7554 = ~UWORD_REG_12_ | ~new_U7553;
  assign new_U7555 = ~new_U2357 | ~new_U7481;
  assign new_U7556 = ~UWORD_REG_13_ | ~new_U7555;
  assign new_U7557 = ~new_U2357 | ~new_U7481;
  assign new_U7558 = ~UWORD_REG_14_ | ~new_U7557;
  assign new_U7559 = ~new_U2357 | ~new_U7481;
  assign new_U7560 = ~LWORD_REG_0_ | ~new_U7559;
  assign new_U7561 = ~new_U2357 | ~new_U7481;
  assign new_U7562 = ~LWORD_REG_1_ | ~new_U7561;
  assign new_U7563 = ~new_U2357 | ~new_U7481;
  assign new_U7564 = ~LWORD_REG_2_ | ~new_U7563;
  assign new_U7565 = ~new_U2357 | ~new_U7481;
  assign new_U7566 = ~LWORD_REG_3_ | ~new_U7565;
  assign new_U7567 = ~new_U2357 | ~new_U7481;
  assign new_U7568 = ~LWORD_REG_4_ | ~new_U7567;
  assign new_U7569 = ~new_U2357 | ~new_U7481;
  assign new_U7570 = ~LWORD_REG_5_ | ~new_U7569;
  assign new_U7571 = ~new_U2357 | ~new_U7481;
  assign new_U7572 = ~LWORD_REG_6_ | ~new_U7571;
  assign new_U7573 = ~new_U2357 | ~new_U7481;
  assign new_U7574 = ~LWORD_REG_7_ | ~new_U7573;
  assign new_U7575 = ~new_U2357 | ~new_U7481;
  assign new_U7576 = ~LWORD_REG_8_ | ~new_U7575;
  assign new_U7577 = ~new_U2357 | ~new_U7481;
  assign new_U7578 = ~LWORD_REG_9_ | ~new_U7577;
  assign new_U7579 = ~new_U2357 | ~new_U7481;
  assign new_U7580 = ~LWORD_REG_10_ | ~new_U7579;
  assign new_U7581 = ~new_U2357 | ~new_U7481;
  assign new_U7582 = ~LWORD_REG_11_ | ~new_U7581;
  assign new_U7583 = ~new_U2357 | ~new_U7481;
  assign new_U7584 = ~LWORD_REG_12_ | ~new_U7583;
  assign new_U7585 = ~new_U2357 | ~new_U7481;
  assign new_U7586 = ~LWORD_REG_13_ | ~new_U7585;
  assign new_U7587 = ~new_U2357 | ~new_U7481;
  assign new_U7588 = ~LWORD_REG_14_ | ~new_U7587;
  assign new_U7589 = ~new_U2357 | ~new_U7481;
  assign new_U7590 = ~LWORD_REG_15_ | ~new_U7589;
  assign new_U7591 = ~new_U4247 | ~new_U7481 | ~new_U3556;
  assign new_U7592 = ~new_U3569 | ~new_U7672 | ~new_U7671;
  assign new_U7593 = ~new_U3855 | ~new_U7481;
  assign new_U7594 = ~new_U7593 | ~new_U3415;
  assign new_U7595 = ~new_U4196 | ~new_U7481;
  assign new_U7596 = ~new_U7595 | ~new_U3434;
  assign new_U7597 = ~new_U3266 | ~new_U3387;
  assign new_U7598 = ~new_U3742 | ~new_U7481;
  assign new_U7599 = ~new_U3743 | ~new_U7598;
  assign new_U7600 = ~INSTQUEUE_REG_0__4_ | ~new_U5404;
  assign new_U7601 = ~new_U2523 | ~INSTQUEUE_REG_0__4_;
  assign new_U7602 = ~new_U2546 | ~INSTQUEUE_REG_0__4_;
  assign new_U7603 = ~new_U4037 | ~new_U4038 | ~new_U4040 | ~new_U4039;
  assign new_U7604 = ~new_U4180 | ~INSTQUEUE_REG_0__4_;
  assign new_U7605 = ~new_U2573 | ~INSTQUEUE_REG_0__4_;
  assign new_U7606 = ~new_U4075 | ~new_U4076 | ~new_U4079 | ~new_U4077;
  assign new_U7607 = ~new_U2592 | ~INSTQUEUE_REG_0__4_;
  assign new_U7608 = ~new_U4121 | ~new_U4122 | ~new_U4124 | ~new_U4123;
  assign new_U7609 = ~new_U3246;
  assign new_U7610 = ~new_U7609 | ~new_U3248;
  assign new_U7611 = ~new_U4346 | ~new_U4349 | ~STATE_REG_1_;
  assign new_U7612 = ~STATE_REG_2_ | ~new_U7456;
  assign new_U7613 = ~STATE_REG_1_ | ~new_U4346;
  assign new_U7614 = ~new_U4490 | ~new_U4498;
  assign new_U7615 = ~new_U5475 | ~new_U4159;
  assign new_U7616 = ~new_U3270 | ~new_U3276;
  assign new_U7617 = ~new_U3379;
  assign new_U7618 = ~new_U4196 | ~new_U7478;
  assign new_U7619 = ~new_U5475 | ~new_U4159;
  assign new_U7620 = ~new_U7619 | ~new_U7618;
  assign new_U7621 = ~BE_N_REG_3_ | ~new_U3236;
  assign new_U7622 = ~BYTEENABLE_REG_3_ | ~new_U4209;
  assign new_U7623 = ~BE_N_REG_2_ | ~new_U3236;
  assign new_U7624 = ~BYTEENABLE_REG_2_ | ~new_U4209;
  assign new_U7625 = ~BE_N_REG_1_ | ~new_U3236;
  assign new_U7626 = ~BYTEENABLE_REG_1_ | ~new_U4209;
  assign new_U7627 = ~BE_N_REG_0_ | ~new_U3236;
  assign new_U7628 = ~BYTEENABLE_REG_0_ | ~new_U4209;
  assign new_U7629 = ~new_U3238 | ~STATE_REG_0_ | ~REQUESTPENDING_REG;
  assign new_U7630 = ~STATE_REG_2_ | ~new_U3246;
  assign new_U7631 = ~new_U7630 | ~new_U7629;
  assign new_U7632 = ~STATE_REG_1_ | ~new_U7612 | ~new_U4349;
  assign new_U7633 = ~new_U7631 | ~new_U3235;
  assign new_U7634 = ~STATE_REG_2_ | ~STATE_REG_0_ | ~new_U3247;
  assign new_U7635 = ~new_U4359 | ~new_U3238;
  assign new_U7636 = STATE_REG_0_ | STATE_REG_1_;
  assign new_U7637 = ~STATE_REG_0_ | ~new_U4246;
  assign new_U7638 = ~new_U3449;
  assign new_U7639 = ~new_U7638 | ~DATAWIDTH_REG_0_;
  assign new_U7640 = ~new_U3450 | ~new_U3449;
  assign new_U7641 = ~new_U3449 | ~new_U4364;
  assign new_U7642 = ~new_U7638 | ~DATAWIDTH_REG_1_;
  assign new_U7643 = ~new_U3252 | ~new_U3529 | ~new_U3528;
  assign new_U7644 = ~INSTQUEUERD_ADDR_REG_1_ | ~new_U3257 | ~INSTQUEUERD_ADDR_REG_2_ | ~INSTQUEUE_REG_7__4_ | ~INSTQUEUERD_ADDR_REG_0_;
  assign new_U7645 = ~new_U3252 | ~new_U3257 | ~INSTQUEUERD_ADDR_REG_2_ | ~INSTQUEUE_REG_5__4_ | ~INSTQUEUERD_ADDR_REG_0_;
  assign new_U7646 = ~INSTQUEUERD_ADDR_REG_1_ | ~new_U3253 | ~new_U3251 | ~INSTQUEUE_REG_2__4_ | ~new_U3257;
  assign new_U7647 = ~new_U3257 | ~new_U3531 | ~new_U3530;
  assign new_U7648 = ~INSTQUEUERD_ADDR_REG_3_ | ~new_U3533 | ~new_U3532;
  assign new_U7649 = ~new_U3252 | ~new_U3535 | ~new_U3534;
  assign new_U7650 = ~INSTQUEUERD_ADDR_REG_1_ | ~new_U3537 | ~new_U3536;
  assign new_U7651 = ~new_U3253 | ~new_U3539 | ~new_U3538;
  assign new_U7652 = ~INSTQUEUERD_ADDR_REG_0_ | ~INSTQUEUERD_ADDR_REG_2_ | ~INSTQUEUERD_ADDR_REG_1_ | ~INSTQUEUE_REG_15__4_ | ~INSTQUEUERD_ADDR_REG_3_;
  assign new_U7653 = ~new_U3257 | ~new_U3253 | ~new_U3252 | ~INSTQUEUE_REG_0__4_ | ~new_U3251;
  assign new_U7654 = ~INSTQUEUERD_ADDR_REG_3_ | ~new_U3253 | ~new_U3252 | ~INSTQUEUE_REG_8__4_ | ~new_U3251;
  assign new_U7655 = ~new_U3253 | ~new_U3251 | ~INSTQUEUERD_ADDR_REG_1_ | ~INSTQUEUE_REG_10__4_ | ~INSTQUEUERD_ADDR_REG_3_;
  assign new_U7656 = ~INSTQUEUERD_ADDR_REG_0_ | ~new_U3541 | ~new_U3540;
  assign new_U7657 = ~new_U3257 | ~new_U3251 | ~INSTQUEUERD_ADDR_REG_1_ | ~INSTQUEUE_REG_3__4_ | ~INSTQUEUERD_ADDR_REG_0_;
  assign new_U7658 = ~INSTQUEUERD_ADDR_REG_3_ | ~new_U3251 | ~INSTQUEUERD_ADDR_REG_1_ | ~INSTQUEUE_REG_11__4_ | ~INSTQUEUERD_ADDR_REG_0_;
  assign new_U7659 = ~new_U3257 | ~new_U3251 | ~INSTQUEUERD_ADDR_REG_1_ | ~INSTQUEUE_REG_3__5_ | ~INSTQUEUERD_ADDR_REG_0_;
  assign new_U7660 = ~INSTQUEUERD_ADDR_REG_3_ | ~new_U3517 | ~new_U3516;
  assign new_U7661 = ~new_U3252 | ~new_U3251 | ~INSTQUEUERD_ADDR_REG_0_ | ~INSTQUEUE_REG_9__6_ | ~INSTQUEUERD_ADDR_REG_3_;
  assign new_U7662 = ~INSTQUEUERD_ADDR_REG_1_ | ~new_U3523 | ~new_U3522;
  assign new_U7663 = ~new_U3253 | ~new_U3251 | ~INSTQUEUERD_ADDR_REG_1_ | ~INSTQUEUE_REG_10__6_ | ~INSTQUEUERD_ADDR_REG_3_;
  assign new_U7664 = ~INSTQUEUERD_ADDR_REG_0_ | ~new_U3251 | ~INSTQUEUERD_ADDR_REG_1_ | ~INSTQUEUE_REG_11__6_ | ~INSTQUEUERD_ADDR_REG_3_;
  assign new_U7665 = ~new_U3257 | ~new_U3253 | ~new_U3252 | ~INSTQUEUE_REG_0__6_ | ~new_U3251;
  assign new_U7666 = ~INSTQUEUERD_ADDR_REG_3_ | ~new_U3253 | ~new_U3252 | ~INSTQUEUE_REG_8__6_ | ~new_U3251;
  assign new_U7667 = ~new_U4482 | ~new_U3424;
  assign new_U7668 = ~new_U7489 | ~new_U3271;
  assign new_U7669 = ~new_U4204 | ~new_R2167_U17;
  assign new_U7670 = ~new_U4494 | ~new_U3260;
  assign new_U7671 = ~STATE2_REG_0_ | ~new_U4500;
  assign new_U7672 = ~new_U4501 | ~new_U3281;
  assign new_U7673 = ~STATE2_REG_3_ | ~new_U3282;
  assign new_U7674 = ~new_U2428 | ~new_U4502;
  assign new_U7675 = STATEBS16_REG | STATE2_REG_0_;
  assign new_U7676 = ~STATE2_REG_0_ | ~new_U7457;
  assign new_U7677 = ~STATE2_REG_0_ | ~new_U4510;
  assign new_U7678 = ~new_U3281 | ~new_U7592 | ~new_U4509;
  assign new_U7679 = ~new_R2144_U49 | ~new_U3300;
  assign new_U7680 = ~new_U4516 | ~new_U3298;
  assign new_U7681 = ~new_U3441;
  assign new_U7682 = ~INSTQUEUEWR_ADDR_REG_2_ | ~new_U3292;
  assign new_U7683 = ~new_U4521 | ~new_U3291;
  assign new_U7684 = ~new_U3442;
  assign new_U7685 = ~new_U4204 | ~new_U3260;
  assign new_U7686 = ~new_R2167_U17 | ~new_U7485;
  assign new_U7687 = ~new_U4420 | ~new_U5454;
  assign new_U7688 = ~new_U5455 | ~new_U4159;
  assign new_U7689 = ~new_U3454 | ~new_U4160;
  assign new_U7690 = ~new_U5464 | ~INSTQUEUERD_ADDR_REG_4_;
  assign new_U7691 = ~new_U4448 | ~new_U3265;
  assign new_U7692 = ~new_U4403 | ~new_U3264;
  assign new_U7693 = ~new_U3258 | ~new_U3402;
  assign new_U7694 = ~new_U4465 | ~new_U5481;
  assign new_U7695 = ~new_U7694 | ~new_U7693;
  assign new_U7696 = ~new_U5464 | ~INSTQUEUERD_ADDR_REG_3_;
  assign new_U7697 = ~new_U5497 | ~new_U4160;
  assign new_U7698 = ~INSTADDRPOINTER_REG_1_ | ~new_U4162;
  assign new_U7699 = ~new_SUB_580_U6 | ~INSTADDRPOINTER_REG_31_;
  assign new_U7700 = ~new_U3457;
  assign new_U7701 = ~INSTADDRPOINTER_REG_0_ | ~new_U4162;
  assign new_U7702 = ~INSTADDRPOINTER_REG_0_ | ~INSTADDRPOINTER_REG_31_;
  assign new_U7703 = ~new_U3458;
  assign new_U7704 = ~new_U5499 | ~new_U5489;
  assign new_U7705 = ~new_U4206 | ~new_U3388;
  assign new_U7706 = ~INSTQUEUERD_ADDR_REG_1_ | ~new_U3251;
  assign new_U7707 = ~INSTQUEUERD_ADDR_REG_2_ | ~new_U3252;
  assign new_U7708 = ~new_U3443;
  assign new_U7709 = ~new_U5464 | ~INSTQUEUERD_ADDR_REG_2_;
  assign new_U7710 = ~new_U5506 | ~new_U4160;
  assign new_U7711 = ~new_U5464 | ~INSTQUEUERD_ADDR_REG_1_;
  assign new_U7712 = ~new_U5517 | ~new_U4160;
  assign new_U7713 = ~new_U4202 | ~INSTQUEUERD_ADDR_REG_0_;
  assign new_U7714 = ~new_U5509 | ~new_U3253;
  assign new_U7715 = ~new_U5464 | ~INSTQUEUERD_ADDR_REG_0_;
  assign new_U7716 = ~new_U5523 | ~new_U4160;
  assign new_U7717 = ~new_U5525 | ~INSTQUEUEWR_ADDR_REG_3_;
  assign new_U7718 = ~new_U5533 | ~new_U3391;
  assign new_U7719 = ~new_U7681 | ~new_U4515;
  assign new_U7720 = ~new_U3441 | ~new_U3301;
  assign new_U7721 = ~new_U7720 | ~new_U7719;
  assign new_U7722 = ~new_U5525 | ~INSTQUEUEWR_ADDR_REG_2_;
  assign new_U7723 = ~new_U5537 | ~new_U3391;
  assign new_U7724 = ~new_U5525 | ~INSTQUEUEWR_ADDR_REG_1_;
  assign new_U7725 = ~new_U5542 | ~new_U3391;
  assign new_U7726 = ~new_U5525 | ~INSTQUEUEWR_ADDR_REG_0_;
  assign new_U7727 = ~new_U5545 | ~new_U3391;
  assign new_U7728 = ~new_U4465 | ~new_U3375;
  assign new_U7729 = ~new_U3258 | ~new_U3268;
  assign new_U7730 = ~new_U4159 | ~new_U3244 | ~new_U7729 | ~new_U7728;
  assign new_U7731 = ~new_U4420 | ~new_R2167_U17 | ~new_U7599;
  assign new_U7732 = ~EAX_REG_31_ | ~new_U3411;
  assign new_U7733 = ~new_U3466 | ~new_U4211;
  assign new_U7734 = ~BYTEENABLE_REG_3_ | ~new_U3420;
  assign new_U7735 = ~new_U3467 | ~new_U4208;
  assign new_U7736 = DATAWIDTH_REG_0_ | DATAWIDTH_REG_1_;
  assign new_U7737 = ~DATAWIDTH_REG_0_ | ~new_U3400;
  assign new_U7738 = ~new_U7737 | ~new_U7736;
  assign new_U7739 = ~new_U7738 | ~new_U3240;
  assign new_U7740 = ~REIP_REG_0_ | ~REIP_REG_1_;
  assign new_U7741 = ~new_U7740 | ~new_U7739;
  assign new_U7742 = ~BYTEENABLE_REG_2_ | ~new_U3420;
  assign new_U7743 = ~new_U7741 | ~new_U4208;
  assign new_U7744 = ~BYTEENABLE_REG_1_ | ~new_U3420;
  assign new_U7745 = ~new_U4208 | ~REIP_REG_1_;
  assign new_U7746 = ~BYTEENABLE_REG_0_ | ~new_U3420;
  assign new_U7747 = ~new_U4208 | ~new_U6587;
  assign new_U7748 = ~new_U4209 | ~new_U3423;
  assign new_U7749 = ~W_R_N_REG | ~new_U3236;
  assign new_U7750 = ~MORE_REG | ~new_U4165;
  assign new_U7751 = ~new_U4225 | ~new_U6588;
  assign new_U7752 = ~new_U7638 | ~STATEBS16_REG;
  assign new_U7753 = ~BS16_N | ~new_U3449;
  assign new_U7754 = ~new_U6591 | ~REQUESTPENDING_REG;
  assign new_U7755 = ~new_U6597 | ~new_U4168;
  assign new_U7756 = ~new_U4209 | ~new_U3422;
  assign new_U7757 = ~D_C_N_REG | ~new_U3236;
  assign new_U7758 = ~M_IO_N_REG | ~new_U3236;
  assign new_U7759 = ~MEMORYFETCH_REG | ~new_U4209;
  assign new_U7760 = ~new_U6602 | ~READREQUEST_REG;
  assign new_U7761 = ~new_U6603 | ~new_U4169;
  assign new_U7762 = ~new_U3475 | ~new_U4170;
  assign new_U7763 = ~new_U5461 | ~INSTQUEUERD_ADDR_REG_4_;
  assign new_U7764 = ~new_U5461 | ~INSTQUEUERD_ADDR_REG_3_;
  assign new_U7765 = ~new_U5494 | ~new_U4170;
  assign new_U7766 = ~new_U5461 | ~INSTQUEUERD_ADDR_REG_2_;
  assign new_U7767 = ~new_U5502 | ~new_U4170;
  assign new_U7768 = ~new_U5461 | ~INSTQUEUERD_ADDR_REG_1_;
  assign new_U7769 = ~new_U5513 | ~new_U4170;
  assign new_U7770 = ~new_U5461 | ~INSTQUEUERD_ADDR_REG_0_;
  assign new_U7771 = ~new_U5519 | ~new_U4170;
  assign new_U7772 = ~new_U2605 | ~new_U3264;
  assign new_U7773 = ~new_U4448 | ~new_U7483;
  assign new_U7774 = ~new_U4191 | ~new_U3288;
  assign new_U7775 = ~INSTQUEUEWR_ADDR_REG_0_ | ~new_U3284;
  assign new_U7776 = ~INSTQUEUERD_ADDR_REG_3_ | ~new_U4171;
  assign new_U7777 = ~new_U7207 | ~new_U3257;
  assign new_U7778 = ~new_U3444;
  assign new_U7779 = ~new_U3263 | ~new_U3271;
  assign new_U7780 = ~new_U7695 | ~new_U4482;
  assign new_U7781 = ~new_U3480 | ~new_U3249;
  assign new_U7782 = ~STATE2_REG_1_ | ~FLUSH_REG | ~new_U7703;
  assign new_ADD_515_U178 = ~new_ADD_515_U103 | ~new_ADD_515_U25;
  assign new_ADD_515_U177 = ~INSTADDRPOINTER_REG_12_ | ~new_ADD_515_U24;
  assign new_ADD_515_U176 = ~new_ADD_515_U104 | ~new_ADD_515_U27;
  assign new_ADD_515_U175 = ~INSTADDRPOINTER_REG_13_ | ~new_ADD_515_U26;
  assign new_ADD_515_U174 = ~new_ADD_515_U105 | ~new_ADD_515_U29;
  assign new_ADD_515_U173 = ~INSTADDRPOINTER_REG_14_ | ~new_ADD_515_U28;
  assign new_ADD_515_U172 = ~new_ADD_515_U106 | ~new_ADD_515_U31;
  assign new_ADD_515_U171 = ~INSTADDRPOINTER_REG_15_ | ~new_ADD_515_U30;
  assign new_ADD_515_U170 = ~new_ADD_515_U107 | ~new_ADD_515_U33;
  assign new_ADD_515_U169 = ~INSTADDRPOINTER_REG_16_ | ~new_ADD_515_U32;
  assign new_ADD_515_U168 = ~new_ADD_515_U108 | ~new_ADD_515_U35;
  assign new_ADD_515_U167 = ~INSTADDRPOINTER_REG_17_ | ~new_ADD_515_U34;
  assign new_ADD_515_U166 = ~new_ADD_515_U109 | ~new_ADD_515_U37;
  assign new_ADD_515_U165 = ~INSTADDRPOINTER_REG_18_ | ~new_ADD_515_U36;
  assign new_ADD_515_U164 = ~new_ADD_515_U110 | ~new_ADD_515_U39;
  assign new_ADD_515_U163 = ~INSTADDRPOINTER_REG_19_ | ~new_ADD_515_U38;
  assign new_ADD_515_U162 = ~new_ADD_515_U111 | ~new_ADD_515_U41;
  assign new_ADD_515_U161 = ~INSTADDRPOINTER_REG_20_ | ~new_ADD_515_U40;
  assign new_ADD_515_U160 = ~new_ADD_515_U112 | ~new_ADD_515_U43;
  assign new_ADD_515_U159 = ~INSTADDRPOINTER_REG_21_ | ~new_ADD_515_U42;
  assign new_ADD_515_U158 = ~new_ADD_515_U113 | ~new_ADD_515_U45;
  assign new_ADD_515_U157 = ~INSTADDRPOINTER_REG_22_ | ~new_ADD_515_U44;
  assign new_ADD_515_U156 = ~new_ADD_515_U114 | ~new_ADD_515_U47;
  assign new_ADD_515_U155 = ~INSTADDRPOINTER_REG_23_ | ~new_ADD_515_U46;
  assign new_ADD_515_U154 = ~new_ADD_515_U115 | ~new_ADD_515_U49;
  assign new_ADD_515_U153 = ~INSTADDRPOINTER_REG_24_ | ~new_ADD_515_U48;
  assign new_ADD_515_U152 = ~new_ADD_515_U116 | ~new_ADD_515_U51;
  assign new_R2027_U5 = ~INSTADDRPOINTER_REG_0_;
  assign new_R2027_U6 = ~INSTADDRPOINTER_REG_2_;
  assign new_R2027_U7 = ~INSTADDRPOINTER_REG_1_;
  assign new_R2027_U8 = ~INSTADDRPOINTER_REG_4_;
  assign new_R2027_U9 = ~INSTADDRPOINTER_REG_3_;
  assign new_R2027_U10 = ~INSTADDRPOINTER_REG_1_ | ~INSTADDRPOINTER_REG_2_ | ~INSTADDRPOINTER_REG_0_;
  assign new_R2027_U11 = ~INSTADDRPOINTER_REG_6_;
  assign new_R2027_U12 = ~INSTADDRPOINTER_REG_5_;
  assign new_R2027_U13 = ~new_R2027_U82 | ~new_R2027_U111;
  assign new_R2027_U14 = ~INSTADDRPOINTER_REG_8_;
  assign new_R2027_U15 = ~INSTADDRPOINTER_REG_7_;
  assign new_R2027_U16 = ~new_R2027_U83 | ~new_R2027_U112;
  assign new_R2027_U17 = ~new_R2027_U84 | ~new_R2027_U118;
  assign new_R2027_U18 = ~INSTADDRPOINTER_REG_9_;
  assign new_R2027_U19 = ~INSTADDRPOINTER_REG_10_;
  assign new_R2027_U20 = ~INSTADDRPOINTER_REG_12_;
  assign new_R2027_U21 = ~INSTADDRPOINTER_REG_11_;
  assign new_R2027_U22 = ~new_R2027_U85 | ~new_R2027_U120;
  assign new_R2027_U23 = ~INSTADDRPOINTER_REG_14_;
  assign new_R2027_U24 = ~INSTADDRPOINTER_REG_13_;
  assign new_R2027_U25 = ~new_R2027_U86 | ~new_R2027_U113;
  assign new_R2027_U26 = ~INSTADDRPOINTER_REG_15_;
  assign new_R2027_U27 = ~new_R2027_U87 | ~new_R2027_U119;
  assign new_R2027_U28 = ~INSTADDRPOINTER_REG_16_;
  assign new_R2027_U29 = ~INSTADDRPOINTER_REG_18_;
  assign new_R2027_U30 = ~INSTADDRPOINTER_REG_17_;
  assign new_R2027_U31 = ~new_R2027_U88 | ~new_R2027_U124;
  assign new_R2027_U32 = ~INSTADDRPOINTER_REG_20_;
  assign new_R2027_U33 = ~INSTADDRPOINTER_REG_19_;
  assign new_R2027_U34 = ~new_R2027_U89 | ~new_R2027_U117;
  assign new_R2027_U35 = ~INSTADDRPOINTER_REG_21_;
  assign new_R2027_U36 = ~new_R2027_U90 | ~new_R2027_U114;
  assign new_R2027_U37 = ~INSTADDRPOINTER_REG_22_;
  assign new_R2027_U38 = ~INSTADDRPOINTER_REG_24_;
  assign new_R2027_U39 = ~INSTADDRPOINTER_REG_23_;
  assign new_R2027_U40 = ~new_R2027_U91 | ~new_R2027_U121;
  assign new_R2027_U41 = ~INSTADDRPOINTER_REG_26_;
  assign new_R2027_U42 = ~INSTADDRPOINTER_REG_25_;
  assign new_R2027_U43 = ~new_R2027_U92 | ~new_R2027_U115;
  assign new_R2027_U44 = ~INSTADDRPOINTER_REG_27_;
  assign new_R2027_U45 = ~INSTADDRPOINTER_REG_28_;
  assign new_R2027_U46 = ~new_R2027_U93 | ~new_R2027_U116;
  assign new_R2027_U47 = ~INSTADDRPOINTER_REG_29_;
  assign new_R2027_U48 = ~new_R2027_U94 | ~new_R2027_U122;
  assign new_R2027_U49 = ~new_R2027_U123 | ~INSTADDRPOINTER_REG_29_;
  assign new_R2027_U50 = ~INSTADDRPOINTER_REG_30_;
  assign new_R2027_U51 = ~new_R2027_U142 | ~new_R2027_U141;
  assign new_R2027_U52 = ~new_R2027_U144 | ~new_R2027_U143;
  assign new_R2027_U53 = ~new_R2027_U146 | ~new_R2027_U145;
  assign new_R2027_U54 = ~new_R2027_U148 | ~new_R2027_U147;
  assign new_R2027_U55 = ~new_R2027_U150 | ~new_R2027_U149;
  assign new_R2027_U56 = ~new_R2027_U152 | ~new_R2027_U151;
  assign new_R2027_U57 = ~new_R2027_U154 | ~new_R2027_U153;
  assign new_R2027_U58 = ~new_R2027_U156 | ~new_R2027_U155;
  assign new_R2027_U59 = ~new_R2027_U158 | ~new_R2027_U157;
  assign new_R2027_U60 = ~new_R2027_U160 | ~new_R2027_U159;
  assign new_R2027_U61 = ~new_R2027_U162 | ~new_R2027_U161;
  assign new_R2027_U62 = ~new_R2027_U164 | ~new_R2027_U163;
  assign new_R2027_U63 = ~new_R2027_U166 | ~new_R2027_U165;
  assign new_R2027_U64 = ~new_R2027_U168 | ~new_R2027_U167;
  assign new_R2027_U65 = ~new_R2027_U170 | ~new_R2027_U169;
  assign new_R2027_U66 = ~new_R2027_U172 | ~new_R2027_U171;
  assign new_R2027_U67 = ~new_R2027_U174 | ~new_R2027_U173;
  assign new_R2027_U68 = ~new_R2027_U176 | ~new_R2027_U175;
  assign new_R2027_U69 = ~new_R2027_U178 | ~new_R2027_U177;
  assign new_R2027_U70 = ~new_R2027_U180 | ~new_R2027_U179;
  assign new_R2027_U71 = ~new_R2027_U182 | ~new_R2027_U181;
  assign new_R2027_U72 = ~new_R2027_U184 | ~new_R2027_U183;
  assign new_R2027_U73 = ~new_R2027_U186 | ~new_R2027_U185;
  assign new_R2027_U74 = ~new_R2027_U188 | ~new_R2027_U187;
  assign new_R2027_U75 = ~new_R2027_U190 | ~new_R2027_U189;
  assign new_R2027_U76 = ~new_R2027_U192 | ~new_R2027_U191;
  assign new_R2027_U77 = ~new_R2027_U194 | ~new_R2027_U193;
  assign new_R2027_U78 = ~new_R2027_U196 | ~new_R2027_U195;
  assign new_R2027_U79 = ~new_R2027_U198 | ~new_R2027_U197;
  assign new_R2027_U80 = ~new_R2027_U200 | ~new_R2027_U199;
  assign new_R2027_U81 = ~new_R2027_U202 | ~new_R2027_U201;
  assign new_R2027_U82 = INSTADDRPOINTER_REG_3_ & INSTADDRPOINTER_REG_4_;
  assign new_R2027_U83 = INSTADDRPOINTER_REG_5_ & INSTADDRPOINTER_REG_6_;
  assign new_R2027_U84 = INSTADDRPOINTER_REG_7_ & INSTADDRPOINTER_REG_8_;
  assign new_R2027_U85 = INSTADDRPOINTER_REG_9_ & INSTADDRPOINTER_REG_10_;
  assign new_R2027_U86 = INSTADDRPOINTER_REG_11_ & INSTADDRPOINTER_REG_12_;
  assign new_R2027_U87 = INSTADDRPOINTER_REG_13_ & INSTADDRPOINTER_REG_14_;
  assign new_R2027_U88 = INSTADDRPOINTER_REG_16_ & INSTADDRPOINTER_REG_15_;
  assign new_R2027_U89 = INSTADDRPOINTER_REG_17_ & INSTADDRPOINTER_REG_18_;
  assign new_R2027_U90 = INSTADDRPOINTER_REG_19_ & INSTADDRPOINTER_REG_20_;
  assign new_R2027_U91 = INSTADDRPOINTER_REG_22_ & INSTADDRPOINTER_REG_21_;
  assign new_R2027_U92 = INSTADDRPOINTER_REG_23_ & INSTADDRPOINTER_REG_24_;
  assign new_R2027_U93 = INSTADDRPOINTER_REG_25_ & INSTADDRPOINTER_REG_26_;
  assign new_R2027_U94 = INSTADDRPOINTER_REG_28_ & INSTADDRPOINTER_REG_27_;
  assign new_R2027_U95 = ~new_R2027_U118 | ~INSTADDRPOINTER_REG_7_;
  assign new_R2027_U96 = ~new_R2027_U112 | ~INSTADDRPOINTER_REG_5_;
  assign new_R2027_U97 = ~new_R2027_U111 | ~INSTADDRPOINTER_REG_3_;
  assign new_R2027_U98 = ~INSTADDRPOINTER_REG_31_;
  assign new_R2027_U99 = ~INSTADDRPOINTER_REG_30_ | ~new_R2027_U128;
  assign new_R2027_U100 = ~INSTADDRPOINTER_REG_1_ | ~INSTADDRPOINTER_REG_0_;
  assign new_R2027_U101 = ~new_R2027_U122 | ~INSTADDRPOINTER_REG_27_;
  assign new_R2027_U102 = ~new_R2027_U116 | ~INSTADDRPOINTER_REG_25_;
  assign new_R2027_U103 = ~new_R2027_U115 | ~INSTADDRPOINTER_REG_23_;
  assign new_R2027_U104 = ~new_R2027_U121 | ~INSTADDRPOINTER_REG_21_;
  assign new_R2027_U105 = ~new_R2027_U114 | ~INSTADDRPOINTER_REG_19_;
  assign new_R2027_U106 = ~new_R2027_U117 | ~INSTADDRPOINTER_REG_17_;
  assign new_R2027_U107 = ~new_R2027_U124 | ~INSTADDRPOINTER_REG_15_;
  assign new_R2027_U108 = ~new_R2027_U119 | ~INSTADDRPOINTER_REG_13_;
  assign new_R2027_U109 = ~new_R2027_U113 | ~INSTADDRPOINTER_REG_11_;
  assign new_R2027_U110 = ~INSTADDRPOINTER_REG_9_ | ~new_R2027_U120;
  assign new_R2027_U111 = ~new_R2027_U10;
  assign new_R2027_U112 = ~new_R2027_U13;
  assign new_R2027_U113 = ~new_R2027_U22;
  assign new_R2027_U114 = ~new_R2027_U34;
  assign new_R2027_U115 = ~new_R2027_U40;
  assign new_R2027_U116 = ~new_R2027_U43;
  assign new_R2027_U117 = ~new_R2027_U31;
  assign new_R2027_U118 = ~new_R2027_U16;
  assign new_R2027_U119 = ~new_R2027_U25;
  assign new_R2027_U120 = ~new_R2027_U17;
  assign new_R2027_U121 = ~new_R2027_U36;
  assign new_R2027_U122 = ~new_R2027_U46;
  assign new_R2027_U123 = ~new_R2027_U48;
  assign new_R2027_U124 = ~new_R2027_U27;
  assign new_R2027_U125 = ~new_R2027_U95;
  assign new_R2027_U126 = ~new_R2027_U96;
  assign new_R2027_U127 = ~new_R2027_U97;
  assign new_R2027_U128 = ~new_R2027_U49;
  assign new_R2027_U129 = ~new_R2027_U99;
  assign new_R2027_U130 = ~new_R2027_U100;
  assign new_R2027_U131 = ~new_R2027_U101;
  assign new_R2027_U132 = ~new_R2027_U102;
  assign new_R2027_U133 = ~new_R2027_U103;
  assign new_R2027_U134 = ~new_R2027_U104;
  assign new_R2027_U135 = ~new_R2027_U105;
  assign new_R2027_U136 = ~new_R2027_U106;
  assign new_R2027_U137 = ~new_R2027_U107;
  assign new_R2027_U138 = ~new_R2027_U108;
  assign new_R2027_U139 = ~new_R2027_U109;
  assign new_R2027_U140 = ~new_R2027_U110;
  assign new_R2027_U141 = ~new_R2027_U120 | ~new_R2027_U18;
  assign new_R2027_U142 = ~INSTADDRPOINTER_REG_9_ | ~new_R2027_U17;
  assign new_R2027_U143 = ~INSTADDRPOINTER_REG_8_ | ~new_R2027_U95;
  assign new_R2027_U144 = ~new_R2027_U125 | ~new_R2027_U14;
  assign new_R2027_U145 = ~new_R2027_U118 | ~new_R2027_U15;
  assign new_R2027_U146 = ~INSTADDRPOINTER_REG_7_ | ~new_R2027_U16;
  assign new_R2027_U147 = ~INSTADDRPOINTER_REG_6_ | ~new_R2027_U96;
  assign new_R2027_U148 = ~new_R2027_U126 | ~new_R2027_U11;
  assign new_R2027_U149 = ~new_R2027_U112 | ~new_R2027_U12;
  assign new_R2027_U150 = ~INSTADDRPOINTER_REG_5_ | ~new_R2027_U13;
  assign new_R2027_U151 = ~INSTADDRPOINTER_REG_4_ | ~new_R2027_U97;
  assign new_R2027_U152 = ~new_R2027_U127 | ~new_R2027_U8;
  assign new_R2027_U153 = ~new_R2027_U111 | ~new_R2027_U9;
  assign new_R2027_U154 = ~INSTADDRPOINTER_REG_3_ | ~new_R2027_U10;
  assign new_R2027_U155 = ~INSTADDRPOINTER_REG_31_ | ~new_R2027_U99;
  assign new_R2027_U156 = ~new_R2027_U129 | ~new_R2027_U98;
  assign new_R2027_U157 = ~INSTADDRPOINTER_REG_30_ | ~new_R2027_U49;
  assign new_R2027_U158 = ~new_R2027_U128 | ~new_R2027_U50;
  assign new_R2027_U159 = ~INSTADDRPOINTER_REG_2_ | ~new_R2027_U100;
  assign new_R2027_U160 = ~new_R2027_U130 | ~new_R2027_U6;
  assign new_R2027_U161 = ~new_R2027_U123 | ~new_R2027_U47;
  assign new_R2027_U162 = ~INSTADDRPOINTER_REG_29_ | ~new_R2027_U48;
  assign new_R2027_U163 = ~INSTADDRPOINTER_REG_28_ | ~new_R2027_U101;
  assign new_R2027_U164 = ~new_R2027_U131 | ~new_R2027_U45;
  assign new_R2027_U165 = ~new_R2027_U122 | ~new_R2027_U44;
  assign new_R2027_U166 = ~INSTADDRPOINTER_REG_27_ | ~new_R2027_U46;
  assign new_R2027_U167 = ~INSTADDRPOINTER_REG_26_ | ~new_R2027_U102;
  assign new_R2027_U168 = ~new_R2027_U132 | ~new_R2027_U41;
  assign new_R2027_U169 = ~new_R2027_U116 | ~new_R2027_U42;
  assign new_R2027_U170 = ~INSTADDRPOINTER_REG_25_ | ~new_R2027_U43;
  assign new_R2027_U171 = ~INSTADDRPOINTER_REG_24_ | ~new_R2027_U103;
  assign new_R2027_U172 = ~new_R2027_U133 | ~new_R2027_U38;
  assign new_R2027_U173 = ~new_R2027_U115 | ~new_R2027_U39;
  assign new_R2027_U174 = ~INSTADDRPOINTER_REG_23_ | ~new_R2027_U40;
  assign new_R2027_U175 = ~INSTADDRPOINTER_REG_22_ | ~new_R2027_U104;
  assign new_R2027_U176 = ~new_R2027_U134 | ~new_R2027_U37;
  assign new_R2027_U177 = ~new_R2027_U121 | ~new_R2027_U35;
  assign new_R2027_U178 = ~INSTADDRPOINTER_REG_21_ | ~new_R2027_U36;
  assign new_R2027_U179 = ~INSTADDRPOINTER_REG_20_ | ~new_R2027_U105;
  assign new_R2027_U180 = ~new_R2027_U135 | ~new_R2027_U32;
  assign new_R2027_U181 = ~INSTADDRPOINTER_REG_0_ | ~new_R2027_U7;
  assign new_R2027_U182 = ~INSTADDRPOINTER_REG_1_ | ~new_R2027_U5;
  assign new_R2027_U183 = ~new_R2027_U114 | ~new_R2027_U33;
  assign new_R2027_U184 = ~INSTADDRPOINTER_REG_19_ | ~new_R2027_U34;
  assign new_R2027_U185 = ~INSTADDRPOINTER_REG_18_ | ~new_R2027_U106;
  assign new_R2027_U186 = ~new_R2027_U136 | ~new_R2027_U29;
  assign new_R2027_U187 = ~new_R2027_U117 | ~new_R2027_U30;
  assign new_R2027_U188 = ~INSTADDRPOINTER_REG_17_ | ~new_R2027_U31;
  assign new_R2027_U189 = ~INSTADDRPOINTER_REG_16_ | ~new_R2027_U107;
  assign new_R2027_U190 = ~new_R2027_U137 | ~new_R2027_U28;
  assign new_R2027_U191 = ~new_R2027_U124 | ~new_R2027_U26;
  assign new_R2027_U192 = ~INSTADDRPOINTER_REG_15_ | ~new_R2027_U27;
  assign new_R2027_U193 = ~INSTADDRPOINTER_REG_14_ | ~new_R2027_U108;
  assign new_R2027_U194 = ~new_R2027_U138 | ~new_R2027_U23;
  assign new_R2027_U195 = ~new_R2027_U119 | ~new_R2027_U24;
  assign new_R2027_U196 = ~INSTADDRPOINTER_REG_13_ | ~new_R2027_U25;
  assign new_R2027_U197 = ~INSTADDRPOINTER_REG_12_ | ~new_R2027_U109;
  assign new_R2027_U198 = ~new_R2027_U139 | ~new_R2027_U20;
  assign new_R2027_U199 = ~new_R2027_U113 | ~new_R2027_U21;
  assign new_R2027_U200 = ~INSTADDRPOINTER_REG_11_ | ~new_R2027_U22;
  assign new_R2027_U201 = ~INSTADDRPOINTER_REG_10_ | ~new_R2027_U110;
  assign new_R2027_U202 = ~new_R2027_U140 | ~new_R2027_U19;
  assign new_R2278_U5 = new_R2278_U217 & new_R2278_U215;
  assign new_R2278_U6 = new_R2278_U227 & new_R2278_U225;
  assign new_R2278_U7 = new_R2278_U6 & new_R2278_U208;
  assign new_R2278_U8 = new_R2278_U7 & new_R2278_U207;
  assign new_R2278_U9 = new_R2278_U235 & new_R2278_U231;
  assign new_R2278_U10 = new_R2278_U9 & new_R2278_U206;
  assign new_R2278_U11 = new_R2278_U10 & new_R2278_U205;
  assign new_R2278_U12 = new_R2278_U11 & new_R2278_U242;
  assign new_R2278_U13 = new_R2278_U12 & new_R2278_U204;
  assign new_R2278_U14 = new_R2278_U250 & new_R2278_U246;
  assign new_R2278_U15 = new_R2278_U14 & new_R2278_U253;
  assign new_R2278_U16 = new_R2278_U15 & new_R2278_U256;
  assign new_R2278_U17 = new_R2278_U292 & new_R2278_U19;
  assign new_R2278_U18 = ~new_U2783 | ~INSTADDRPOINTER_REG_4_;
  assign new_R2278_U19 = ~new_U2787 | ~INSTADDRPOINTER_REG_0_;
  assign new_R2278_U20 = ~new_U2782 | ~INSTADDRPOINTER_REG_5_;
  assign new_R2278_U21 = ~INSTADDRPOINTER_REG_30_;
  assign new_R2278_U22 = ~new_U2770;
  assign new_R2278_U23 = ~new_U2770 | ~INSTADDRPOINTER_REG_19_;
  assign new_R2278_U24 = ~new_U2771 | ~INSTADDRPOINTER_REG_16_;
  assign new_R2278_U25 = ~new_R2278_U40 | ~new_R2278_U207;
  assign new_R2278_U26 = ~new_U2779 | ~INSTADDRPOINTER_REG_8_;
  assign new_R2278_U27 = ~new_U2778 | ~INSTADDRPOINTER_REG_9_;
  assign new_R2278_U28 = ~new_U2777 | ~INSTADDRPOINTER_REG_10_;
  assign new_R2278_U29 = ~new_U2775 | ~INSTADDRPOINTER_REG_12_;
  assign new_R2278_U30 = ~new_U2773 | ~INSTADDRPOINTER_REG_14_;
  assign new_R2278_U31 = ~new_U2774 | ~INSTADDRPOINTER_REG_13_;
  assign new_R2278_U32 = ~INSTADDRPOINTER_REG_29_;
  assign new_R2278_U33 = ~new_U2770;
  assign new_R2278_U34 = ~INSTADDRPOINTER_REG_28_;
  assign new_R2278_U35 = ~new_U2770;
  assign new_R2278_U36 = ~new_U2770 | ~INSTADDRPOINTER_REG_26_;
  assign new_R2278_U37 = ~new_R2278_U328 | ~new_R2278_U257;
  assign new_R2278_U38 = ~new_R2278_U325 | ~new_R2278_U254;
  assign new_R2278_U39 = ~new_R2278_U322 | ~new_R2278_U251;
  assign new_R2278_U40 = ~new_R2278_U306 | ~new_R2278_U229;
  assign new_R2278_U41 = ~new_R2278_U304 | ~new_R2278_U228;
  assign new_R2278_U42 = ~new_R2278_U402 | ~new_R2278_U401;
  assign new_R2278_U43 = new_R2278_U178 & new_R2278_U162;
  assign new_R2278_U44 = new_R2278_U303 & new_R2278_U179;
  assign new_R2278_U45 = new_R2278_U182 & new_R2278_U163;
  assign new_R2278_U46 = new_R2278_U302 & new_R2278_U301;
  assign new_R2278_U47 = INSTADDRPOINTER_REG_20_ & new_U2770;
  assign new_R2278_U48 = new_R2278_U178 & new_R2278_U162;
  assign new_R2278_U49 = new_R2278_U337 & new_R2278_U179;
  assign new_R2278_U50 = new_R2278_U182 & new_R2278_U301 & new_R2278_U163;
  assign new_R2278_U51 = new_R2278_U189 & new_R2278_U185;
  assign new_R2278_U52 = new_R2278_U5 & new_R2278_U51;
  assign new_R2278_U53 = new_R2278_U186 & new_R2278_U189;
  assign new_R2278_U54 = new_R2278_U295 & new_R2278_U296 & new_R2278_U293 & new_R2278_U216;
  assign new_R2278_U55 = new_R2278_U209 & new_R2278_U221 & new_R2278_U211 & new_R2278_U213;
  assign new_R2278_U56 = new_R2278_U297 & new_R2278_U298 & new_R2278_U294 & new_R2278_U210;
  assign new_R2278_U57 = new_R2278_U13 & new_R2278_U8;
  assign new_R2278_U58 = new_R2278_U332 & new_R2278_U245;
  assign new_R2278_U59 = new_R2278_U58 & new_R2278_U333 & new_R2278_U320;
  assign new_R2278_U60 = new_R2278_U16 & new_R2278_U259;
  assign new_R2278_U61 = new_R2278_U331 & new_R2278_U260;
  assign new_R2278_U62 = ~new_R2278_U364 | ~new_R2278_U363;
  assign new_R2278_U63 = ~new_R2278_U369 | ~new_R2278_U368;
  assign new_R2278_U64 = ~new_R2278_U376 | ~new_R2278_U375;
  assign new_R2278_U65 = ~new_R2278_U381 | ~new_R2278_U380;
  assign new_R2278_U66 = new_R2278_U25 & new_R2278_U23;
  assign new_R2278_U67 = new_R2278_U318 & new_R2278_U243;
  assign new_R2278_U68 = new_R2278_U315 & new_R2278_U240;
  assign new_R2278_U69 = new_R2278_U312 & new_R2278_U238;
  assign new_R2278_U70 = new_R2278_U310 & new_R2278_U236;
  assign new_R2278_U71 = new_R2278_U295 & new_R2278_U296 & new_R2278_U293 & new_R2278_U216;
  assign new_R2278_U72 = ~new_R2278_U26 | ~new_R2278_U187;
  assign new_R2278_U73 = ~new_R2278_U189 | ~new_R2278_U27;
  assign new_R2278_U74 = new_R2278_U350 & new_R2278_U349;
  assign new_R2278_U75 = ~new_R2278_U45 | ~new_R2278_U46 | ~new_R2278_U183;
  assign new_R2278_U76 = ~new_R2278_U185 | ~new_R2278_U26;
  assign new_R2278_U77 = new_R2278_U352 & new_R2278_U351;
  assign new_R2278_U78 = ~new_R2278_U197 | ~new_R2278_U165;
  assign new_R2278_U79 = ~new_R2278_U162 | ~new_R2278_U163;
  assign new_R2278_U80 = new_R2278_U354 & new_R2278_U353;
  assign new_R2278_U81 = ~new_R2278_U20 | ~new_R2278_U195;
  assign new_R2278_U82 = ~new_R2278_U165 | ~new_R2278_U164;
  assign new_R2278_U83 = new_R2278_U356 & new_R2278_U355;
  assign new_R2278_U84 = ~new_R2278_U18 | ~new_R2278_U193;
  assign new_R2278_U85 = ~new_R2278_U179 | ~new_R2278_U20;
  assign new_R2278_U86 = new_R2278_U358 & new_R2278_U357;
  assign new_R2278_U87 = ~new_R2278_U175 | ~new_R2278_U176;
  assign new_R2278_U88 = ~new_R2278_U178 | ~new_R2278_U18;
  assign new_R2278_U89 = new_R2278_U360 & new_R2278_U359;
  assign new_R2278_U90 = ~new_R2278_U172 | ~new_R2278_U173;
  assign new_R2278_U91 = ~new_R2278_U166 | ~new_R2278_U175;
  assign new_R2278_U92 = new_R2278_U362 & new_R2278_U361;
  assign new_R2278_U93 = ~new_U2769;
  assign new_R2278_U94 = ~INSTADDRPOINTER_REG_31_;
  assign new_R2278_U95 = ~new_R2278_U61 | ~new_R2278_U330;
  assign new_R2278_U96 = new_R2278_U367 & new_R2278_U366;
  assign new_R2278_U97 = ~new_R2278_U329 | ~new_R2278_U327;
  assign new_R2278_U98 = new_R2278_U372 & new_R2278_U371;
  assign new_R2278_U99 = ~new_R2278_U169 | ~new_R2278_U170;
  assign new_R2278_U100 = ~new_R2278_U167 | ~new_R2278_U172;
  assign new_R2278_U101 = new_R2278_U374 & new_R2278_U373;
  assign new_R2278_U102 = ~new_R2278_U326 | ~new_R2278_U324;
  assign new_R2278_U103 = new_R2278_U379 & new_R2278_U378;
  assign new_R2278_U104 = ~new_R2278_U323 | ~new_R2278_U321;
  assign new_R2278_U105 = new_R2278_U384 & new_R2278_U383;
  assign new_R2278_U106 = ~new_R2278_U36 | ~new_R2278_U248;
  assign new_R2278_U107 = ~new_R2278_U250 | ~new_R2278_U251;
  assign new_R2278_U108 = new_R2278_U386 & new_R2278_U385;
  assign new_R2278_U109 = ~new_R2278_U246 | ~new_R2278_U36;
  assign new_R2278_U110 = ~new_R2278_U59 | ~new_R2278_U347;
  assign new_R2278_U111 = new_R2278_U388 & new_R2278_U387;
  assign new_R2278_U112 = ~new_R2278_U67 | ~new_R2278_U316;
  assign new_R2278_U113 = ~new_R2278_U204 | ~new_R2278_U245;
  assign new_R2278_U114 = new_R2278_U390 & new_R2278_U389;
  assign new_R2278_U115 = ~new_R2278_U68 | ~new_R2278_U313;
  assign new_R2278_U116 = ~new_R2278_U243 | ~new_R2278_U242;
  assign new_R2278_U117 = new_R2278_U392 & new_R2278_U391;
  assign new_R2278_U118 = ~new_R2278_U69 | ~new_R2278_U311;
  assign new_R2278_U119 = ~new_R2278_U240 | ~new_R2278_U205;
  assign new_R2278_U120 = new_R2278_U394 & new_R2278_U393;
  assign new_R2278_U121 = ~new_R2278_U70 | ~new_R2278_U309;
  assign new_R2278_U122 = ~new_R2278_U238 | ~new_R2278_U206;
  assign new_R2278_U123 = new_R2278_U396 & new_R2278_U395;
  assign new_R2278_U124 = ~new_R2278_U232 | ~new_R2278_U233;
  assign new_R2278_U125 = ~new_R2278_U236 | ~new_R2278_U235;
  assign new_R2278_U126 = new_R2278_U398 & new_R2278_U397;
  assign new_R2278_U127 = ~new_R2278_U231 | ~new_R2278_U232;
  assign new_R2278_U128 = ~new_R2278_U66 | ~new_R2278_U345;
  assign new_R2278_U129 = new_R2278_U400 & new_R2278_U399;
  assign new_R2278_U130 = ~new_R2278_U168 | ~new_R2278_U169;
  assign new_R2278_U131 = ~new_R2278_U207 | ~new_R2278_U23;
  assign new_R2278_U132 = ~new_R2278_U307 | ~new_R2278_U343;
  assign new_R2278_U133 = new_R2278_U404 & new_R2278_U403;
  assign new_R2278_U134 = ~new_R2278_U208 | ~new_R2278_U229;
  assign new_R2278_U135 = ~new_R2278_U305 | ~new_R2278_U341;
  assign new_R2278_U136 = new_R2278_U406 & new_R2278_U405;
  assign new_R2278_U137 = ~new_R2278_U227 | ~new_R2278_U228;
  assign new_R2278_U138 = ~new_R2278_U339 | ~new_R2278_U24;
  assign new_R2278_U139 = new_R2278_U408 & new_R2278_U407;
  assign new_R2278_U140 = ~new_R2278_U223 | ~new_R2278_U56;
  assign new_R2278_U141 = ~new_R2278_U225 | ~new_R2278_U24;
  assign new_R2278_U142 = new_R2278_U410 & new_R2278_U409;
  assign new_R2278_U143 = ~new_R2278_U280 | ~new_R2278_U30;
  assign new_R2278_U144 = ~new_R2278_U209 | ~new_R2278_U210;
  assign new_R2278_U145 = new_R2278_U412 & new_R2278_U411;
  assign new_R2278_U146 = ~new_R2278_U31 | ~new_R2278_U278;
  assign new_R2278_U147 = ~new_R2278_U30 | ~new_R2278_U211;
  assign new_R2278_U148 = new_R2278_U414 & new_R2278_U413;
  assign new_R2278_U149 = ~new_R2278_U29 | ~new_R2278_U276;
  assign new_R2278_U150 = ~new_R2278_U213 | ~new_R2278_U31;
  assign new_R2278_U151 = new_R2278_U416 & new_R2278_U415;
  assign new_R2278_U152 = ~new_R2278_U219 | ~new_R2278_U71;
  assign new_R2278_U153 = ~new_R2278_U221 | ~new_R2278_U29;
  assign new_R2278_U154 = new_R2278_U418 & new_R2278_U417;
  assign new_R2278_U155 = ~new_R2278_U288 | ~new_R2278_U28;
  assign new_R2278_U156 = ~new_R2278_U215 | ~new_R2278_U216;
  assign new_R2278_U157 = new_R2278_U420 & new_R2278_U419;
  assign new_R2278_U158 = ~new_R2278_U27 | ~new_R2278_U286;
  assign new_R2278_U159 = ~new_R2278_U28 | ~new_R2278_U217;
  assign new_R2278_U160 = new_R2278_U422 & new_R2278_U421;
  assign new_R2278_U161 = ~new_R2278_U19;
  assign new_R2278_U162 = INSTADDRPOINTER_REG_7_ | new_U2780;
  assign new_R2278_U163 = ~new_U2780 | ~INSTADDRPOINTER_REG_7_;
  assign new_R2278_U164 = INSTADDRPOINTER_REG_6_ | new_U2781;
  assign new_R2278_U165 = ~new_U2781 | ~INSTADDRPOINTER_REG_6_;
  assign new_R2278_U166 = INSTADDRPOINTER_REG_3_ | new_U2784;
  assign new_R2278_U167 = INSTADDRPOINTER_REG_2_ | new_U2785;
  assign new_R2278_U168 = INSTADDRPOINTER_REG_1_ | new_U2786;
  assign new_R2278_U169 = ~new_U2786 | ~INSTADDRPOINTER_REG_1_;
  assign new_R2278_U170 = ~new_R2278_U161 | ~new_R2278_U168;
  assign new_R2278_U171 = ~new_R2278_U99;
  assign new_R2278_U172 = ~new_U2785 | ~INSTADDRPOINTER_REG_2_;
  assign new_R2278_U173 = ~new_R2278_U99 | ~new_R2278_U299;
  assign new_R2278_U174 = ~new_R2278_U90;
  assign new_R2278_U175 = ~new_U2784 | ~INSTADDRPOINTER_REG_3_;
  assign new_R2278_U176 = ~new_R2278_U300 | ~new_R2278_U166;
  assign new_R2278_U177 = ~new_R2278_U87;
  assign new_R2278_U178 = INSTADDRPOINTER_REG_4_ | new_U2783;
  assign new_R2278_U179 = INSTADDRPOINTER_REG_5_ | new_U2782;
  assign new_R2278_U180 = ~new_R2278_U20;
  assign new_R2278_U181 = ~new_R2278_U18;
  assign new_R2278_U182 = ~new_R2278_U162 | ~new_R2278_U164 | ~new_R2278_U181 | ~new_R2278_U179;
  assign new_R2278_U183 = ~new_R2278_U44 | ~new_R2278_U43 | ~new_R2278_U87;
  assign new_R2278_U184 = ~new_R2278_U75;
  assign new_R2278_U185 = INSTADDRPOINTER_REG_8_ | new_U2779;
  assign new_R2278_U186 = ~new_R2278_U26;
  assign new_R2278_U187 = ~new_R2278_U185 | ~new_R2278_U75;
  assign new_R2278_U188 = ~new_R2278_U72;
  assign new_R2278_U189 = INSTADDRPOINTER_REG_9_ | new_U2778;
  assign new_R2278_U190 = ~new_R2278_U27;
  assign new_R2278_U191 = ~new_R2278_U73;
  assign new_R2278_U192 = ~new_R2278_U76;
  assign new_R2278_U193 = ~new_R2278_U178 | ~new_R2278_U87;
  assign new_R2278_U194 = ~new_R2278_U84;
  assign new_R2278_U195 = ~new_R2278_U84 | ~new_R2278_U179;
  assign new_R2278_U196 = ~new_R2278_U81;
  assign new_R2278_U197 = ~new_R2278_U81 | ~new_R2278_U164;
  assign new_R2278_U198 = ~new_R2278_U78;
  assign new_R2278_U199 = ~new_R2278_U79;
  assign new_R2278_U200 = ~new_R2278_U82;
  assign new_R2278_U201 = ~new_R2278_U85;
  assign new_R2278_U202 = ~new_R2278_U88;
  assign new_R2278_U203 = ~new_R2278_U91;
  assign new_R2278_U204 = INSTADDRPOINTER_REG_25_ | new_U2770;
  assign new_R2278_U205 = INSTADDRPOINTER_REG_23_ | new_U2770;
  assign new_R2278_U206 = INSTADDRPOINTER_REG_22_ | new_U2770;
  assign new_R2278_U207 = INSTADDRPOINTER_REG_19_ | new_U2770;
  assign new_R2278_U208 = INSTADDRPOINTER_REG_18_ | new_U2770;
  assign new_R2278_U209 = INSTADDRPOINTER_REG_15_ | new_U2772;
  assign new_R2278_U210 = ~new_U2772 | ~INSTADDRPOINTER_REG_15_;
  assign new_R2278_U211 = INSTADDRPOINTER_REG_14_ | new_U2773;
  assign new_R2278_U212 = ~new_R2278_U30;
  assign new_R2278_U213 = INSTADDRPOINTER_REG_13_ | new_U2774;
  assign new_R2278_U214 = ~new_R2278_U31;
  assign new_R2278_U215 = INSTADDRPOINTER_REG_11_ | new_U2776;
  assign new_R2278_U216 = ~new_U2776 | ~INSTADDRPOINTER_REG_11_;
  assign new_R2278_U217 = INSTADDRPOINTER_REG_10_ | new_U2777;
  assign new_R2278_U218 = ~new_R2278_U28;
  assign new_R2278_U219 = ~new_R2278_U52 | ~new_R2278_U335;
  assign new_R2278_U220 = ~new_R2278_U152;
  assign new_R2278_U221 = INSTADDRPOINTER_REG_12_ | new_U2775;
  assign new_R2278_U222 = ~new_R2278_U29;
  assign new_R2278_U223 = ~new_R2278_U55 | ~new_R2278_U338;
  assign new_R2278_U224 = ~new_R2278_U140;
  assign new_R2278_U225 = INSTADDRPOINTER_REG_16_ | new_U2771;
  assign new_R2278_U226 = ~new_R2278_U24;
  assign new_R2278_U227 = INSTADDRPOINTER_REG_17_ | new_U2770;
  assign new_R2278_U228 = ~new_U2770 | ~INSTADDRPOINTER_REG_17_;
  assign new_R2278_U229 = ~new_U2770 | ~INSTADDRPOINTER_REG_18_;
  assign new_R2278_U230 = ~new_R2278_U23;
  assign new_R2278_U231 = INSTADDRPOINTER_REG_20_ | new_U2770;
  assign new_R2278_U232 = ~new_U2770 | ~INSTADDRPOINTER_REG_20_;
  assign new_R2278_U233 = ~new_R2278_U231 | ~new_R2278_U128;
  assign new_R2278_U234 = ~new_R2278_U124;
  assign new_R2278_U235 = INSTADDRPOINTER_REG_21_ | new_U2770;
  assign new_R2278_U236 = ~new_U2770 | ~INSTADDRPOINTER_REG_21_;
  assign new_R2278_U237 = ~new_R2278_U121;
  assign new_R2278_U238 = ~new_U2770 | ~INSTADDRPOINTER_REG_22_;
  assign new_R2278_U239 = ~new_R2278_U118;
  assign new_R2278_U240 = ~new_U2770 | ~INSTADDRPOINTER_REG_23_;
  assign new_R2278_U241 = ~new_R2278_U115;
  assign new_R2278_U242 = INSTADDRPOINTER_REG_24_ | new_U2770;
  assign new_R2278_U243 = ~new_U2770 | ~INSTADDRPOINTER_REG_24_;
  assign new_R2278_U244 = ~new_R2278_U112;
  assign new_R2278_U245 = ~new_U2770 | ~INSTADDRPOINTER_REG_25_;
  assign new_R2278_U246 = INSTADDRPOINTER_REG_26_ | new_U2770;
  assign new_R2278_U247 = ~new_R2278_U36;
  assign new_R2278_U248 = ~new_R2278_U246 | ~new_R2278_U110;
  assign new_R2278_U249 = ~new_R2278_U106;
  assign new_R2278_U250 = INSTADDRPOINTER_REG_27_ | new_U2770;
  assign new_R2278_U251 = ~new_U2770 | ~INSTADDRPOINTER_REG_27_;
  assign new_R2278_U252 = ~new_R2278_U104;
  assign new_R2278_U253 = INSTADDRPOINTER_REG_28_ | new_U2770;
  assign new_R2278_U254 = ~new_U2770 | ~INSTADDRPOINTER_REG_28_;
  assign new_R2278_U255 = ~new_R2278_U102;
  assign new_R2278_U256 = INSTADDRPOINTER_REG_29_ | new_U2770;
  assign new_R2278_U257 = ~new_U2770 | ~INSTADDRPOINTER_REG_29_;
  assign new_R2278_U258 = ~new_R2278_U97;
  assign new_R2278_U259 = INSTADDRPOINTER_REG_30_ | new_U2770;
  assign new_R2278_U260 = ~new_U2770 | ~INSTADDRPOINTER_REG_30_;
  assign new_R2278_U261 = ~new_R2278_U95;
  assign new_R2278_U262 = ~new_R2278_U100;
  assign new_R2278_U263 = ~new_R2278_U107;
  assign new_R2278_U264 = ~new_R2278_U109;
  assign new_R2278_U265 = ~new_R2278_U113;
  assign new_R2278_U266 = ~new_R2278_U116;
  assign new_R2278_U267 = ~new_R2278_U119;
  assign new_R2278_U268 = ~new_R2278_U122;
  assign new_R2278_U269 = ~new_R2278_U125;
  assign new_R2278_U270 = ~new_R2278_U127;
  assign new_R2278_U271 = ~new_R2278_U130;
  assign new_R2278_U272 = ~new_R2278_U131;
  assign new_R2278_U273 = ~new_R2278_U134;
  assign new_R2278_U274 = ~new_R2278_U137;
  assign new_R2278_U275 = ~new_R2278_U141;
  assign new_R2278_U276 = ~new_R2278_U221 | ~new_R2278_U152;
  assign new_R2278_U277 = ~new_R2278_U149;
  assign new_R2278_U278 = ~new_R2278_U149 | ~new_R2278_U213;
  assign new_R2278_U279 = ~new_R2278_U146;
  assign new_R2278_U280 = ~new_R2278_U146 | ~new_R2278_U211;
  assign new_R2278_U281 = ~new_R2278_U143;
  assign new_R2278_U282 = ~new_R2278_U144;
  assign new_R2278_U283 = ~new_R2278_U147;
  assign new_R2278_U284 = ~new_R2278_U150;
  assign new_R2278_U285 = ~new_R2278_U153;
  assign new_R2278_U286 = ~new_R2278_U189 | ~new_R2278_U72;
  assign new_R2278_U287 = ~new_R2278_U158;
  assign new_R2278_U288 = ~new_R2278_U158 | ~new_R2278_U217;
  assign new_R2278_U289 = ~new_R2278_U155;
  assign new_R2278_U290 = ~new_R2278_U156;
  assign new_R2278_U291 = ~new_R2278_U159;
  assign new_R2278_U292 = INSTADDRPOINTER_REG_0_ | new_U2787;
  assign new_R2278_U293 = ~new_R2278_U53 | ~new_R2278_U5;
  assign new_R2278_U294 = ~new_R2278_U209 | ~new_R2278_U211 | ~new_R2278_U222 | ~new_R2278_U213;
  assign new_R2278_U295 = ~new_R2278_U190 | ~new_R2278_U5;
  assign new_R2278_U296 = ~new_R2278_U218 | ~new_R2278_U5;
  assign new_R2278_U297 = ~new_R2278_U212 | ~new_R2278_U209;
  assign new_R2278_U298 = ~new_R2278_U209 | ~new_R2278_U211 | ~new_R2278_U214;
  assign new_R2278_U299 = INSTADDRPOINTER_REG_2_ | new_U2785;
  assign new_R2278_U300 = ~new_R2278_U172 | ~new_R2278_U173;
  assign new_R2278_U301 = ~new_U2781 | ~INSTADDRPOINTER_REG_6_ | ~new_R2278_U162;
  assign new_R2278_U302 = ~new_R2278_U164 | ~new_R2278_U180 | ~new_R2278_U162;
  assign new_R2278_U303 = INSTADDRPOINTER_REG_6_ | new_U2781;
  assign new_R2278_U304 = ~new_R2278_U226 | ~new_R2278_U227;
  assign new_R2278_U305 = ~new_R2278_U41;
  assign new_R2278_U306 = ~new_R2278_U41 | ~new_R2278_U208;
  assign new_R2278_U307 = ~new_R2278_U40;
  assign new_R2278_U308 = ~new_R2278_U25;
  assign new_R2278_U309 = ~new_R2278_U9 | ~new_R2278_U128;
  assign new_R2278_U310 = ~new_R2278_U47 | ~new_R2278_U235;
  assign new_R2278_U311 = ~new_R2278_U10 | ~new_R2278_U128;
  assign new_R2278_U312 = ~new_R2278_U334 | ~new_R2278_U206;
  assign new_R2278_U313 = ~new_R2278_U11 | ~new_R2278_U128;
  assign new_R2278_U314 = ~new_R2278_U312 | ~new_R2278_U238;
  assign new_R2278_U315 = ~new_R2278_U314 | ~new_R2278_U205;
  assign new_R2278_U316 = ~new_R2278_U12 | ~new_R2278_U128;
  assign new_R2278_U317 = ~new_R2278_U315 | ~new_R2278_U240;
  assign new_R2278_U318 = ~new_R2278_U317 | ~new_R2278_U242;
  assign new_R2278_U319 = ~new_R2278_U318 | ~new_R2278_U243;
  assign new_R2278_U320 = ~new_R2278_U319 | ~new_R2278_U204;
  assign new_R2278_U321 = ~new_R2278_U14 | ~new_R2278_U110;
  assign new_R2278_U322 = ~new_R2278_U247 | ~new_R2278_U250;
  assign new_R2278_U323 = ~new_R2278_U39;
  assign new_R2278_U324 = ~new_R2278_U15 | ~new_R2278_U110;
  assign new_R2278_U325 = ~new_R2278_U39 | ~new_R2278_U253;
  assign new_R2278_U326 = ~new_R2278_U38;
  assign new_R2278_U327 = ~new_R2278_U16 | ~new_R2278_U110;
  assign new_R2278_U328 = ~new_R2278_U38 | ~new_R2278_U256;
  assign new_R2278_U329 = ~new_R2278_U37;
  assign new_R2278_U330 = ~new_R2278_U60 | ~new_R2278_U110;
  assign new_R2278_U331 = ~new_R2278_U37 | ~new_R2278_U259;
  assign new_R2278_U332 = ~new_R2278_U230 | ~new_R2278_U13;
  assign new_R2278_U333 = ~new_R2278_U308 | ~new_R2278_U13;
  assign new_R2278_U334 = ~new_R2278_U310 | ~new_R2278_U236;
  assign new_R2278_U335 = ~new_R2278_U50 | ~new_R2278_U336 | ~new_R2278_U302;
  assign new_R2278_U336 = ~new_R2278_U49 | ~new_R2278_U48 | ~new_R2278_U87;
  assign new_R2278_U337 = INSTADDRPOINTER_REG_6_ | new_U2781;
  assign new_R2278_U338 = ~new_R2278_U219 | ~new_R2278_U54;
  assign new_R2278_U339 = ~new_R2278_U225 | ~new_R2278_U140;
  assign new_R2278_U340 = ~new_R2278_U138;
  assign new_R2278_U341 = ~new_R2278_U6 | ~new_R2278_U140;
  assign new_R2278_U342 = ~new_R2278_U135;
  assign new_R2278_U343 = ~new_R2278_U7 | ~new_R2278_U140;
  assign new_R2278_U344 = ~new_R2278_U132;
  assign new_R2278_U345 = ~new_R2278_U8 | ~new_R2278_U140;
  assign new_R2278_U346 = ~new_R2278_U128;
  assign new_R2278_U347 = ~new_R2278_U57 | ~new_R2278_U140;
  assign new_R2278_U348 = ~new_R2278_U110;
  assign new_R2278_U349 = ~new_R2278_U188 | ~new_R2278_U73;
  assign new_R2278_U350 = ~new_R2278_U191 | ~new_R2278_U72;
  assign new_R2278_U351 = ~new_R2278_U184 | ~new_R2278_U76;
  assign new_R2278_U352 = ~new_R2278_U192 | ~new_R2278_U75;
  assign new_R2278_U353 = ~new_R2278_U198 | ~new_R2278_U79;
  assign new_R2278_U354 = ~new_R2278_U199 | ~new_R2278_U78;
  assign new_R2278_U355 = ~new_R2278_U196 | ~new_R2278_U82;
  assign new_R2278_U356 = ~new_R2278_U200 | ~new_R2278_U81;
  assign new_R2278_U357 = ~new_R2278_U194 | ~new_R2278_U85;
  assign new_R2278_U358 = ~new_R2278_U201 | ~new_R2278_U84;
  assign new_R2278_U359 = ~new_R2278_U177 | ~new_R2278_U88;
  assign new_R2278_U360 = ~new_R2278_U202 | ~new_R2278_U87;
  assign new_R2278_U361 = ~new_R2278_U174 | ~new_R2278_U91;
  assign new_R2278_U362 = ~new_R2278_U203 | ~new_R2278_U90;
  assign new_R2278_U363 = ~new_U2769 | ~new_R2278_U94;
  assign new_R2278_U364 = ~INSTADDRPOINTER_REG_31_ | ~new_R2278_U93;
  assign new_R2278_U365 = ~new_R2278_U62;
  assign new_R2278_U366 = ~new_R2278_U261 | ~new_R2278_U365;
  assign new_R2278_U367 = ~new_R2278_U62 | ~new_R2278_U95;
  assign new_R2278_U368 = ~new_U2770 | ~new_R2278_U21;
  assign new_R2278_U369 = ~INSTADDRPOINTER_REG_30_ | ~new_R2278_U22;
  assign new_R2278_U370 = ~new_R2278_U63;
  assign new_R2278_U371 = ~new_R2278_U258 | ~new_R2278_U370;
  assign new_R2278_U372 = ~new_R2278_U63 | ~new_R2278_U97;
  assign new_R2278_U373 = ~new_R2278_U171 | ~new_R2278_U100;
  assign new_R2278_U374 = ~new_R2278_U262 | ~new_R2278_U99;
  assign new_R2278_U375 = ~new_U2770 | ~new_R2278_U32;
  assign new_R2278_U376 = ~INSTADDRPOINTER_REG_29_ | ~new_R2278_U33;
  assign new_R2278_U377 = ~new_R2278_U64;
  assign new_R2278_U378 = ~new_R2278_U255 | ~new_R2278_U377;
  assign new_R2278_U379 = ~new_R2278_U64 | ~new_R2278_U102;
  assign new_R2278_U380 = ~new_U2770 | ~new_R2278_U34;
  assign new_R2278_U381 = ~INSTADDRPOINTER_REG_28_ | ~new_R2278_U35;
  assign new_R2278_U382 = ~new_R2278_U65;
  assign new_R2278_U383 = ~new_R2278_U252 | ~new_R2278_U382;
  assign new_R2278_U384 = ~new_R2278_U65 | ~new_R2278_U104;
  assign new_R2278_U385 = ~new_R2278_U249 | ~new_R2278_U107;
  assign new_R2278_U386 = ~new_R2278_U263 | ~new_R2278_U106;
  assign new_R2278_U387 = ~new_R2278_U264 | ~new_R2278_U110;
  assign new_R2278_U388 = ~new_R2278_U348 | ~new_R2278_U109;
  assign new_R2278_U389 = ~new_R2278_U244 | ~new_R2278_U113;
  assign new_R2278_U390 = ~new_R2278_U265 | ~new_R2278_U112;
  assign new_R2278_U391 = ~new_R2278_U241 | ~new_R2278_U116;
  assign new_R2278_U392 = ~new_R2278_U266 | ~new_R2278_U115;
  assign new_R2278_U393 = ~new_R2278_U239 | ~new_R2278_U119;
  assign new_R2278_U394 = ~new_R2278_U267 | ~new_R2278_U118;
  assign new_R2278_U395 = ~new_R2278_U237 | ~new_R2278_U122;
  assign new_R2278_U396 = ~new_R2278_U268 | ~new_R2278_U121;
  assign new_R2278_U397 = ~new_R2278_U234 | ~new_R2278_U125;
  assign new_R2278_U398 = ~new_R2278_U269 | ~new_R2278_U124;
  assign new_R2278_U399 = ~new_R2278_U270 | ~new_R2278_U128;
  assign new_R2278_U400 = ~new_R2278_U346 | ~new_R2278_U127;
  assign new_R2278_U401 = ~new_R2278_U161 | ~new_R2278_U130;
  assign new_R2278_U402 = ~new_R2278_U271 | ~new_R2278_U19;
  assign new_R2278_U403 = ~new_R2278_U272 | ~new_R2278_U132;
  assign new_R2278_U404 = ~new_R2278_U344 | ~new_R2278_U131;
  assign new_R2278_U405 = ~new_R2278_U273 | ~new_R2278_U135;
  assign new_R2278_U406 = ~new_R2278_U342 | ~new_R2278_U134;
  assign new_R2278_U407 = ~new_R2278_U274 | ~new_R2278_U138;
  assign new_R2278_U408 = ~new_R2278_U340 | ~new_R2278_U137;
  assign new_R2278_U409 = ~new_R2278_U224 | ~new_R2278_U141;
  assign new_R2278_U410 = ~new_R2278_U275 | ~new_R2278_U140;
  assign new_R2278_U411 = ~new_R2278_U281 | ~new_R2278_U144;
  assign new_R2278_U412 = ~new_R2278_U282 | ~new_R2278_U143;
  assign new_R2278_U413 = ~new_R2278_U279 | ~new_R2278_U147;
  assign new_R2278_U414 = ~new_R2278_U283 | ~new_R2278_U146;
  assign new_R2278_U415 = ~new_R2278_U277 | ~new_R2278_U150;
  assign new_R2278_U416 = ~new_R2278_U284 | ~new_R2278_U149;
  assign new_R2278_U417 = ~new_R2278_U220 | ~new_R2278_U153;
  assign new_R2278_U418 = ~new_R2278_U285 | ~new_R2278_U152;
  assign new_R2278_U419 = ~new_R2278_U289 | ~new_R2278_U156;
  assign new_R2278_U420 = ~new_R2278_U290 | ~new_R2278_U155;
  assign new_R2278_U421 = ~new_R2278_U287 | ~new_R2278_U159;
  assign new_R2278_U422 = ~new_R2278_U291 | ~new_R2278_U158;
  assign new_R2358_U5 = new_R2358_U281 & new_R2358_U282 & new_R2358_U293 & new_R2358_U285;
  assign new_R2358_U6 = new_R2358_U329 & new_R2358_U325;
  assign new_R2358_U7 = new_R2358_U141 & new_R2358_U6 & new_R2358_U324;
  assign new_R2358_U8 = new_R2358_U135 & new_R2358_U5;
  assign new_R2358_U9 = new_R2358_U296 & new_R2358_U294;
  assign new_R2358_U10 = new_R2358_U304 & new_R2358_U253;
  assign new_R2358_U11 = new_R2358_U303 & new_R2358_U301;
  assign new_R2358_U12 = new_R2358_U8 & new_R2358_U7;
  assign new_R2358_U13 = new_R2358_U528 & new_R2358_U527;
  assign new_R2358_U14 = new_R2358_U379 & new_R2358_U378;
  assign new_R2358_U15 = new_R2358_U376 & new_R2358_U374;
  assign new_R2358_U16 = new_R2358_U370 & new_R2358_U367;
  assign new_R2358_U17 = new_R2358_U360 & new_R2358_U359;
  assign new_R2358_U18 = new_R2358_U354 & new_R2358_U352;
  assign new_R2358_U19 = new_R2358_U336 & new_R2358_U335;
  assign new_R2358_U20 = new_R2358_U276 & new_R2358_U274;
  assign new_R2358_U21 = new_R2358_U266 & new_R2358_U262;
  assign new_R2358_U22 = ~new_U2352;
  assign new_R2358_U23 = ~new_U2643;
  assign new_R2358_U24 = ~new_U2644;
  assign new_R2358_U25 = ~new_U2645;
  assign new_R2358_U26 = ~new_U2646;
  assign new_R2358_U27 = ~new_U2649;
  assign new_R2358_U28 = ~new_U2648;
  assign new_R2358_U29 = ~new_U2650;
  assign new_R2358_U30 = ~new_U2647;
  assign new_R2358_U31 = ~new_U2644 | ~new_R2358_U77;
  assign new_R2358_U32 = ~new_U2642;
  assign new_R2358_U33 = ~new_U2641;
  assign new_R2358_U34 = ~new_R2358_U246 | ~new_R2358_U259;
  assign new_R2358_U35 = ~new_U2620;
  assign new_R2358_U36 = ~new_U2625;
  assign new_R2358_U37 = ~new_U2624;
  assign new_R2358_U38 = ~new_U2622;
  assign new_R2358_U39 = ~new_U2623;
  assign new_R2358_U40 = ~new_U2621;
  assign new_R2358_U41 = ~new_U2626;
  assign new_R2358_U42 = ~new_U2627;
  assign new_R2358_U43 = ~new_U2628;
  assign new_R2358_U44 = ~new_U2629;
  assign new_R2358_U45 = ~new_U2630;
  assign new_R2358_U46 = ~new_U2630 | ~new_R2358_U78;
  assign new_R2358_U47 = ~new_U2639;
  assign new_R2358_U48 = ~new_U2640;
  assign new_R2358_U49 = ~new_U2642 | ~new_R2358_U490;
  assign new_R2358_U50 = ~new_U2637;
  assign new_R2358_U51 = ~new_U2637 | ~new_R2358_U80;
  assign new_R2358_U52 = ~new_U2638;
  assign new_R2358_U53 = ~new_U2638 | ~new_R2358_U531;
  assign new_R2358_U54 = ~new_U2636;
  assign new_R2358_U55 = ~new_R2358_U142 | ~new_R2358_U9;
  assign new_R2358_U56 = ~new_U2631;
  assign new_R2358_U57 = ~new_U2632;
  assign new_R2358_U58 = ~new_U2633;
  assign new_R2358_U59 = ~new_U2633 | ~new_R2358_U607;
  assign new_R2358_U60 = ~new_U2634;
  assign new_R2358_U61 = ~new_U2634 | ~new_R2358_U601;
  assign new_R2358_U62 = ~new_R2358_U438 | ~new_R2358_U320;
  assign new_R2358_U63 = ~new_R2358_U280 | ~new_R2358_U291;
  assign new_R2358_U64 = ~new_R2358_U233 | ~new_R2358_U270;
  assign new_R2358_U65 = ~new_R2358_U64 | ~new_R2358_U229;
  assign new_R2358_U66 = ~new_R2358_U417 | ~new_R2358_U316;
  assign new_R2358_U67 = ~new_R2358_U146 | ~new_R2358_U410 | ~new_R2358_U219;
  assign new_R2358_U68 = ~new_R2358_U418 | ~new_R2358_U416;
  assign new_R2358_U69 = ~new_R2358_U408 | ~new_R2358_U407 | ~new_R2358_U295;
  assign new_R2358_U70 = ~new_R2358_U313 | ~new_R2358_U67;
  assign new_R2358_U71 = ~new_U2635;
  assign new_R2358_U72 = ~new_R2358_U51 | ~new_R2358_U364;
  assign new_R2358_U73 = ~new_R2358_U414 | ~new_R2358_U305;
  assign new_R2358_U74 = ~new_R2358_U423 | ~new_R2358_U413;
  assign new_R2358_U75 = ~new_R2358_U74 | ~new_R2358_U301;
  assign new_R2358_U76 = ~new_R2358_U441 | ~new_R2358_U440;
  assign new_R2358_U77 = ~new_R2358_U454 | ~new_R2358_U453;
  assign new_R2358_U78 = ~new_R2358_U552 | ~new_R2358_U551;
  assign new_R2358_U79 = ~new_R2358_U520 | ~new_R2358_U519;
  assign new_R2358_U80 = ~new_R2358_U525 | ~new_R2358_U524;
  assign new_R2358_U81 = ~new_R2358_U533 | ~new_R2358_U532;
  assign new_R2358_U82 = ~new_R2358_U654 | ~new_R2358_U653;
  assign new_R2358_U83 = ~new_R2358_U492 | ~new_R2358_U491;
  assign new_R2358_U84 = new_R2358_U49 & new_R2358_U253;
  assign new_R2358_U85 = ~new_R2358_U494 | ~new_R2358_U493;
  assign new_R2358_U86 = ~new_R2358_U499 | ~new_R2358_U498;
  assign new_R2358_U87 = new_R2358_U246 & new_R2358_U243;
  assign new_R2358_U88 = ~new_R2358_U501 | ~new_R2358_U500;
  assign new_R2358_U89 = new_R2358_U247 & new_R2358_U244;
  assign new_R2358_U90 = ~new_R2358_U503 | ~new_R2358_U502;
  assign new_R2358_U91 = ~new_R2358_U609 | ~new_R2358_U608;
  assign new_R2358_U92 = new_R2358_U278 & new_R2358_U277;
  assign new_R2358_U93 = ~new_R2358_U611 | ~new_R2358_U610;
  assign new_R2358_U94 = new_R2358_U280 & new_R2358_U279;
  assign new_R2358_U95 = ~new_R2358_U613 | ~new_R2358_U612;
  assign new_R2358_U96 = new_R2358_U288 & new_R2358_U281;
  assign new_R2358_U97 = ~new_R2358_U615 | ~new_R2358_U614;
  assign new_R2358_U98 = new_R2358_U289 & new_R2358_U282;
  assign new_R2358_U99 = ~new_R2358_U617 | ~new_R2358_U616;
  assign new_R2358_U100 = new_R2358_U285 & new_R2358_U284;
  assign new_R2358_U101 = ~new_R2358_U619 | ~new_R2358_U618;
  assign new_R2358_U102 = new_R2358_U293 & new_R2358_U283;
  assign new_R2358_U103 = ~new_R2358_U621 | ~new_R2358_U620;
  assign new_R2358_U104 = new_R2358_U320 & new_R2358_U319;
  assign new_R2358_U105 = ~new_R2358_U623 | ~new_R2358_U622;
  assign new_R2358_U106 = new_R2358_U322 & new_R2358_U321;
  assign new_R2358_U107 = ~new_R2358_U625 | ~new_R2358_U624;
  assign new_R2358_U108 = new_R2358_U324 & new_R2358_U323;
  assign new_R2358_U109 = ~new_R2358_U627 | ~new_R2358_U626;
  assign new_R2358_U110 = ~new_R2358_U632 | ~new_R2358_U631;
  assign new_R2358_U111 = new_R2358_U233 & new_R2358_U232;
  assign new_R2358_U112 = ~new_R2358_U634 | ~new_R2358_U633;
  assign new_R2358_U113 = new_R2358_U317 & new_R2358_U316;
  assign new_R2358_U114 = ~new_R2358_U636 | ~new_R2358_U635;
  assign new_R2358_U115 = new_R2358_U295 & new_R2358_U294;
  assign new_R2358_U116 = ~new_R2358_U638 | ~new_R2358_U637;
  assign new_R2358_U117 = new_R2358_U59 & new_R2358_U296;
  assign new_R2358_U118 = ~new_R2358_U640 | ~new_R2358_U639;
  assign new_R2358_U119 = ~new_R2358_U645 | ~new_R2358_U644;
  assign new_R2358_U120 = ~new_R2358_U650 | ~new_R2358_U649;
  assign new_R2358_U121 = new_R2358_U310 & new_R2358_U53;
  assign new_R2358_U122 = ~new_R2358_U652 | ~new_R2358_U651;
  assign new_R2358_U123 = new_R2358_U235 & new_R2358_U232;
  assign new_R2358_U124 = new_R2358_U231 & new_R2358_U229;
  assign new_R2358_U125 = new_R2358_U244 & new_R2358_U243;
  assign new_R2358_U126 = new_R2358_U249 & new_R2358_U245;
  assign new_R2358_U127 = new_R2358_U245 & new_R2358_U222;
  assign new_R2358_U128 = new_R2358_U265 & new_R2358_U31;
  assign new_R2358_U129 = new_R2358_U231 & new_R2358_U230;
  assign new_R2358_U130 = new_R2358_U285 & new_R2358_U282;
  assign new_R2358_U131 = new_R2358_U288 & new_R2358_U289;
  assign new_R2358_U132 = new_R2358_U281 & new_R2358_U279;
  assign new_R2358_U133 = new_R2358_U326 & new_R2358_U323;
  assign new_R2358_U134 = new_R2358_U322 & new_R2358_U319;
  assign new_R2358_U135 = new_R2358_U279 & new_R2358_U277;
  assign new_R2358_U136 = new_R2358_U11 & new_R2358_U10;
  assign new_R2358_U137 = new_R2358_U432 & new_R2358_U425;
  assign new_R2358_U138 = new_R2358_U310 & new_R2358_U224;
  assign new_R2358_U139 = new_R2358_U415 & new_R2358_U311;
  assign new_R2358_U140 = new_R2358_U420 & new_R2358_U411;
  assign new_R2358_U141 = new_R2358_U322 & new_R2358_U319;
  assign new_R2358_U142 = new_R2358_U317 & new_R2358_U313;
  assign new_R2358_U143 = new_R2358_U12 & new_R2358_U426;
  assign new_R2358_U144 = new_R2358_U402 & new_R2358_U278;
  assign new_R2358_U145 = new_R2358_U430 & new_R2358_U144 & new_R2358_U406;
  assign new_R2358_U146 = new_R2358_U420 & new_R2358_U411;
  assign new_R2358_U147 = new_R2358_U313 & new_R2358_U317;
  assign new_R2358_U148 = new_R2358_U7 & new_R2358_U149;
  assign new_R2358_U149 = new_R2358_U9 & new_R2358_U147;
  assign new_R2358_U150 = new_R2358_U422 & new_R2358_U439;
  assign new_R2358_U151 = new_R2358_U5 & new_R2358_U279;
  assign new_R2358_U152 = new_R2358_U293 & new_R2358_U285 & new_R2358_U282;
  assign new_R2358_U153 = new_R2358_U289 & new_R2358_U287;
  assign new_R2358_U154 = new_R2358_U284 & new_R2358_U283;
  assign new_R2358_U155 = new_R2358_U156 & new_R2358_U434;
  assign new_R2358_U156 = new_R2358_U6 & new_R2358_U324;
  assign new_R2358_U157 = new_R2358_U418 & new_R2358_U46;
  assign new_R2358_U158 = new_R2358_U6 & new_R2358_U326;
  assign new_R2358_U159 = new_R2358_U313 & new_R2358_U9;
  assign new_R2358_U160 = new_R2358_U300 & new_R2358_U299 & new_R2358_U224;
  assign new_R2358_U161 = new_R2358_U369 & new_R2358_U227;
  assign new_R2358_U162 = new_R2358_U303 & new_R2358_U302;
  assign new_R2358_U163 = new_R2358_U375 & new_R2358_U307;
  assign new_R2358_U164 = ~new_U2612;
  assign new_R2358_U165 = new_R2358_U444 & new_R2358_U443;
  assign new_R2358_U166 = ~new_U2610;
  assign new_R2358_U167 = ~new_U2609;
  assign new_R2358_U168 = ~new_U2667;
  assign new_R2358_U169 = ~new_U2668;
  assign new_R2358_U170 = ~new_U2670;
  assign new_R2358_U171 = ~new_U2671;
  assign new_R2358_U172 = ~new_U2672;
  assign new_R2358_U173 = ~new_U2669;
  assign new_R2358_U174 = ~new_U2611;
  assign new_R2358_U175 = ~new_R2358_U49 | ~new_R2358_U255;
  assign new_R2358_U176 = ~new_R2358_U126 | ~new_R2358_U251 | ~new_R2358_U250;
  assign new_R2358_U177 = ~new_R2358_U247 | ~new_R2358_U257;
  assign new_R2358_U178 = ~new_R2358_U230 | ~new_R2358_U240;
  assign new_R2358_U179 = ~new_U2651;
  assign new_R2358_U180 = new_R2358_U505 & new_R2358_U504;
  assign new_R2358_U181 = ~new_U2613;
  assign new_R2358_U182 = ~new_U2614;
  assign new_R2358_U183 = ~new_U2617;
  assign new_R2358_U184 = ~new_U2615;
  assign new_R2358_U185 = ~new_U2616;
  assign new_R2358_U186 = ~new_U2618;
  assign new_R2358_U187 = ~new_U2664;
  assign new_R2358_U188 = ~new_U2665;
  assign new_R2358_U189 = ~new_U2666;
  assign new_R2358_U190 = ~new_U2663;
  assign new_R2358_U191 = ~new_U2658;
  assign new_R2358_U192 = ~new_U2659;
  assign new_R2358_U193 = ~new_U2660;
  assign new_R2358_U194 = ~new_U2661;
  assign new_R2358_U195 = ~new_U2662;
  assign new_R2358_U196 = ~new_U2654;
  assign new_R2358_U197 = ~new_U2655;
  assign new_R2358_U198 = ~new_U2656;
  assign new_R2358_U199 = ~new_U2657;
  assign new_R2358_U200 = ~new_U2652;
  assign new_R2358_U201 = ~new_U2653;
  assign new_R2358_U202 = ~new_R2358_U145 | ~new_R2358_U429;
  assign new_R2358_U203 = ~new_R2358_U292 | ~new_R2358_U332;
  assign new_R2358_U204 = ~new_R2358_U338 | ~new_R2358_U337;
  assign new_R2358_U205 = ~new_R2358_U153 | ~new_R2358_U340;
  assign new_R2358_U206 = ~new_R2358_U344 | ~new_R2358_U285;
  assign new_R2358_U207 = ~new_R2358_U283 | ~new_R2358_U342;
  assign new_R2358_U208 = ~new_R2358_U150 | ~new_R2358_U421;
  assign new_R2358_U209 = ~new_R2358_U321 | ~new_R2358_U347;
  assign new_R2358_U210 = ~new_R2358_U345 | ~new_R2358_U437;
  assign new_R2358_U211 = ~new_R2358_U350 | ~new_R2358_U325;
  assign new_R2358_U212 = ~new_R2358_U236 | ~new_R2358_U268;
  assign new_R2358_U213 = ~new_R2358_U412 | ~new_R2358_U409;
  assign new_R2358_U214 = ~new_R2358_U356 | ~new_R2358_U59;
  assign new_R2358_U215 = ~new_R2358_U61 | ~new_R2358_U70;
  assign new_R2358_U216 = ~new_R2358_U53 | ~new_R2358_U361;
  assign new_R2358_U217 = ~new_R2358_U137 | ~new_R2358_U431;
  assign new_R2358_U218 = ~new_R2358_U236 | ~new_R2358_U235;
  assign new_R2358_U219 = ~new_R2358_U139 | ~new_R2358_U138 | ~new_R2358_U217;
  assign new_R2358_U220 = ~new_R2358_U211;
  assign new_R2358_U221 = ~new_R2358_U206;
  assign new_R2358_U222 = ~new_R2358_U404 | ~new_R2358_U403;
  assign new_R2358_U223 = ~new_R2358_U51;
  assign new_R2358_U224 = ~new_R2358_U521 | ~new_R2358_U54;
  assign new_R2358_U225 = ~new_R2358_U46;
  assign new_R2358_U226 = ~new_R2358_U349 | ~new_R2358_U329;
  assign new_R2358_U227 = ~new_U2636 | ~new_R2358_U79;
  assign new_R2358_U228 = ~new_R2358_U31;
  assign new_R2358_U229 = ~new_R2358_U28 | ~new_R2358_U480 | ~new_R2358_U479;
  assign new_R2358_U230 = ~new_U2647 | ~new_R2358_U485;
  assign new_R2358_U231 = ~new_R2358_U30 | ~new_R2358_U482 | ~new_R2358_U481;
  assign new_R2358_U232 = ~new_R2358_U27 | ~new_R2358_U476 | ~new_R2358_U475;
  assign new_R2358_U233 = ~new_U2649 | ~new_R2358_U471;
  assign new_R2358_U234 = ~new_U2648 | ~new_R2358_U468;
  assign new_R2358_U235 = ~new_R2358_U29 | ~new_R2358_U478 | ~new_R2358_U477;
  assign new_R2358_U236 = ~new_U2650 | ~new_R2358_U474;
  assign new_R2358_U237 = ~new_R2358_U236 | ~new_R2358_U22;
  assign new_R2358_U238 = ~new_R2358_U123 | ~new_R2358_U237;
  assign new_R2358_U239 = ~new_R2358_U234 | ~new_R2358_U238 | ~new_R2358_U233;
  assign new_R2358_U240 = ~new_R2358_U124 | ~new_R2358_U239;
  assign new_R2358_U241 = ~new_R2358_U178;
  assign new_R2358_U242 = ~new_R2358_U23 | ~new_R2358_U452 | ~new_R2358_U451;
  assign new_R2358_U243 = ~new_R2358_U25 | ~new_R2358_U463 | ~new_R2358_U462;
  assign new_R2358_U244 = ~new_R2358_U26 | ~new_R2358_U465 | ~new_R2358_U464;
  assign new_R2358_U245 = ~new_U2643 | ~new_R2358_U450;
  assign new_R2358_U246 = ~new_U2645 | ~new_R2358_U458;
  assign new_R2358_U247 = ~new_U2646 | ~new_R2358_U461;
  assign new_R2358_U248 = ~new_R2358_U247 | ~new_R2358_U246;
  assign new_R2358_U249 = ~new_R2358_U222 | ~new_R2358_U243 | ~new_R2358_U248;
  assign new_R2358_U250 = ~new_R2358_U222 | ~new_R2358_U178 | ~new_R2358_U125;
  assign new_R2358_U251 = ~new_R2358_U228 | ~new_R2358_U242;
  assign new_R2358_U252 = ~new_R2358_U176;
  assign new_R2358_U253 = ~new_R2358_U32 | ~new_R2358_U487 | ~new_R2358_U486;
  assign new_R2358_U254 = ~new_R2358_U49;
  assign new_R2358_U255 = ~new_R2358_U253 | ~new_R2358_U176;
  assign new_R2358_U256 = ~new_R2358_U175;
  assign new_R2358_U257 = ~new_R2358_U244 | ~new_R2358_U178;
  assign new_R2358_U258 = ~new_R2358_U177;
  assign new_R2358_U259 = ~new_R2358_U177 | ~new_R2358_U243;
  assign new_R2358_U260 = ~new_R2358_U34;
  assign new_R2358_U261 = ~new_R2358_U260 | ~new_R2358_U31;
  assign new_R2358_U262 = ~new_R2358_U127 | ~new_R2358_U261;
  assign new_R2358_U263 = ~new_R2358_U455 | ~new_R2358_U24;
  assign new_R2358_U264 = ~new_R2358_U263 | ~new_R2358_U34;
  assign new_R2358_U265 = ~new_R2358_U245 | ~new_R2358_U242;
  assign new_R2358_U266 = ~new_R2358_U128 | ~new_R2358_U264;
  assign new_R2358_U267 = ~new_R2358_U455 | ~new_R2358_U24;
  assign new_R2358_U268 = ~new_U2352 | ~new_R2358_U235;
  assign new_R2358_U269 = ~new_R2358_U212;
  assign new_R2358_U270 = ~new_R2358_U212 | ~new_R2358_U232;
  assign new_R2358_U271 = ~new_R2358_U64;
  assign new_R2358_U272 = ~new_R2358_U65;
  assign new_R2358_U273 = ~new_R2358_U65 | ~new_R2358_U234;
  assign new_R2358_U274 = ~new_R2358_U129 | ~new_R2358_U273;
  assign new_R2358_U275 = ~new_R2358_U231 | ~new_R2358_U230;
  assign new_R2358_U276 = ~new_R2358_U275 | ~new_R2358_U65 | ~new_R2358_U234;
  assign new_R2358_U277 = ~new_R2358_U35 | ~new_R2358_U563 | ~new_R2358_U562;
  assign new_R2358_U278 = ~new_U2620 | ~new_R2358_U580;
  assign new_R2358_U279 = ~new_R2358_U40 | ~new_R2358_U565 | ~new_R2358_U564;
  assign new_R2358_U280 = ~new_U2621 | ~new_R2358_U595;
  assign new_R2358_U281 = ~new_R2358_U38 | ~new_R2358_U555 | ~new_R2358_U554;
  assign new_R2358_U282 = ~new_R2358_U39 | ~new_R2358_U557 | ~new_R2358_U556;
  assign new_R2358_U283 = ~new_U2625 | ~new_R2358_U583;
  assign new_R2358_U284 = ~new_U2624 | ~new_R2358_U586;
  assign new_R2358_U285 = ~new_R2358_U37 | ~new_R2358_U559 | ~new_R2358_U558;
  assign new_R2358_U286 = ~new_R2358_U284 | ~new_R2358_U283;
  assign new_R2358_U287 = ~new_R2358_U130 | ~new_R2358_U286;
  assign new_R2358_U288 = ~new_U2622 | ~new_R2358_U592;
  assign new_R2358_U289 = ~new_U2623 | ~new_R2358_U589;
  assign new_R2358_U290 = ~new_R2358_U131 | ~new_R2358_U287;
  assign new_R2358_U291 = ~new_R2358_U132 | ~new_R2358_U290;
  assign new_R2358_U292 = ~new_R2358_U63;
  assign new_R2358_U293 = ~new_R2358_U36 | ~new_R2358_U561 | ~new_R2358_U560;
  assign new_R2358_U294 = ~new_R2358_U57 | ~new_R2358_U536 | ~new_R2358_U535;
  assign new_R2358_U295 = ~new_U2632 | ~new_R2358_U604;
  assign new_R2358_U296 = ~new_R2358_U58 | ~new_R2358_U538 | ~new_R2358_U537;
  assign new_R2358_U297 = ~new_R2358_U59;
  assign new_R2358_U298 = ~new_R2358_U61;
  assign new_R2358_U299 = ~new_R2358_U13 | ~new_R2358_U71;
  assign new_R2358_U300 = ~new_U2635 | ~new_R2358_U81;
  assign new_R2358_U301 = ~new_R2358_U48 | ~new_R2358_U510 | ~new_R2358_U509;
  assign new_R2358_U302 = ~new_U2639 | ~new_R2358_U515;
  assign new_R2358_U303 = ~new_R2358_U47 | ~new_R2358_U512 | ~new_R2358_U511;
  assign new_R2358_U304 = ~new_R2358_U442 | ~new_R2358_U33;
  assign new_R2358_U305 = ~new_U2641 | ~new_R2358_U76;
  assign new_R2358_U306 = ~new_R2358_U74;
  assign new_R2358_U307 = ~new_U2640 | ~new_R2358_U518;
  assign new_R2358_U308 = ~new_R2358_U217;
  assign new_R2358_U309 = ~new_R2358_U53;
  assign new_R2358_U310 = ~new_R2358_U52 | ~new_R2358_U523 | ~new_R2358_U522;
  assign new_R2358_U311 = ~new_R2358_U526 | ~new_R2358_U50;
  assign new_R2358_U312 = ~new_R2358_U67;
  assign new_R2358_U313 = ~new_R2358_U60 | ~new_R2358_U540 | ~new_R2358_U539;
  assign new_R2358_U314 = ~new_R2358_U70;
  assign new_R2358_U315 = ~new_R2358_U213;
  assign new_R2358_U316 = ~new_U2631 | ~new_R2358_U598;
  assign new_R2358_U317 = ~new_R2358_U56 | ~new_R2358_U542 | ~new_R2358_U541;
  assign new_R2358_U318 = ~new_R2358_U68;
  assign new_R2358_U319 = ~new_R2358_U41 | ~new_R2358_U544 | ~new_R2358_U543;
  assign new_R2358_U320 = ~new_U2626 | ~new_R2358_U568;
  assign new_R2358_U321 = ~new_U2627 | ~new_R2358_U571;
  assign new_R2358_U322 = ~new_R2358_U42 | ~new_R2358_U546 | ~new_R2358_U545;
  assign new_R2358_U323 = ~new_U2628 | ~new_R2358_U574;
  assign new_R2358_U324 = ~new_R2358_U43 | ~new_R2358_U548 | ~new_R2358_U547;
  assign new_R2358_U325 = ~new_R2358_U44 | ~new_R2358_U550 | ~new_R2358_U549;
  assign new_R2358_U326 = ~new_U2629 | ~new_R2358_U577;
  assign new_R2358_U327 = ~new_R2358_U225 | ~new_R2358_U325;
  assign new_R2358_U328 = ~new_R2358_U437 | ~new_R2358_U321;
  assign new_R2358_U329 = ~new_R2358_U553 | ~new_R2358_U45;
  assign new_R2358_U330 = ~new_R2358_U202;
  assign new_R2358_U331 = ~new_R2358_U208;
  assign new_R2358_U332 = ~new_R2358_U151 | ~new_R2358_U208;
  assign new_R2358_U333 = ~new_R2358_U203;
  assign new_R2358_U334 = ~new_R2358_U234 | ~new_R2358_U229;
  assign new_R2358_U335 = ~new_R2358_U271 | ~new_R2358_U334;
  assign new_R2358_U336 = ~new_R2358_U272 | ~new_R2358_U234;
  assign new_R2358_U337 = ~new_R2358_U290 | ~new_R2358_U281;
  assign new_R2358_U338 = ~new_R2358_U5 | ~new_R2358_U208;
  assign new_R2358_U339 = ~new_R2358_U204;
  assign new_R2358_U340 = ~new_R2358_U152 | ~new_R2358_U208;
  assign new_R2358_U341 = ~new_R2358_U205;
  assign new_R2358_U342 = ~new_R2358_U208 | ~new_R2358_U293;
  assign new_R2358_U343 = ~new_R2358_U207;
  assign new_R2358_U344 = ~new_R2358_U154 | ~new_R2358_U342;
  assign new_R2358_U345 = ~new_R2358_U433 | ~new_R2358_U155;
  assign new_R2358_U346 = ~new_R2358_U210;
  assign new_R2358_U347 = ~new_R2358_U210 | ~new_R2358_U322;
  assign new_R2358_U348 = ~new_R2358_U209;
  assign new_R2358_U349 = ~new_R2358_U157 | ~new_R2358_U416;
  assign new_R2358_U350 = ~new_R2358_U326 | ~new_R2358_U226;
  assign new_R2358_U351 = ~new_R2358_U318 | ~new_R2358_U46;
  assign new_R2358_U352 = ~new_R2358_U158 | ~new_R2358_U351;
  assign new_R2358_U353 = ~new_R2358_U326 | ~new_R2358_U325;
  assign new_R2358_U354 = ~new_R2358_U226 | ~new_R2358_U353;
  assign new_R2358_U355 = ~new_R2358_U215;
  assign new_R2358_U356 = ~new_R2358_U215 | ~new_R2358_U296;
  assign new_R2358_U357 = ~new_R2358_U214;
  assign new_R2358_U358 = ~new_R2358_U313 | ~new_R2358_U61;
  assign new_R2358_U359 = ~new_R2358_U312 | ~new_R2358_U358;
  assign new_R2358_U360 = ~new_R2358_U314 | ~new_R2358_U61;
  assign new_R2358_U361 = ~new_R2358_U310 | ~new_R2358_U217;
  assign new_R2358_U362 = ~new_R2358_U216;
  assign new_R2358_U363 = ~new_R2358_U526 | ~new_R2358_U50;
  assign new_R2358_U364 = ~new_R2358_U363 | ~new_R2358_U216;
  assign new_R2358_U365 = ~new_R2358_U72;
  assign new_R2358_U366 = ~new_R2358_U365 | ~new_R2358_U227;
  assign new_R2358_U367 = ~new_R2358_U160 | ~new_R2358_U366;
  assign new_R2358_U368 = ~new_R2358_U72 | ~new_R2358_U224;
  assign new_R2358_U369 = ~new_R2358_U300 | ~new_R2358_U299;
  assign new_R2358_U370 = ~new_R2358_U161 | ~new_R2358_U368;
  assign new_R2358_U371 = ~new_R2358_U526 | ~new_R2358_U50;
  assign new_R2358_U372 = ~new_R2358_U75;
  assign new_R2358_U373 = ~new_R2358_U75 | ~new_R2358_U307;
  assign new_R2358_U374 = ~new_R2358_U162 | ~new_R2358_U373;
  assign new_R2358_U375 = ~new_R2358_U303 | ~new_R2358_U302;
  assign new_R2358_U376 = ~new_R2358_U163 | ~new_R2358_U75;
  assign new_R2358_U377 = ~new_R2358_U307 | ~new_R2358_U301;
  assign new_R2358_U378 = ~new_R2358_U306 | ~new_R2358_U377;
  assign new_R2358_U379 = ~new_R2358_U372 | ~new_R2358_U307;
  assign new_R2358_U380 = ~new_R2358_U218;
  assign new_R2358_U381 = ~new_R2358_U49 | ~new_R2358_U253;
  assign new_R2358_U382 = ~new_R2358_U267 | ~new_R2358_U31;
  assign new_R2358_U383 = ~new_R2358_U246 | ~new_R2358_U243;
  assign new_R2358_U384 = ~new_R2358_U247 | ~new_R2358_U244;
  assign new_R2358_U385 = ~new_R2358_U278 | ~new_R2358_U277;
  assign new_R2358_U386 = ~new_R2358_U280 | ~new_R2358_U279;
  assign new_R2358_U387 = ~new_R2358_U288 | ~new_R2358_U281;
  assign new_R2358_U388 = ~new_R2358_U289 | ~new_R2358_U282;
  assign new_R2358_U389 = ~new_R2358_U285 | ~new_R2358_U284;
  assign new_R2358_U390 = ~new_R2358_U293 | ~new_R2358_U283;
  assign new_R2358_U391 = ~new_R2358_U320 | ~new_R2358_U319;
  assign new_R2358_U392 = ~new_R2358_U322 | ~new_R2358_U321;
  assign new_R2358_U393 = ~new_R2358_U324 | ~new_R2358_U323;
  assign new_R2358_U394 = ~new_R2358_U329 | ~new_R2358_U46;
  assign new_R2358_U395 = ~new_R2358_U233 | ~new_R2358_U232;
  assign new_R2358_U396 = ~new_R2358_U317 | ~new_R2358_U316;
  assign new_R2358_U397 = ~new_R2358_U295 | ~new_R2358_U294;
  assign new_R2358_U398 = ~new_R2358_U59 | ~new_R2358_U296;
  assign new_R2358_U399 = ~new_R2358_U227 | ~new_R2358_U224;
  assign new_R2358_U400 = ~new_R2358_U371 | ~new_R2358_U51;
  assign new_R2358_U401 = ~new_R2358_U310 | ~new_R2358_U53;
  assign new_R2358_U402 = ~new_R2358_U63 | ~new_R2358_U277;
  assign new_R2358_U403 = ~new_R2358_U77 | ~new_R2358_U242;
  assign new_R2358_U404 = ~new_U2644 | ~new_R2358_U242;
  assign new_R2358_U405 = ~new_U2640 | ~new_R2358_U518;
  assign new_R2358_U406 = ~new_R2358_U8 | ~new_R2358_U62;
  assign new_R2358_U407 = ~new_R2358_U297 | ~new_R2358_U9;
  assign new_R2358_U408 = ~new_R2358_U298 | ~new_R2358_U9;
  assign new_R2358_U409 = ~new_R2358_U159 | ~new_R2358_U67;
  assign new_R2358_U410 = ~new_R2358_U299 | ~new_R2358_U223 | ~new_R2358_U224;
  assign new_R2358_U411 = ~new_R2358_U299 | ~new_R2358_U224 | ~new_R2358_U309 | ~new_R2358_U311;
  assign new_R2358_U412 = ~new_R2358_U69;
  assign new_R2358_U413 = ~new_R2358_U10 | ~new_R2358_U176;
  assign new_R2358_U414 = ~new_R2358_U254 | ~new_R2358_U304;
  assign new_R2358_U415 = ~new_R2358_U13 | ~new_R2358_U71;
  assign new_R2358_U416 = ~new_R2358_U426 | ~new_R2358_U67;
  assign new_R2358_U417 = ~new_R2358_U69 | ~new_R2358_U317;
  assign new_R2358_U418 = ~new_R2358_U66;
  assign new_R2358_U419 = ~new_R2358_U13 | ~new_R2358_U71;
  assign new_R2358_U420 = ~new_R2358_U428 | ~new_R2358_U427 | ~new_R2358_U419;
  assign new_R2358_U421 = ~new_R2358_U67 | ~new_R2358_U148;
  assign new_R2358_U422 = ~new_R2358_U66 | ~new_R2358_U7;
  assign new_R2358_U423 = ~new_R2358_U73;
  assign new_R2358_U424 = ~new_R2358_U405 | ~new_R2358_U302;
  assign new_R2358_U425 = ~new_R2358_U424 | ~new_R2358_U303;
  assign new_R2358_U426 = ~new_R2358_U55;
  assign new_R2358_U427 = ~new_R2358_U227 | ~new_R2358_U71;
  assign new_R2358_U428 = ~new_R2358_U534 | ~new_R2358_U227;
  assign new_R2358_U429 = ~new_R2358_U143 | ~new_R2358_U435;
  assign new_R2358_U430 = ~new_R2358_U12 | ~new_R2358_U66;
  assign new_R2358_U431 = ~new_R2358_U136 | ~new_R2358_U176;
  assign new_R2358_U432 = ~new_R2358_U11 | ~new_R2358_U73;
  assign new_R2358_U433 = ~new_R2358_U312 | ~new_R2358_U418;
  assign new_R2358_U434 = ~new_R2358_U418 | ~new_R2358_U55;
  assign new_R2358_U435 = ~new_R2358_U140 | ~new_R2358_U410 | ~new_R2358_U219;
  assign new_R2358_U436 = ~new_R2358_U133 | ~new_R2358_U327;
  assign new_R2358_U437 = ~new_R2358_U436 | ~new_R2358_U324;
  assign new_R2358_U438 = ~new_R2358_U134 | ~new_R2358_U328;
  assign new_R2358_U439 = ~new_R2358_U62;
  assign new_R2358_U440 = ~new_U2352 | ~new_R2358_U164;
  assign new_R2358_U441 = ~new_U2612 | ~new_R2358_U22;
  assign new_R2358_U442 = ~new_R2358_U76;
  assign new_R2358_U443 = ~new_R2358_U442 | ~new_U2641;
  assign new_R2358_U444 = ~new_R2358_U76 | ~new_R2358_U33;
  assign new_R2358_U445 = ~new_R2358_U442 | ~new_U2641;
  assign new_R2358_U446 = ~new_R2358_U76 | ~new_R2358_U33;
  assign new_R2358_U447 = ~new_R2358_U446 | ~new_R2358_U445;
  assign new_R2358_U448 = ~new_U2352 | ~new_R2358_U166;
  assign new_R2358_U449 = ~new_U2610 | ~new_R2358_U22;
  assign new_R2358_U450 = ~new_R2358_U449 | ~new_R2358_U448;
  assign new_R2358_U451 = ~new_U2352 | ~new_R2358_U166;
  assign new_R2358_U452 = ~new_U2610 | ~new_R2358_U22;
  assign new_R2358_U453 = ~new_U2352 | ~new_R2358_U167;
  assign new_R2358_U454 = ~new_U2609 | ~new_R2358_U22;
  assign new_R2358_U455 = ~new_R2358_U77;
  assign new_R2358_U456 = ~new_U2352 | ~new_R2358_U168;
  assign new_R2358_U457 = ~new_U2667 | ~new_R2358_U22;
  assign new_R2358_U458 = ~new_R2358_U457 | ~new_R2358_U456;
  assign new_R2358_U459 = ~new_U2352 | ~new_R2358_U169;
  assign new_R2358_U460 = ~new_U2668 | ~new_R2358_U22;
  assign new_R2358_U461 = ~new_R2358_U460 | ~new_R2358_U459;
  assign new_R2358_U462 = ~new_U2352 | ~new_R2358_U168;
  assign new_R2358_U463 = ~new_U2667 | ~new_R2358_U22;
  assign new_R2358_U464 = ~new_U2352 | ~new_R2358_U169;
  assign new_R2358_U465 = ~new_U2668 | ~new_R2358_U22;
  assign new_R2358_U466 = ~new_U2352 | ~new_R2358_U170;
  assign new_R2358_U467 = ~new_U2670 | ~new_R2358_U22;
  assign new_R2358_U468 = ~new_R2358_U467 | ~new_R2358_U466;
  assign new_R2358_U469 = ~new_U2352 | ~new_R2358_U171;
  assign new_R2358_U470 = ~new_U2671 | ~new_R2358_U22;
  assign new_R2358_U471 = ~new_R2358_U470 | ~new_R2358_U469;
  assign new_R2358_U472 = ~new_U2352 | ~new_R2358_U172;
  assign new_R2358_U473 = ~new_U2672 | ~new_R2358_U22;
  assign new_R2358_U474 = ~new_R2358_U473 | ~new_R2358_U472;
  assign new_R2358_U475 = ~new_U2352 | ~new_R2358_U171;
  assign new_R2358_U476 = ~new_U2671 | ~new_R2358_U22;
  assign new_R2358_U477 = ~new_U2352 | ~new_R2358_U172;
  assign new_R2358_U478 = ~new_U2672 | ~new_R2358_U22;
  assign new_R2358_U479 = ~new_U2352 | ~new_R2358_U170;
  assign new_R2358_U480 = ~new_U2670 | ~new_R2358_U22;
  assign new_R2358_U481 = ~new_U2352 | ~new_R2358_U173;
  assign new_R2358_U482 = ~new_U2669 | ~new_R2358_U22;
  assign new_R2358_U483 = ~new_U2352 | ~new_R2358_U173;
  assign new_R2358_U484 = ~new_U2669 | ~new_R2358_U22;
  assign new_R2358_U485 = ~new_R2358_U484 | ~new_R2358_U483;
  assign new_R2358_U486 = ~new_U2352 | ~new_R2358_U174;
  assign new_R2358_U487 = ~new_U2611 | ~new_R2358_U22;
  assign new_R2358_U488 = ~new_U2352 | ~new_R2358_U174;
  assign new_R2358_U489 = ~new_U2611 | ~new_R2358_U22;
  assign new_R2358_U490 = ~new_R2358_U489 | ~new_R2358_U488;
  assign new_R2358_U491 = ~new_R2358_U165 | ~new_R2358_U175;
  assign new_R2358_U492 = ~new_R2358_U256 | ~new_R2358_U447;
  assign new_R2358_U493 = ~new_R2358_U381 | ~new_R2358_U176;
  assign new_R2358_U494 = ~new_R2358_U84 | ~new_R2358_U252;
  assign new_R2358_U495 = ~new_R2358_U455 | ~new_U2644;
  assign new_R2358_U496 = ~new_R2358_U77 | ~new_R2358_U24;
  assign new_R2358_U497 = ~new_R2358_U496 | ~new_R2358_U495;
  assign new_R2358_U498 = ~new_R2358_U382 | ~new_R2358_U34;
  assign new_R2358_U499 = ~new_R2358_U497 | ~new_R2358_U260;
  assign new_R2358_U500 = ~new_R2358_U383 | ~new_R2358_U177;
  assign new_R2358_U501 = ~new_R2358_U87 | ~new_R2358_U258;
  assign new_R2358_U502 = ~new_R2358_U384 | ~new_R2358_U178;
  assign new_R2358_U503 = ~new_R2358_U89 | ~new_R2358_U241;
  assign new_R2358_U504 = ~new_U2352 | ~new_R2358_U179;
  assign new_R2358_U505 = ~new_U2651 | ~new_R2358_U22;
  assign new_R2358_U506 = ~new_U2352 | ~new_R2358_U179;
  assign new_R2358_U507 = ~new_U2651 | ~new_R2358_U22;
  assign new_R2358_U508 = ~new_R2358_U507 | ~new_R2358_U506;
  assign new_R2358_U509 = ~new_U2352 | ~new_R2358_U181;
  assign new_R2358_U510 = ~new_U2613 | ~new_R2358_U22;
  assign new_R2358_U511 = ~new_U2352 | ~new_R2358_U182;
  assign new_R2358_U512 = ~new_U2614 | ~new_R2358_U22;
  assign new_R2358_U513 = ~new_U2352 | ~new_R2358_U182;
  assign new_R2358_U514 = ~new_U2614 | ~new_R2358_U22;
  assign new_R2358_U515 = ~new_R2358_U514 | ~new_R2358_U513;
  assign new_R2358_U516 = ~new_U2352 | ~new_R2358_U181;
  assign new_R2358_U517 = ~new_U2613 | ~new_R2358_U22;
  assign new_R2358_U518 = ~new_R2358_U517 | ~new_R2358_U516;
  assign new_R2358_U519 = ~new_U2352 | ~new_R2358_U183;
  assign new_R2358_U520 = ~new_U2617 | ~new_R2358_U22;
  assign new_R2358_U521 = ~new_R2358_U79;
  assign new_R2358_U522 = ~new_U2352 | ~new_R2358_U184;
  assign new_R2358_U523 = ~new_U2615 | ~new_R2358_U22;
  assign new_R2358_U524 = ~new_U2352 | ~new_R2358_U185;
  assign new_R2358_U525 = ~new_U2616 | ~new_R2358_U22;
  assign new_R2358_U526 = ~new_R2358_U80;
  assign new_R2358_U527 = ~new_U2352 | ~new_R2358_U186;
  assign new_R2358_U528 = ~new_U2618 | ~new_R2358_U22;
  assign new_R2358_U529 = ~new_U2352 | ~new_R2358_U184;
  assign new_R2358_U530 = ~new_U2615 | ~new_R2358_U22;
  assign new_R2358_U531 = ~new_R2358_U530 | ~new_R2358_U529;
  assign new_R2358_U532 = ~new_U2352 | ~new_R2358_U186;
  assign new_R2358_U533 = ~new_U2618 | ~new_R2358_U22;
  assign new_R2358_U534 = ~new_R2358_U81;
  assign new_R2358_U535 = ~new_U2352 | ~new_R2358_U187;
  assign new_R2358_U536 = ~new_U2664 | ~new_R2358_U22;
  assign new_R2358_U537 = ~new_U2352 | ~new_R2358_U188;
  assign new_R2358_U538 = ~new_U2665 | ~new_R2358_U22;
  assign new_R2358_U539 = ~new_U2352 | ~new_R2358_U189;
  assign new_R2358_U540 = ~new_U2666 | ~new_R2358_U22;
  assign new_R2358_U541 = ~new_U2352 | ~new_R2358_U190;
  assign new_R2358_U542 = ~new_U2663 | ~new_R2358_U22;
  assign new_R2358_U543 = ~new_U2352 | ~new_R2358_U191;
  assign new_R2358_U544 = ~new_U2658 | ~new_R2358_U22;
  assign new_R2358_U545 = ~new_U2352 | ~new_R2358_U192;
  assign new_R2358_U546 = ~new_U2659 | ~new_R2358_U22;
  assign new_R2358_U547 = ~new_U2352 | ~new_R2358_U193;
  assign new_R2358_U548 = ~new_U2660 | ~new_R2358_U22;
  assign new_R2358_U549 = ~new_U2352 | ~new_R2358_U194;
  assign new_R2358_U550 = ~new_U2661 | ~new_R2358_U22;
  assign new_R2358_U551 = ~new_U2352 | ~new_R2358_U195;
  assign new_R2358_U552 = ~new_U2662 | ~new_R2358_U22;
  assign new_R2358_U553 = ~new_R2358_U78;
  assign new_R2358_U554 = ~new_U2352 | ~new_R2358_U196;
  assign new_R2358_U555 = ~new_U2654 | ~new_R2358_U22;
  assign new_R2358_U556 = ~new_U2352 | ~new_R2358_U197;
  assign new_R2358_U557 = ~new_U2655 | ~new_R2358_U22;
  assign new_R2358_U558 = ~new_U2352 | ~new_R2358_U198;
  assign new_R2358_U559 = ~new_U2656 | ~new_R2358_U22;
  assign new_R2358_U560 = ~new_U2352 | ~new_R2358_U199;
  assign new_R2358_U561 = ~new_U2657 | ~new_R2358_U22;
  assign new_R2358_U562 = ~new_U2352 | ~new_R2358_U200;
  assign new_R2358_U563 = ~new_U2652 | ~new_R2358_U22;
  assign new_R2358_U564 = ~new_U2352 | ~new_R2358_U201;
  assign new_R2358_U565 = ~new_U2653 | ~new_R2358_U22;
  assign new_R2358_U566 = ~new_U2352 | ~new_R2358_U191;
  assign new_R2358_U567 = ~new_U2658 | ~new_R2358_U22;
  assign new_R2358_U568 = ~new_R2358_U567 | ~new_R2358_U566;
  assign new_R2358_U569 = ~new_U2352 | ~new_R2358_U192;
  assign new_R2358_U570 = ~new_U2659 | ~new_R2358_U22;
  assign new_R2358_U571 = ~new_R2358_U570 | ~new_R2358_U569;
  assign new_R2358_U572 = ~new_U2352 | ~new_R2358_U193;
  assign new_R2358_U573 = ~new_U2660 | ~new_R2358_U22;
  assign new_R2358_U574 = ~new_R2358_U573 | ~new_R2358_U572;
  assign new_R2358_U575 = ~new_U2352 | ~new_R2358_U194;
  assign new_R2358_U576 = ~new_U2661 | ~new_R2358_U22;
  assign new_R2358_U577 = ~new_R2358_U576 | ~new_R2358_U575;
  assign new_R2358_U578 = ~new_U2352 | ~new_R2358_U200;
  assign new_R2358_U579 = ~new_U2652 | ~new_R2358_U22;
  assign new_R2358_U580 = ~new_R2358_U579 | ~new_R2358_U578;
  assign new_R2358_U581 = ~new_U2352 | ~new_R2358_U199;
  assign new_R2358_U582 = ~new_U2657 | ~new_R2358_U22;
  assign new_R2358_U583 = ~new_R2358_U582 | ~new_R2358_U581;
  assign new_R2358_U584 = ~new_U2352 | ~new_R2358_U198;
  assign new_R2358_U585 = ~new_U2656 | ~new_R2358_U22;
  assign new_R2358_U586 = ~new_R2358_U585 | ~new_R2358_U584;
  assign new_R2358_U587 = ~new_U2352 | ~new_R2358_U197;
  assign new_R2358_U588 = ~new_U2655 | ~new_R2358_U22;
  assign new_R2358_U589 = ~new_R2358_U588 | ~new_R2358_U587;
  assign new_R2358_U590 = ~new_U2352 | ~new_R2358_U196;
  assign new_R2358_U591 = ~new_U2654 | ~new_R2358_U22;
  assign new_R2358_U592 = ~new_R2358_U591 | ~new_R2358_U590;
  assign new_R2358_U593 = ~new_U2352 | ~new_R2358_U201;
  assign new_R2358_U594 = ~new_U2653 | ~new_R2358_U22;
  assign new_R2358_U595 = ~new_R2358_U594 | ~new_R2358_U593;
  assign new_R2358_U596 = ~new_U2352 | ~new_R2358_U190;
  assign new_R2358_U597 = ~new_U2663 | ~new_R2358_U22;
  assign new_R2358_U598 = ~new_R2358_U597 | ~new_R2358_U596;
  assign new_R2358_U599 = ~new_U2352 | ~new_R2358_U189;
  assign new_R2358_U600 = ~new_U2666 | ~new_R2358_U22;
  assign new_R2358_U601 = ~new_R2358_U600 | ~new_R2358_U599;
  assign new_R2358_U602 = ~new_U2352 | ~new_R2358_U187;
  assign new_R2358_U603 = ~new_U2664 | ~new_R2358_U22;
  assign new_R2358_U604 = ~new_R2358_U603 | ~new_R2358_U602;
  assign new_R2358_U605 = ~new_U2352 | ~new_R2358_U188;
  assign new_R2358_U606 = ~new_U2665 | ~new_R2358_U22;
  assign new_R2358_U607 = ~new_R2358_U606 | ~new_R2358_U605;
  assign new_R2358_U608 = ~new_R2358_U180 | ~new_R2358_U202;
  assign new_R2358_U609 = ~new_R2358_U330 | ~new_R2358_U508;
  assign new_R2358_U610 = ~new_R2358_U385 | ~new_R2358_U203;
  assign new_R2358_U611 = ~new_R2358_U92 | ~new_R2358_U333;
  assign new_R2358_U612 = ~new_R2358_U386 | ~new_R2358_U204;
  assign new_R2358_U613 = ~new_R2358_U94 | ~new_R2358_U339;
  assign new_R2358_U614 = ~new_R2358_U387 | ~new_R2358_U205;
  assign new_R2358_U615 = ~new_R2358_U96 | ~new_R2358_U341;
  assign new_R2358_U616 = ~new_R2358_U221 | ~new_R2358_U388;
  assign new_R2358_U617 = ~new_R2358_U98 | ~new_R2358_U206;
  assign new_R2358_U618 = ~new_R2358_U389 | ~new_R2358_U207;
  assign new_R2358_U619 = ~new_R2358_U100 | ~new_R2358_U343;
  assign new_R2358_U620 = ~new_R2358_U390 | ~new_R2358_U208;
  assign new_R2358_U621 = ~new_R2358_U102 | ~new_R2358_U331;
  assign new_R2358_U622 = ~new_R2358_U391 | ~new_R2358_U209;
  assign new_R2358_U623 = ~new_R2358_U104 | ~new_R2358_U348;
  assign new_R2358_U624 = ~new_R2358_U392 | ~new_R2358_U210;
  assign new_R2358_U625 = ~new_R2358_U106 | ~new_R2358_U346;
  assign new_R2358_U626 = ~new_R2358_U220 | ~new_R2358_U393;
  assign new_R2358_U627 = ~new_R2358_U108 | ~new_R2358_U211;
  assign new_R2358_U628 = ~new_R2358_U553 | ~new_U2630;
  assign new_R2358_U629 = ~new_R2358_U78 | ~new_R2358_U45;
  assign new_R2358_U630 = ~new_R2358_U629 | ~new_R2358_U628;
  assign new_R2358_U631 = ~new_R2358_U394 | ~new_R2358_U68;
  assign new_R2358_U632 = ~new_R2358_U630 | ~new_R2358_U318;
  assign new_R2358_U633 = ~new_R2358_U395 | ~new_R2358_U212;
  assign new_R2358_U634 = ~new_R2358_U111 | ~new_R2358_U269;
  assign new_R2358_U635 = ~new_R2358_U396 | ~new_R2358_U213;
  assign new_R2358_U636 = ~new_R2358_U113 | ~new_R2358_U315;
  assign new_R2358_U637 = ~new_R2358_U397 | ~new_R2358_U214;
  assign new_R2358_U638 = ~new_R2358_U115 | ~new_R2358_U357;
  assign new_R2358_U639 = ~new_R2358_U398 | ~new_R2358_U215;
  assign new_R2358_U640 = ~new_R2358_U117 | ~new_R2358_U355;
  assign new_R2358_U641 = ~new_R2358_U521 | ~new_U2636;
  assign new_R2358_U642 = ~new_R2358_U79 | ~new_R2358_U54;
  assign new_R2358_U643 = ~new_R2358_U642 | ~new_R2358_U641;
  assign new_R2358_U644 = ~new_R2358_U399 | ~new_R2358_U72;
  assign new_R2358_U645 = ~new_R2358_U643 | ~new_R2358_U365;
  assign new_R2358_U646 = ~new_R2358_U526 | ~new_U2637;
  assign new_R2358_U647 = ~new_R2358_U80 | ~new_R2358_U50;
  assign new_R2358_U648 = ~new_R2358_U647 | ~new_R2358_U646;
  assign new_R2358_U649 = ~new_R2358_U400 | ~new_R2358_U216;
  assign new_R2358_U650 = ~new_R2358_U362 | ~new_R2358_U648;
  assign new_R2358_U651 = ~new_R2358_U401 | ~new_R2358_U217;
  assign new_R2358_U652 = ~new_R2358_U121 | ~new_R2358_U308;
  assign new_R2358_U653 = ~new_U2352 | ~new_R2358_U218;
  assign new_R2358_U654 = ~new_R2358_U380 | ~new_R2358_U22;
  assign new_R2337_U5 = ~PHYADDRPOINTER_REG_1_;
  assign new_R2337_U6 = ~PHYADDRPOINTER_REG_5_;
  assign new_R2337_U7 = ~PHYADDRPOINTER_REG_4_;
  assign new_R2337_U8 = ~PHYADDRPOINTER_REG_3_;
  assign new_R2337_U9 = ~PHYADDRPOINTER_REG_2_;
  assign new_R2337_U10 = ~PHYADDRPOINTER_REG_3_ | ~PHYADDRPOINTER_REG_2_ | ~PHYADDRPOINTER_REG_4_ | ~PHYADDRPOINTER_REG_5_ | ~PHYADDRPOINTER_REG_1_;
  assign new_R2337_U11 = ~PHYADDRPOINTER_REG_7_;
  assign new_R2337_U12 = ~PHYADDRPOINTER_REG_6_;
  assign new_R2337_U13 = ~new_R2337_U81 | ~new_R2337_U108;
  assign new_R2337_U14 = ~PHYADDRPOINTER_REG_8_;
  assign new_R2337_U15 = ~PHYADDRPOINTER_REG_9_;
  assign new_R2337_U16 = ~PHYADDRPOINTER_REG_2_ | ~PHYADDRPOINTER_REG_3_ | ~PHYADDRPOINTER_REG_1_;
  assign new_R2337_U17 = ~new_R2337_U82 | ~new_R2337_U110;
  assign new_R2337_U18 = ~PHYADDRPOINTER_REG_11_;
  assign new_R2337_U19 = ~PHYADDRPOINTER_REG_10_;
  assign new_R2337_U20 = ~new_R2337_U83 | ~new_R2337_U112;
  assign new_R2337_U21 = ~PHYADDRPOINTER_REG_13_;
  assign new_R2337_U22 = ~PHYADDRPOINTER_REG_12_;
  assign new_R2337_U23 = ~new_R2337_U84 | ~new_R2337_U114;
  assign new_R2337_U24 = ~PHYADDRPOINTER_REG_15_;
  assign new_R2337_U25 = ~PHYADDRPOINTER_REG_14_;
  assign new_R2337_U26 = ~new_R2337_U85 | ~new_R2337_U116;
  assign new_R2337_U27 = ~PHYADDRPOINTER_REG_17_;
  assign new_R2337_U28 = ~PHYADDRPOINTER_REG_16_;
  assign new_R2337_U29 = ~new_R2337_U86 | ~new_R2337_U118;
  assign new_R2337_U30 = ~PHYADDRPOINTER_REG_19_;
  assign new_R2337_U31 = ~PHYADDRPOINTER_REG_18_;
  assign new_R2337_U32 = ~new_R2337_U87 | ~new_R2337_U120;
  assign new_R2337_U33 = ~PHYADDRPOINTER_REG_21_;
  assign new_R2337_U34 = ~PHYADDRPOINTER_REG_20_;
  assign new_R2337_U35 = ~new_R2337_U88 | ~new_R2337_U122;
  assign new_R2337_U36 = ~PHYADDRPOINTER_REG_23_;
  assign new_R2337_U37 = ~PHYADDRPOINTER_REG_22_;
  assign new_R2337_U38 = ~new_R2337_U89 | ~new_R2337_U124;
  assign new_R2337_U39 = ~PHYADDRPOINTER_REG_25_;
  assign new_R2337_U40 = ~PHYADDRPOINTER_REG_24_;
  assign new_R2337_U41 = ~new_R2337_U90 | ~new_R2337_U126;
  assign new_R2337_U42 = ~PHYADDRPOINTER_REG_26_;
  assign new_R2337_U43 = ~PHYADDRPOINTER_REG_26_ | ~new_R2337_U128;
  assign new_R2337_U44 = ~PHYADDRPOINTER_REG_27_;
  assign new_R2337_U45 = ~PHYADDRPOINTER_REG_27_ | ~new_R2337_U129;
  assign new_R2337_U46 = ~PHYADDRPOINTER_REG_28_;
  assign new_R2337_U47 = ~PHYADDRPOINTER_REG_28_ | ~new_R2337_U130;
  assign new_R2337_U48 = ~PHYADDRPOINTER_REG_29_;
  assign new_R2337_U49 = ~PHYADDRPOINTER_REG_29_ | ~new_R2337_U131;
  assign new_R2337_U50 = ~PHYADDRPOINTER_REG_30_;
  assign new_R2337_U51 = ~new_R2337_U135 | ~new_R2337_U134;
  assign new_R2337_U52 = ~new_R2337_U137 | ~new_R2337_U136;
  assign new_R2337_U53 = ~new_R2337_U139 | ~new_R2337_U138;
  assign new_R2337_U54 = ~new_R2337_U141 | ~new_R2337_U140;
  assign new_R2337_U55 = ~new_R2337_U143 | ~new_R2337_U142;
  assign new_R2337_U56 = ~new_R2337_U145 | ~new_R2337_U144;
  assign new_R2337_U57 = ~new_R2337_U147 | ~new_R2337_U146;
  assign new_R2337_U58 = ~new_R2337_U149 | ~new_R2337_U148;
  assign new_R2337_U59 = ~new_R2337_U151 | ~new_R2337_U150;
  assign new_R2337_U60 = ~new_R2337_U153 | ~new_R2337_U152;
  assign new_R2337_U61 = ~new_R2337_U155 | ~new_R2337_U154;
  assign new_R2337_U62 = ~new_R2337_U157 | ~new_R2337_U156;
  assign new_R2337_U63 = ~new_R2337_U159 | ~new_R2337_U158;
  assign new_R2337_U64 = ~new_R2337_U161 | ~new_R2337_U160;
  assign new_R2337_U65 = ~new_R2337_U163 | ~new_R2337_U162;
  assign new_R2337_U66 = ~new_R2337_U165 | ~new_R2337_U164;
  assign new_R2337_U67 = ~new_R2337_U167 | ~new_R2337_U166;
  assign new_R2337_U68 = ~new_R2337_U169 | ~new_R2337_U168;
  assign new_R2337_U69 = ~new_R2337_U171 | ~new_R2337_U170;
  assign new_R2337_U70 = ~new_R2337_U173 | ~new_R2337_U172;
  assign new_R2337_U71 = ~new_R2337_U175 | ~new_R2337_U174;
  assign new_R2337_U72 = ~new_R2337_U177 | ~new_R2337_U176;
  assign new_R2337_U73 = ~new_R2337_U179 | ~new_R2337_U178;
  assign new_R2337_U74 = ~new_R2337_U181 | ~new_R2337_U180;
  assign new_R2337_U75 = ~new_R2337_U183 | ~new_R2337_U182;
  assign new_R2337_U76 = ~new_R2337_U185 | ~new_R2337_U184;
  assign new_R2337_U77 = ~new_R2337_U187 | ~new_R2337_U186;
  assign new_R2337_U78 = ~new_R2337_U189 | ~new_R2337_U188;
  assign new_R2337_U79 = ~new_R2337_U191 | ~new_R2337_U190;
  assign new_R2337_U80 = ~new_R2337_U193 | ~new_R2337_U192;
  assign new_R2337_U81 = PHYADDRPOINTER_REG_7_ & PHYADDRPOINTER_REG_6_;
  assign new_R2337_U82 = PHYADDRPOINTER_REG_8_ & PHYADDRPOINTER_REG_9_;
  assign new_R2337_U83 = PHYADDRPOINTER_REG_11_ & PHYADDRPOINTER_REG_10_;
  assign new_R2337_U84 = PHYADDRPOINTER_REG_13_ & PHYADDRPOINTER_REG_12_;
  assign new_R2337_U85 = PHYADDRPOINTER_REG_15_ & PHYADDRPOINTER_REG_14_;
  assign new_R2337_U86 = PHYADDRPOINTER_REG_17_ & PHYADDRPOINTER_REG_16_;
  assign new_R2337_U87 = PHYADDRPOINTER_REG_19_ & PHYADDRPOINTER_REG_18_;
  assign new_R2337_U88 = PHYADDRPOINTER_REG_21_ & PHYADDRPOINTER_REG_20_;
  assign new_R2337_U89 = PHYADDRPOINTER_REG_23_ & PHYADDRPOINTER_REG_22_;
  assign new_R2337_U90 = PHYADDRPOINTER_REG_25_ & PHYADDRPOINTER_REG_24_;
  assign new_R2337_U91 = ~PHYADDRPOINTER_REG_8_ | ~new_R2337_U110;
  assign new_R2337_U92 = ~PHYADDRPOINTER_REG_6_ | ~new_R2337_U108;
  assign new_R2337_U93 = ~new_R2337_U106 | ~PHYADDRPOINTER_REG_4_;
  assign new_R2337_U94 = ~PHYADDRPOINTER_REG_2_ | ~PHYADDRPOINTER_REG_1_;
  assign new_R2337_U95 = ~PHYADDRPOINTER_REG_31_;
  assign new_R2337_U96 = ~PHYADDRPOINTER_REG_30_ | ~new_R2337_U132;
  assign new_R2337_U97 = ~PHYADDRPOINTER_REG_24_ | ~new_R2337_U126;
  assign new_R2337_U98 = ~PHYADDRPOINTER_REG_22_ | ~new_R2337_U124;
  assign new_R2337_U99 = ~PHYADDRPOINTER_REG_20_ | ~new_R2337_U122;
  assign new_R2337_U100 = ~PHYADDRPOINTER_REG_18_ | ~new_R2337_U120;
  assign new_R2337_U101 = ~PHYADDRPOINTER_REG_16_ | ~new_R2337_U118;
  assign new_R2337_U102 = ~PHYADDRPOINTER_REG_14_ | ~new_R2337_U116;
  assign new_R2337_U103 = ~PHYADDRPOINTER_REG_12_ | ~new_R2337_U114;
  assign new_R2337_U104 = ~PHYADDRPOINTER_REG_10_ | ~new_R2337_U112;
  assign new_R2337_U105 = ~new_R2337_U94;
  assign new_R2337_U106 = ~new_R2337_U16;
  assign new_R2337_U107 = ~new_R2337_U93;
  assign new_R2337_U108 = ~new_R2337_U10;
  assign new_R2337_U109 = ~new_R2337_U92;
  assign new_R2337_U110 = ~new_R2337_U13;
  assign new_R2337_U111 = ~new_R2337_U91;
  assign new_R2337_U112 = ~new_R2337_U17;
  assign new_R2337_U113 = ~new_R2337_U104;
  assign new_R2337_U114 = ~new_R2337_U20;
  assign new_R2337_U115 = ~new_R2337_U103;
  assign new_R2337_U116 = ~new_R2337_U23;
  assign new_R2337_U117 = ~new_R2337_U102;
  assign new_R2337_U118 = ~new_R2337_U26;
  assign new_R2337_U119 = ~new_R2337_U101;
  assign new_R2337_U120 = ~new_R2337_U29;
  assign new_R2337_U121 = ~new_R2337_U100;
  assign new_R2337_U122 = ~new_R2337_U32;
  assign new_R2337_U123 = ~new_R2337_U99;
  assign new_R2337_U124 = ~new_R2337_U35;
  assign new_R2337_U125 = ~new_R2337_U98;
  assign new_R2337_U126 = ~new_R2337_U38;
  assign new_R2337_U127 = ~new_R2337_U97;
  assign new_R2337_U128 = ~new_R2337_U41;
  assign new_R2337_U129 = ~new_R2337_U43;
  assign new_R2337_U130 = ~new_R2337_U45;
  assign new_R2337_U131 = ~new_R2337_U47;
  assign new_R2337_U132 = ~new_R2337_U49;
  assign new_R2337_U133 = ~new_R2337_U96;
  assign new_R2337_U134 = ~PHYADDRPOINTER_REG_9_ | ~new_R2337_U91;
  assign new_R2337_U135 = ~new_R2337_U111 | ~new_R2337_U15;
  assign new_R2337_U136 = ~PHYADDRPOINTER_REG_8_ | ~new_R2337_U13;
  assign new_R2337_U137 = ~new_R2337_U110 | ~new_R2337_U14;
  assign new_R2337_U138 = ~PHYADDRPOINTER_REG_7_ | ~new_R2337_U92;
  assign new_R2337_U139 = ~new_R2337_U109 | ~new_R2337_U11;
  assign new_R2337_U140 = ~PHYADDRPOINTER_REG_6_ | ~new_R2337_U10;
  assign new_R2337_U141 = ~new_R2337_U108 | ~new_R2337_U12;
  assign new_R2337_U142 = ~PHYADDRPOINTER_REG_5_ | ~new_R2337_U93;
  assign new_R2337_U143 = ~new_R2337_U107 | ~new_R2337_U6;
  assign new_R2337_U144 = ~PHYADDRPOINTER_REG_4_ | ~new_R2337_U16;
  assign new_R2337_U145 = ~new_R2337_U106 | ~new_R2337_U7;
  assign new_R2337_U146 = ~PHYADDRPOINTER_REG_3_ | ~new_R2337_U94;
  assign new_R2337_U147 = ~new_R2337_U105 | ~new_R2337_U8;
  assign new_R2337_U148 = ~PHYADDRPOINTER_REG_31_ | ~new_R2337_U96;
  assign new_R2337_U149 = ~new_R2337_U133 | ~new_R2337_U95;
  assign new_R2337_U150 = ~PHYADDRPOINTER_REG_30_ | ~new_R2337_U49;
  assign new_R2337_U151 = ~new_R2337_U132 | ~new_R2337_U50;
  assign new_R2337_U152 = ~PHYADDRPOINTER_REG_1_ | ~new_R2337_U9;
  assign new_R2337_U153 = ~PHYADDRPOINTER_REG_2_ | ~new_R2337_U5;
  assign new_R2337_U154 = ~PHYADDRPOINTER_REG_29_ | ~new_R2337_U47;
  assign new_R2337_U155 = ~new_R2337_U131 | ~new_R2337_U48;
  assign new_R2337_U156 = ~PHYADDRPOINTER_REG_28_ | ~new_R2337_U45;
  assign new_R2337_U157 = ~new_R2337_U130 | ~new_R2337_U46;
  assign new_R2337_U158 = ~PHYADDRPOINTER_REG_27_ | ~new_R2337_U43;
  assign new_R2337_U159 = ~new_R2337_U129 | ~new_R2337_U44;
  assign new_R2337_U160 = ~PHYADDRPOINTER_REG_26_ | ~new_R2337_U41;
  assign new_R2337_U161 = ~new_R2337_U128 | ~new_R2337_U42;
  assign new_R2337_U162 = ~PHYADDRPOINTER_REG_25_ | ~new_R2337_U97;
  assign new_R2337_U163 = ~new_R2337_U127 | ~new_R2337_U39;
  assign new_R2337_U164 = ~PHYADDRPOINTER_REG_24_ | ~new_R2337_U38;
  assign new_R2337_U165 = ~new_R2337_U126 | ~new_R2337_U40;
  assign new_R2337_U166 = ~PHYADDRPOINTER_REG_23_ | ~new_R2337_U98;
  assign new_R2337_U167 = ~new_R2337_U125 | ~new_R2337_U36;
  assign new_R2337_U168 = ~PHYADDRPOINTER_REG_22_ | ~new_R2337_U35;
  assign new_R2337_U169 = ~new_R2337_U124 | ~new_R2337_U37;
  assign new_R2337_U170 = ~PHYADDRPOINTER_REG_21_ | ~new_R2337_U99;
  assign new_R2337_U171 = ~new_R2337_U123 | ~new_R2337_U33;
  assign new_R2337_U172 = ~PHYADDRPOINTER_REG_20_ | ~new_R2337_U32;
  assign new_R2337_U173 = ~new_R2337_U122 | ~new_R2337_U34;
  assign new_R2337_U174 = ~PHYADDRPOINTER_REG_19_ | ~new_R2337_U100;
  assign new_R2337_U175 = ~new_R2337_U121 | ~new_R2337_U30;
  assign new_R2337_U176 = ~PHYADDRPOINTER_REG_18_ | ~new_R2337_U29;
  assign new_R2337_U177 = ~new_R2337_U120 | ~new_R2337_U31;
  assign new_R2337_U178 = ~PHYADDRPOINTER_REG_17_ | ~new_R2337_U101;
  assign new_R2337_U179 = ~new_R2337_U119 | ~new_R2337_U27;
  assign new_R2337_U180 = ~PHYADDRPOINTER_REG_16_ | ~new_R2337_U26;
  assign new_R2337_U181 = ~new_R2337_U118 | ~new_R2337_U28;
  assign new_R2337_U182 = ~PHYADDRPOINTER_REG_15_ | ~new_R2337_U102;
  assign new_R2337_U183 = ~new_R2337_U117 | ~new_R2337_U24;
  assign new_R2337_U184 = ~PHYADDRPOINTER_REG_14_ | ~new_R2337_U23;
  assign new_R2337_U185 = ~new_R2337_U116 | ~new_R2337_U25;
  assign new_R2337_U186 = ~PHYADDRPOINTER_REG_13_ | ~new_R2337_U103;
  assign new_R2337_U187 = ~new_R2337_U115 | ~new_R2337_U21;
  assign new_R2337_U188 = ~PHYADDRPOINTER_REG_12_ | ~new_R2337_U20;
  assign new_R2337_U189 = ~new_R2337_U114 | ~new_R2337_U22;
  assign new_R2337_U190 = ~PHYADDRPOINTER_REG_11_ | ~new_R2337_U104;
  assign new_R2337_U191 = ~new_R2337_U113 | ~new_R2337_U18;
  assign new_R2337_U192 = ~PHYADDRPOINTER_REG_10_ | ~new_R2337_U17;
  assign new_R2337_U193 = ~new_R2337_U112 | ~new_R2337_U19;
  assign new_R2182_U5 = new_R2182_U47 & new_U2740;
  assign new_R2182_U6 = new_R2182_U60 & new_R2182_U16;
  assign new_R2182_U7 = ~new_U2744;
  assign new_R2182_U8 = ~new_U3233;
  assign new_R2182_U9 = ~new_U3233 | ~new_U2744;
  assign new_R2182_U10 = ~new_U2742;
  assign new_R2182_U11 = ~new_U2741;
  assign new_R2182_U12 = ~new_U2740;
  assign new_R2182_U13 = ~new_R2182_U35 | ~new_R2182_U41;
  assign new_R2182_U14 = ~new_U2737;
  assign new_R2182_U15 = ~new_U2738;
  assign new_R2182_U16 = ~new_U2723 | ~new_U2739;
  assign new_R2182_U17 = ~new_U2736;
  assign new_R2182_U18 = ~new_U2735;
  assign new_R2182_U19 = ~new_R2182_U36 | ~new_R2182_U49;
  assign new_R2182_U20 = ~new_U2734;
  assign new_R2182_U21 = ~new_R2182_U37 | ~new_R2182_U46;
  assign new_R2182_U22 = ~new_R2182_U48 | ~new_U2734;
  assign new_R2182_U23 = ~new_U2733;
  assign new_R2182_U24 = ~new_R2182_U64 | ~new_R2182_U63;
  assign new_R2182_U25 = ~new_R2182_U66 | ~new_R2182_U65;
  assign new_R2182_U26 = ~new_R2182_U68 | ~new_R2182_U67;
  assign new_R2182_U27 = ~new_R2182_U72 | ~new_R2182_U71;
  assign new_R2182_U28 = ~new_R2182_U74 | ~new_R2182_U73;
  assign new_R2182_U29 = ~new_R2182_U76 | ~new_R2182_U75;
  assign new_R2182_U30 = ~new_R2182_U78 | ~new_R2182_U77;
  assign new_R2182_U31 = ~new_R2182_U80 | ~new_R2182_U79;
  assign new_R2182_U32 = ~new_R2182_U82 | ~new_R2182_U81;
  assign new_R2182_U33 = ~new_R2182_U84 | ~new_R2182_U83;
  assign new_R2182_U34 = ~new_R2182_U86 | ~new_R2182_U85;
  assign new_R2182_U35 = new_U2742 & new_U2741;
  assign new_R2182_U36 = new_U2738 & new_U2737;
  assign new_R2182_U37 = new_U2735 & new_U2736;
  assign new_R2182_U38 = ~new_U2742 | ~new_R2182_U41;
  assign new_R2182_U39 = ~new_U2732;
  assign new_R2182_U40 = ~new_U2733 | ~new_R2182_U56;
  assign new_R2182_U41 = ~new_R2182_U52 | ~new_R2182_U53;
  assign new_R2182_U42 = new_R2182_U70 & new_R2182_U69;
  assign new_R2182_U43 = ~new_R2182_U46 | ~new_U2736;
  assign new_R2182_U44 = ~new_R2182_U49 | ~new_U2738;
  assign new_R2182_U45 = ~new_R2182_U51 | ~new_R2182_U62;
  assign new_R2182_U46 = ~new_R2182_U19;
  assign new_R2182_U47 = ~new_R2182_U13;
  assign new_R2182_U48 = ~new_R2182_U21;
  assign new_R2182_U49 = ~new_R2182_U16;
  assign new_R2182_U50 = ~new_R2182_U9;
  assign new_R2182_U51 = new_U2743 | new_U2731;
  assign new_R2182_U52 = ~new_U2731 | ~new_U2743;
  assign new_R2182_U53 = ~new_R2182_U50 | ~new_R2182_U51;
  assign new_R2182_U54 = ~new_R2182_U41;
  assign new_R2182_U55 = ~new_R2182_U38;
  assign new_R2182_U56 = ~new_R2182_U22;
  assign new_R2182_U57 = ~new_R2182_U40;
  assign new_R2182_U58 = ~new_R2182_U43;
  assign new_R2182_U59 = ~new_R2182_U44;
  assign new_R2182_U60 = new_U2739 | new_U2723;
  assign new_R2182_U61 = ~new_R2182_U45;
  assign new_R2182_U62 = ~new_U2731 | ~new_U2743;
  assign new_R2182_U63 = ~new_R2182_U47 | ~new_R2182_U12;
  assign new_R2182_U64 = ~new_U2740 | ~new_R2182_U13;
  assign new_R2182_U65 = ~new_U2741 | ~new_R2182_U38;
  assign new_R2182_U66 = ~new_R2182_U55 | ~new_R2182_U11;
  assign new_R2182_U67 = ~new_U2732 | ~new_R2182_U40;
  assign new_R2182_U68 = ~new_R2182_U57 | ~new_R2182_U39;
  assign new_R2182_U69 = ~new_U2742 | ~new_R2182_U41;
  assign new_R2182_U70 = ~new_R2182_U54 | ~new_R2182_U10;
  assign new_R2182_U71 = ~new_U2733 | ~new_R2182_U22;
  assign new_R2182_U72 = ~new_R2182_U56 | ~new_R2182_U23;
  assign new_R2182_U73 = ~new_R2182_U48 | ~new_R2182_U20;
  assign new_R2182_U74 = ~new_U2734 | ~new_R2182_U21;
  assign new_R2182_U75 = ~new_U2735 | ~new_R2182_U43;
  assign new_R2182_U76 = ~new_R2182_U58 | ~new_R2182_U18;
  assign new_R2182_U77 = ~new_R2182_U46 | ~new_R2182_U17;
  assign new_R2182_U78 = ~new_U2736 | ~new_R2182_U19;
  assign new_R2182_U79 = ~new_U2737 | ~new_R2182_U44;
  assign new_R2182_U80 = ~new_R2182_U59 | ~new_R2182_U14;
  assign new_R2182_U81 = ~new_R2182_U49 | ~new_R2182_U15;
  assign new_R2182_U82 = ~new_U2738 | ~new_R2182_U16;
  assign new_R2182_U83 = ~new_R2182_U50 | ~new_R2182_U45;
  assign new_R2182_U84 = ~new_R2182_U61 | ~new_R2182_U9;
  assign new_R2182_U85 = ~new_U3233 | ~new_R2182_U7;
  assign new_R2182_U86 = ~new_U2744 | ~new_R2182_U8;
  assign new_R2144_U5 = new_R2144_U104 & new_R2144_U103;
  assign new_R2144_U6 = new_R2144_U29 & new_R2144_U27 & new_R2144_U36 & new_R2144_U35;
  assign new_R2144_U7 = new_R2144_U104 & new_R2144_U81;
  assign new_R2144_U8 = new_R2144_U138 & new_R2144_U136;
  assign new_R2144_U9 = new_R2144_U128 & new_R2144_U127;
  assign new_R2144_U10 = new_R2144_U82 & new_R2144_U213 & new_R2144_U212;
  assign new_R2144_U11 = ~new_R2144_U144 | ~new_R2144_U146;
  assign new_R2144_U12 = ~new_U2355;
  assign new_R2144_U13 = ~new_U2750;
  assign new_R2144_U14 = ~new_U2751;
  assign new_R2144_U15 = ~new_U2752;
  assign new_R2144_U16 = ~new_U2749;
  assign new_R2144_U17 = ~new_U2745;
  assign new_R2144_U18 = ~new_U2748;
  assign new_R2144_U19 = ~new_U2748 | ~new_R2144_U178;
  assign new_R2144_U20 = ~new_U2747;
  assign new_R2144_U21 = ~new_U2747 | ~new_R2144_U170;
  assign new_R2144_U22 = ~new_U2746;
  assign new_R2144_U23 = ~new_U2746 | ~new_R2144_U173;
  assign new_R2144_U24 = ~new_R2144_U79 | ~new_R2144_U63;
  assign new_R2144_U25 = ~new_R2144_U6 | ~new_R2144_U79;
  assign new_R2144_U26 = ~new_R2144_U65 | ~new_R2144_U141;
  assign new_R2144_U27 = ~new_R2144_U206 | ~new_R2144_U205;
  assign new_R2144_U28 = ~new_R2144_U186 | ~new_R2144_U185;
  assign new_R2144_U29 = ~new_R2144_U203 | ~new_R2144_U202;
  assign new_R2144_U30 = ~new_R2144_U209 | ~new_R2144_U208;
  assign new_R2144_U31 = ~new_R2144_U224 | ~new_R2144_U223;
  assign new_R2144_U32 = ~new_R2144_U221 | ~new_R2144_U220;
  assign new_R2144_U33 = ~new_R2144_U227 | ~new_R2144_U226;
  assign new_R2144_U34 = ~new_R2144_U230 | ~new_R2144_U229;
  assign new_R2144_U35 = ~new_R2144_U233 | ~new_R2144_U232;
  assign new_R2144_U36 = ~new_R2144_U236 | ~new_R2144_U235;
  assign new_R2144_U37 = ~new_R2144_U248 | ~new_R2144_U247;
  assign new_R2144_U38 = ~new_R2144_U250 | ~new_R2144_U249;
  assign new_R2144_U39 = ~new_R2144_U252 | ~new_R2144_U251;
  assign new_R2144_U40 = ~new_R2144_U254 | ~new_R2144_U253;
  assign new_R2144_U41 = ~new_R2144_U256 | ~new_R2144_U255;
  assign new_R2144_U42 = ~new_R2144_U258 | ~new_R2144_U257;
  assign new_R2144_U43 = ~new_R2144_U260 | ~new_R2144_U259;
  assign new_R2144_U44 = new_R2144_U21 & new_R2144_U105;
  assign new_R2144_U45 = ~new_R2144_U217 | ~new_R2144_U216;
  assign new_R2144_U46 = new_R2144_U19 & new_R2144_U106;
  assign new_R2144_U47 = ~new_R2144_U219 | ~new_R2144_U218;
  assign new_R2144_U48 = new_R2144_U162 & new_R2144_U109;
  assign new_R2144_U49 = ~new_R2144_U239 | ~new_R2144_U238;
  assign new_R2144_U50 = ~new_R2144_U246 | ~new_R2144_U245;
  assign new_R2144_U51 = new_R2144_U110 & new_R2144_U109;
  assign new_R2144_U52 = new_R2144_U106 & new_R2144_U105;
  assign new_R2144_U53 = new_R2144_U7 & new_R2144_U52;
  assign new_R2144_U54 = new_R2144_U152 & new_R2144_U153 & new_R2144_U103 & new_R2144_U151;
  assign new_R2144_U55 = new_R2144_U109 & new_R2144_U106;
  assign new_R2144_U56 = new_R2144_U159 & new_R2144_U19;
  assign new_R2144_U57 = new_R2144_U156 & new_R2144_U21;
  assign new_R2144_U58 = new_R2144_U159 & new_R2144_U19 & new_R2144_U21;
  assign new_R2144_U59 = new_R2144_U5 & new_R2144_U105;
  assign new_R2144_U60 = new_R2144_U126 & new_R2144_U21;
  assign new_R2144_U61 = new_R2144_U23 & new_R2144_U81;
  assign new_R2144_U62 = new_R2144_U111 & new_R2144_U110;
  assign new_R2144_U63 = new_R2144_U6 & new_R2144_U64;
  assign new_R2144_U64 = new_R2144_U32 & new_R2144_U31 & new_R2144_U34 & new_R2144_U33;
  assign new_R2144_U65 = new_R2144_U34 & new_R2144_U33;
  assign new_R2144_U66 = new_R2144_U29 & new_R2144_U36 & new_R2144_U27;
  assign new_R2144_U67 = new_R2144_U29 & new_R2144_U27;
  assign new_R2144_U68 = ~new_U2762;
  assign new_R2144_U69 = ~new_U2761;
  assign new_R2144_U70 = ~new_U2763;
  assign new_R2144_U71 = ~new_U2764;
  assign new_R2144_U72 = ~new_U2766;
  assign new_R2144_U73 = ~new_U2767;
  assign new_R2144_U74 = ~new_U2768;
  assign new_R2144_U75 = ~new_U2765;
  assign new_R2144_U76 = ~new_U2760;
  assign new_R2144_U77 = ~new_U2759;
  assign new_R2144_U78 = ~new_R2144_U29 | ~new_R2144_U79;
  assign new_R2144_U79 = ~new_R2144_U99 | ~new_R2144_U54;
  assign new_R2144_U80 = new_R2144_U211 & new_R2144_U210;
  assign new_R2144_U81 = ~new_R2144_U22 | ~new_R2144_U165 | ~new_R2144_U164;
  assign new_R2144_U82 = new_R2144_U215 & new_R2144_U214;
  assign new_R2144_U83 = ~new_R2144_U56 | ~new_R2144_U158;
  assign new_R2144_U84 = ~new_R2144_U111 | ~new_R2144_U118;
  assign new_R2144_U85 = ~new_U2754;
  assign new_R2144_U86 = ~new_U2753;
  assign new_R2144_U87 = ~new_U2755;
  assign new_R2144_U88 = ~new_U2756;
  assign new_R2144_U89 = ~new_U2757;
  assign new_R2144_U90 = ~new_U2758;
  assign new_R2144_U91 = ~new_R2144_U100 | ~new_R2144_U132;
  assign new_R2144_U92 = new_R2144_U241 & new_R2144_U240;
  assign new_R2144_U93 = ~new_R2144_U129 | ~new_R2144_U113;
  assign new_R2144_U94 = ~new_R2144_U143 | ~new_R2144_U32;
  assign new_R2144_U95 = ~new_R2144_U141 | ~new_R2144_U34;
  assign new_R2144_U96 = ~new_R2144_U79 | ~new_R2144_U66;
  assign new_R2144_U97 = ~new_R2144_U67 | ~new_R2144_U79;
  assign new_R2144_U98 = ~new_R2144_U113 | ~new_R2144_U112;
  assign new_R2144_U99 = ~new_R2144_U53 | ~new_R2144_U84;
  assign new_R2144_U100 = ~new_U2751 | ~new_R2144_U28;
  assign new_R2144_U101 = ~new_R2144_U24;
  assign new_R2144_U102 = ~new_R2144_U81;
  assign new_R2144_U103 = ~new_U2745 | ~new_R2144_U181;
  assign new_R2144_U104 = ~new_R2144_U17 | ~new_R2144_U167 | ~new_R2144_U166;
  assign new_R2144_U105 = ~new_R2144_U20 | ~new_R2144_U175 | ~new_R2144_U174;
  assign new_R2144_U106 = ~new_R2144_U18 | ~new_R2144_U201 | ~new_R2144_U200;
  assign new_R2144_U107 = ~new_R2144_U21;
  assign new_R2144_U108 = ~new_R2144_U23;
  assign new_R2144_U109 = ~new_R2144_U13 | ~new_R2144_U194 | ~new_R2144_U193;
  assign new_R2144_U110 = ~new_R2144_U16 | ~new_R2144_U196 | ~new_R2144_U195;
  assign new_R2144_U111 = ~new_U2749 | ~new_R2144_U199;
  assign new_R2144_U112 = ~new_R2144_U15 | ~new_R2144_U189 | ~new_R2144_U188;
  assign new_R2144_U113 = ~new_U2752 | ~new_R2144_U192;
  assign new_R2144_U114 = ~new_R2144_U187 | ~new_R2144_U14;
  assign new_R2144_U115 = ~new_U2355 | ~new_R2144_U112;
  assign new_R2144_U116 = ~new_U2750 | ~new_R2144_U184;
  assign new_R2144_U117 = ~new_R2144_U155 | ~new_R2144_U157;
  assign new_R2144_U118 = ~new_R2144_U51 | ~new_R2144_U117;
  assign new_R2144_U119 = ~new_R2144_U84;
  assign new_R2144_U120 = ~new_R2144_U19;
  assign new_R2144_U121 = ~new_R2144_U79;
  assign new_R2144_U122 = ~new_R2144_U78;
  assign new_R2144_U123 = ~new_R2144_U83;
  assign new_R2144_U124 = ~new_R2144_U83 | ~new_R2144_U105;
  assign new_R2144_U125 = ~new_R2144_U21 | ~new_R2144_U124;
  assign new_R2144_U126 = ~new_R2144_U23 | ~new_R2144_U81;
  assign new_R2144_U127 = ~new_R2144_U60 | ~new_R2144_U124;
  assign new_R2144_U128 = ~new_R2144_U61 | ~new_R2144_U125;
  assign new_R2144_U129 = ~new_U2355 | ~new_R2144_U112;
  assign new_R2144_U130 = ~new_R2144_U93;
  assign new_R2144_U131 = ~new_R2144_U187 | ~new_R2144_U14;
  assign new_R2144_U132 = ~new_R2144_U131 | ~new_R2144_U93;
  assign new_R2144_U133 = ~new_R2144_U91;
  assign new_R2144_U134 = ~new_R2144_U91 | ~new_R2144_U109;
  assign new_R2144_U135 = ~new_R2144_U134 | ~new_R2144_U116;
  assign new_R2144_U136 = ~new_R2144_U62 | ~new_R2144_U135;
  assign new_R2144_U137 = ~new_R2144_U161 | ~new_R2144_U110;
  assign new_R2144_U138 = ~new_R2144_U137 | ~new_R2144_U134 | ~new_R2144_U116;
  assign new_R2144_U139 = ~new_R2144_U97;
  assign new_R2144_U140 = ~new_R2144_U96;
  assign new_R2144_U141 = ~new_R2144_U25;
  assign new_R2144_U142 = ~new_R2144_U95;
  assign new_R2144_U143 = ~new_R2144_U26;
  assign new_R2144_U144 = ~new_U2355 | ~new_R2144_U24;
  assign new_R2144_U145 = ~new_R2144_U144;
  assign new_R2144_U146 = ~new_R2144_U101 | ~new_R2144_U12;
  assign new_R2144_U147 = ~new_R2144_U94;
  assign new_R2144_U148 = ~new_R2144_U98;
  assign new_R2144_U149 = ~new_R2144_U21 | ~new_R2144_U105;
  assign new_R2144_U150 = ~new_R2144_U19 | ~new_R2144_U106;
  assign new_R2144_U151 = ~new_R2144_U7 | ~new_R2144_U120 | ~new_R2144_U105;
  assign new_R2144_U152 = ~new_R2144_U107 | ~new_R2144_U7;
  assign new_R2144_U153 = ~new_R2144_U108 | ~new_R2144_U7;
  assign new_R2144_U154 = ~new_R2144_U100 | ~new_R2144_U113 | ~new_R2144_U115;
  assign new_R2144_U155 = ~new_R2144_U154 | ~new_R2144_U114;
  assign new_R2144_U156 = ~new_R2144_U104 | ~new_R2144_U103;
  assign new_R2144_U157 = ~new_U2750 | ~new_R2144_U184;
  assign new_R2144_U158 = ~new_R2144_U55 | ~new_R2144_U117 | ~new_R2144_U110;
  assign new_R2144_U159 = ~new_R2144_U199 | ~new_U2749 | ~new_R2144_U106;
  assign new_R2144_U160 = ~new_R2144_U58 | ~new_R2144_U158;
  assign new_R2144_U161 = ~new_U2749 | ~new_R2144_U199;
  assign new_R2144_U162 = ~new_U2750 | ~new_R2144_U184;
  assign new_R2144_U163 = ~new_R2144_U116 | ~new_R2144_U109;
  assign new_R2144_U164 = ~new_U2355 | ~new_R2144_U68;
  assign new_R2144_U165 = ~new_U2762 | ~new_R2144_U12;
  assign new_R2144_U166 = ~new_U2355 | ~new_R2144_U69;
  assign new_R2144_U167 = ~new_U2761 | ~new_R2144_U12;
  assign new_R2144_U168 = ~new_U2355 | ~new_R2144_U70;
  assign new_R2144_U169 = ~new_U2763 | ~new_R2144_U12;
  assign new_R2144_U170 = ~new_R2144_U169 | ~new_R2144_U168;
  assign new_R2144_U171 = ~new_U2355 | ~new_R2144_U68;
  assign new_R2144_U172 = ~new_U2762 | ~new_R2144_U12;
  assign new_R2144_U173 = ~new_R2144_U172 | ~new_R2144_U171;
  assign new_R2144_U174 = ~new_U2355 | ~new_R2144_U70;
  assign new_R2144_U175 = ~new_U2763 | ~new_R2144_U12;
  assign new_R2144_U176 = ~new_U2355 | ~new_R2144_U71;
  assign new_R2144_U177 = ~new_U2764 | ~new_R2144_U12;
  assign new_R2144_U178 = ~new_R2144_U177 | ~new_R2144_U176;
  assign new_R2144_U179 = ~new_U2355 | ~new_R2144_U69;
  assign new_R2144_U180 = ~new_U2761 | ~new_R2144_U12;
  assign new_R2144_U181 = ~new_R2144_U180 | ~new_R2144_U179;
  assign new_R2144_U182 = ~new_U2355 | ~new_R2144_U72;
  assign new_R2144_U183 = ~new_U2766 | ~new_R2144_U12;
  assign new_R2144_U184 = ~new_R2144_U183 | ~new_R2144_U182;
  assign new_R2144_U185 = ~new_U2355 | ~new_R2144_U73;
  assign new_R2144_U186 = ~new_U2767 | ~new_R2144_U12;
  assign new_R2144_U187 = ~new_R2144_U28;
  assign new_R2144_U188 = ~new_U2355 | ~new_R2144_U74;
  assign new_R2144_U189 = ~new_U2768 | ~new_R2144_U12;
  assign new_R2144_U190 = ~new_U2355 | ~new_R2144_U74;
  assign new_R2144_U191 = ~new_U2768 | ~new_R2144_U12;
  assign new_R2144_U192 = ~new_R2144_U191 | ~new_R2144_U190;
  assign new_R2144_U193 = ~new_U2355 | ~new_R2144_U72;
  assign new_R2144_U194 = ~new_U2766 | ~new_R2144_U12;
  assign new_R2144_U195 = ~new_U2355 | ~new_R2144_U75;
  assign new_R2144_U196 = ~new_U2765 | ~new_R2144_U12;
  assign new_R2144_U197 = ~new_U2355 | ~new_R2144_U75;
  assign new_R2144_U198 = ~new_U2765 | ~new_R2144_U12;
  assign new_R2144_U199 = ~new_R2144_U198 | ~new_R2144_U197;
  assign new_R2144_U200 = ~new_U2355 | ~new_R2144_U71;
  assign new_R2144_U201 = ~new_U2764 | ~new_R2144_U12;
  assign new_R2144_U202 = ~new_U2355 | ~new_R2144_U76;
  assign new_R2144_U203 = ~new_U2760 | ~new_R2144_U12;
  assign new_R2144_U204 = ~new_R2144_U29;
  assign new_R2144_U205 = ~new_U2355 | ~new_R2144_U77;
  assign new_R2144_U206 = ~new_U2759 | ~new_R2144_U12;
  assign new_R2144_U207 = ~new_R2144_U27;
  assign new_R2144_U208 = ~new_R2144_U122 | ~new_R2144_U207;
  assign new_R2144_U209 = ~new_R2144_U27 | ~new_R2144_U78;
  assign new_R2144_U210 = ~new_R2144_U121 | ~new_R2144_U204;
  assign new_R2144_U211 = ~new_R2144_U29 | ~new_R2144_U79;
  assign new_R2144_U212 = ~new_R2144_U23 | ~new_R2144_U57 | ~new_R2144_U124;
  assign new_R2144_U213 = ~new_R2144_U5 | ~new_R2144_U108;
  assign new_R2144_U214 = ~new_R2144_U102 | ~new_R2144_U156;
  assign new_R2144_U215 = ~new_R2144_U81 | ~new_R2144_U59 | ~new_R2144_U160;
  assign new_R2144_U216 = ~new_R2144_U149 | ~new_R2144_U83;
  assign new_R2144_U217 = ~new_R2144_U44 | ~new_R2144_U123;
  assign new_R2144_U218 = ~new_R2144_U150 | ~new_R2144_U84;
  assign new_R2144_U219 = ~new_R2144_U46 | ~new_R2144_U119;
  assign new_R2144_U220 = ~new_U2355 | ~new_R2144_U85;
  assign new_R2144_U221 = ~new_U2754 | ~new_R2144_U12;
  assign new_R2144_U222 = ~new_R2144_U32;
  assign new_R2144_U223 = ~new_U2355 | ~new_R2144_U86;
  assign new_R2144_U224 = ~new_U2753 | ~new_R2144_U12;
  assign new_R2144_U225 = ~new_R2144_U31;
  assign new_R2144_U226 = ~new_U2355 | ~new_R2144_U87;
  assign new_R2144_U227 = ~new_U2755 | ~new_R2144_U12;
  assign new_R2144_U228 = ~new_R2144_U33;
  assign new_R2144_U229 = ~new_U2355 | ~new_R2144_U88;
  assign new_R2144_U230 = ~new_U2756 | ~new_R2144_U12;
  assign new_R2144_U231 = ~new_R2144_U34;
  assign new_R2144_U232 = ~new_U2355 | ~new_R2144_U89;
  assign new_R2144_U233 = ~new_U2757 | ~new_R2144_U12;
  assign new_R2144_U234 = ~new_R2144_U35;
  assign new_R2144_U235 = ~new_U2355 | ~new_R2144_U90;
  assign new_R2144_U236 = ~new_U2758 | ~new_R2144_U12;
  assign new_R2144_U237 = ~new_R2144_U36;
  assign new_R2144_U238 = ~new_R2144_U163 | ~new_R2144_U91;
  assign new_R2144_U239 = ~new_R2144_U48 | ~new_R2144_U133;
  assign new_R2144_U240 = ~new_R2144_U187 | ~new_U2751;
  assign new_R2144_U241 = ~new_R2144_U28 | ~new_R2144_U14;
  assign new_R2144_U242 = ~new_R2144_U187 | ~new_U2751;
  assign new_R2144_U243 = ~new_R2144_U28 | ~new_R2144_U14;
  assign new_R2144_U244 = ~new_R2144_U243 | ~new_R2144_U242;
  assign new_R2144_U245 = ~new_R2144_U92 | ~new_R2144_U93;
  assign new_R2144_U246 = ~new_R2144_U130 | ~new_R2144_U244;
  assign new_R2144_U247 = ~new_R2144_U147 | ~new_R2144_U225;
  assign new_R2144_U248 = ~new_R2144_U31 | ~new_R2144_U94;
  assign new_R2144_U249 = ~new_R2144_U222 | ~new_R2144_U143;
  assign new_R2144_U250 = ~new_R2144_U32 | ~new_R2144_U26;
  assign new_R2144_U251 = ~new_R2144_U142 | ~new_R2144_U228;
  assign new_R2144_U252 = ~new_R2144_U33 | ~new_R2144_U95;
  assign new_R2144_U253 = ~new_R2144_U231 | ~new_R2144_U141;
  assign new_R2144_U254 = ~new_R2144_U34 | ~new_R2144_U25;
  assign new_R2144_U255 = ~new_R2144_U140 | ~new_R2144_U234;
  assign new_R2144_U256 = ~new_R2144_U35 | ~new_R2144_U96;
  assign new_R2144_U257 = ~new_R2144_U139 | ~new_R2144_U237;
  assign new_R2144_U258 = ~new_R2144_U36 | ~new_R2144_U97;
  assign new_R2144_U259 = ~new_U2355 | ~new_R2144_U98;
  assign new_R2144_U260 = ~new_R2144_U148 | ~new_R2144_U12;
  assign new_LT_589_U6 = new_LT_589_U8 | new_U2673;
  assign new_LT_589_U7 = new_R584_U7 & new_R584_U6;
  assign new_LT_589_U8 = ~new_R584_U8 & ~new_LT_589_U7 & ~new_R584_U9;
  assign new_R584_U6 = ~new_U2676;
  assign new_R584_U7 = ~new_U2677;
  assign new_R584_U8 = ~new_U2674;
  assign new_R584_U9 = ~new_U2675;
  assign new_R2099_U4 = ~new_U4178;
  assign new_R2099_U5 = ~new_U4177;
  assign new_R2099_U6 = ~new_U2678;
  assign new_R2099_U7 = ~new_R2099_U88 | ~new_R2099_U137;
  assign new_R2099_U8 = ~new_R2099_U89 | ~new_R2099_U155;
  assign new_R2099_U9 = ~new_R2099_U90 | ~new_R2099_U157;
  assign new_R2099_U10 = ~new_R2099_U91 | ~new_R2099_U159;
  assign new_R2099_U11 = ~new_R2099_U92 | ~new_R2099_U161;
  assign new_R2099_U12 = ~new_R2099_U93 | ~new_R2099_U163;
  assign new_R2099_U13 = ~new_R2099_U94 | ~new_R2099_U165;
  assign new_R2099_U14 = ~new_R2099_U95 | ~new_R2099_U167;
  assign new_R2099_U15 = ~new_R2099_U169 | ~new_R2099_U55;
  assign new_R2099_U16 = ~new_R2099_U170 | ~new_R2099_U54;
  assign new_R2099_U17 = ~new_R2099_U171 | ~new_R2099_U53;
  assign new_R2099_U18 = ~new_R2099_U172 | ~new_R2099_U52;
  assign new_R2099_U19 = ~new_R2099_U173 | ~new_R2099_U51;
  assign new_R2099_U20 = ~new_R2099_U174 | ~new_R2099_U50;
  assign new_R2099_U21 = ~new_R2099_U175 | ~new_R2099_U49;
  assign new_R2099_U22 = ~new_R2099_U176 | ~new_R2099_U48;
  assign new_R2099_U23 = ~new_R2099_U177 | ~new_R2099_U47;
  assign new_R2099_U24 = ~new_R2099_U178 | ~new_R2099_U46;
  assign new_R2099_U25 = ~new_R2099_U179 | ~new_R2099_U45;
  assign new_R2099_U26 = ~new_R2099_U210 | ~new_R2099_U209;
  assign new_R2099_U27 = ~new_R2099_U183 | ~new_R2099_U182;
  assign new_R2099_U28 = ~new_R2099_U204 | ~new_R2099_U203;
  assign new_R2099_U29 = ~new_R2099_U207 | ~new_R2099_U206;
  assign new_R2099_U30 = ~new_R2099_U198 | ~new_R2099_U197;
  assign new_R2099_U31 = ~new_R2099_U201 | ~new_R2099_U200;
  assign new_R2099_U32 = ~new_R2099_U186 | ~new_R2099_U185;
  assign new_R2099_U33 = ~new_R2099_U189 | ~new_R2099_U188;
  assign new_R2099_U34 = ~new_R2099_U195 | ~new_R2099_U194;
  assign new_R2099_U35 = ~new_R2099_U192 | ~new_R2099_U191;
  assign new_R2099_U36 = ~new_R2099_U213 | ~new_R2099_U212;
  assign new_R2099_U37 = ~new_R2099_U215 | ~new_R2099_U214;
  assign new_R2099_U38 = ~new_R2099_U217 | ~new_R2099_U216;
  assign new_R2099_U39 = ~new_R2099_U219 | ~new_R2099_U218;
  assign new_R2099_U40 = ~new_R2099_U221 | ~new_R2099_U220;
  assign new_R2099_U41 = ~new_R2099_U223 | ~new_R2099_U222;
  assign new_R2099_U42 = ~new_R2099_U225 | ~new_R2099_U224;
  assign new_R2099_U43 = ~new_R2099_U284 | ~new_R2099_U283;
  assign new_R2099_U44 = ~new_R2099_U287 | ~new_R2099_U286;
  assign new_R2099_U45 = ~new_R2099_U227 | ~new_R2099_U226;
  assign new_R2099_U46 = ~new_R2099_U230 | ~new_R2099_U229;
  assign new_R2099_U47 = ~new_R2099_U233 | ~new_R2099_U232;
  assign new_R2099_U48 = ~new_R2099_U236 | ~new_R2099_U235;
  assign new_R2099_U49 = ~new_R2099_U239 | ~new_R2099_U238;
  assign new_R2099_U50 = ~new_R2099_U242 | ~new_R2099_U241;
  assign new_R2099_U51 = ~new_R2099_U245 | ~new_R2099_U244;
  assign new_R2099_U52 = ~new_R2099_U248 | ~new_R2099_U247;
  assign new_R2099_U53 = ~new_R2099_U251 | ~new_R2099_U250;
  assign new_R2099_U54 = ~new_R2099_U254 | ~new_R2099_U253;
  assign new_R2099_U55 = ~new_R2099_U257 | ~new_R2099_U256;
  assign new_R2099_U56 = ~new_R2099_U278 | ~new_R2099_U277;
  assign new_R2099_U57 = ~new_R2099_U281 | ~new_R2099_U280;
  assign new_R2099_U58 = ~new_R2099_U272 | ~new_R2099_U271;
  assign new_R2099_U59 = ~new_R2099_U275 | ~new_R2099_U274;
  assign new_R2099_U60 = ~new_R2099_U266 | ~new_R2099_U265;
  assign new_R2099_U61 = ~new_R2099_U269 | ~new_R2099_U268;
  assign new_R2099_U62 = ~new_R2099_U260 | ~new_R2099_U259;
  assign new_R2099_U63 = ~new_R2099_U263 | ~new_R2099_U262;
  assign new_R2099_U64 = ~new_R2099_U293 | ~new_R2099_U292;
  assign new_R2099_U65 = ~new_R2099_U295 | ~new_R2099_U294;
  assign new_R2099_U66 = ~new_R2099_U299 | ~new_R2099_U298;
  assign new_R2099_U67 = ~new_R2099_U301 | ~new_R2099_U300;
  assign new_R2099_U68 = ~new_R2099_U303 | ~new_R2099_U302;
  assign new_R2099_U69 = ~new_R2099_U305 | ~new_R2099_U304;
  assign new_R2099_U70 = ~new_R2099_U307 | ~new_R2099_U306;
  assign new_R2099_U71 = ~new_R2099_U309 | ~new_R2099_U308;
  assign new_R2099_U72 = ~new_R2099_U311 | ~new_R2099_U310;
  assign new_R2099_U73 = ~new_R2099_U313 | ~new_R2099_U312;
  assign new_R2099_U74 = ~new_R2099_U315 | ~new_R2099_U314;
  assign new_R2099_U75 = ~new_R2099_U317 | ~new_R2099_U316;
  assign new_R2099_U76 = ~new_R2099_U326 | ~new_R2099_U325;
  assign new_R2099_U77 = ~new_R2099_U328 | ~new_R2099_U327;
  assign new_R2099_U78 = ~new_R2099_U330 | ~new_R2099_U329;
  assign new_R2099_U79 = ~new_R2099_U332 | ~new_R2099_U331;
  assign new_R2099_U80 = ~new_R2099_U334 | ~new_R2099_U333;
  assign new_R2099_U81 = ~new_R2099_U336 | ~new_R2099_U335;
  assign new_R2099_U82 = ~new_R2099_U338 | ~new_R2099_U337;
  assign new_R2099_U83 = ~new_R2099_U340 | ~new_R2099_U339;
  assign new_R2099_U84 = ~new_R2099_U342 | ~new_R2099_U341;
  assign new_R2099_U85 = ~new_R2099_U344 | ~new_R2099_U343;
  assign new_R2099_U86 = ~new_R2099_U349 | ~new_R2099_U348;
  assign new_R2099_U87 = ~new_R2099_U324 | ~new_R2099_U323;
  assign new_R2099_U88 = new_R2099_U34 & new_R2099_U35;
  assign new_R2099_U89 = new_R2099_U31 & new_R2099_U30;
  assign new_R2099_U90 = new_R2099_U29 & new_R2099_U28;
  assign new_R2099_U91 = new_R2099_U26 & new_R2099_U27;
  assign new_R2099_U92 = new_R2099_U63 & new_R2099_U62;
  assign new_R2099_U93 = new_R2099_U61 & new_R2099_U60;
  assign new_R2099_U94 = new_R2099_U59 & new_R2099_U58;
  assign new_R2099_U95 = new_R2099_U57 & new_R2099_U56;
  assign new_R2099_U96 = new_R2099_U44 & new_R2099_U43;
  assign new_R2099_U97 = ~new_R2099_U290 | ~new_R2099_U289;
  assign new_R2099_U98 = ~new_R2099_U346 | ~new_R2099_U345;
  assign new_R2099_U99 = ~new_U2702;
  assign new_R2099_U100 = ~new_U2710;
  assign new_R2099_U101 = ~new_U2709;
  assign new_R2099_U102 = ~new_U2708;
  assign new_R2099_U103 = ~new_U2707;
  assign new_R2099_U104 = ~new_U2706;
  assign new_R2099_U105 = ~new_U2705;
  assign new_R2099_U106 = ~new_U2704;
  assign new_R2099_U107 = ~new_U2703;
  assign new_R2099_U108 = ~new_U2701;
  assign new_R2099_U109 = ~new_R2099_U159 | ~new_R2099_U27;
  assign new_R2099_U110 = ~new_R2099_U157 | ~new_R2099_U28;
  assign new_R2099_U111 = ~new_R2099_U155 | ~new_R2099_U30;
  assign new_R2099_U112 = ~new_R2099_U35 | ~new_R2099_U137;
  assign new_R2099_U113 = ~new_U2682;
  assign new_R2099_U114 = ~new_U2683;
  assign new_R2099_U115 = ~new_U2684;
  assign new_R2099_U116 = ~new_U2685;
  assign new_R2099_U117 = ~new_U2686;
  assign new_R2099_U118 = ~new_U2687;
  assign new_R2099_U119 = ~new_U2688;
  assign new_R2099_U120 = ~new_U2689;
  assign new_R2099_U121 = ~new_U2690;
  assign new_R2099_U122 = ~new_U2691;
  assign new_R2099_U123 = ~new_U2692;
  assign new_R2099_U124 = ~new_U2700;
  assign new_R2099_U125 = ~new_U2699;
  assign new_R2099_U126 = ~new_U2698;
  assign new_R2099_U127 = ~new_U2697;
  assign new_R2099_U128 = ~new_U2696;
  assign new_R2099_U129 = ~new_U2695;
  assign new_R2099_U130 = ~new_U2694;
  assign new_R2099_U131 = ~new_U2693;
  assign new_R2099_U132 = ~new_U2680;
  assign new_R2099_U133 = ~new_U2681;
  assign new_R2099_U134 = ~new_U2679;
  assign new_R2099_U135 = ~new_R2099_U96 | ~new_R2099_U180;
  assign new_R2099_U136 = ~new_R2099_U180 | ~new_R2099_U44;
  assign new_R2099_U137 = ~new_R2099_U152 | ~new_R2099_U151;
  assign new_R2099_U138 = new_R2099_U297 & new_R2099_U296;
  assign new_R2099_U139 = new_R2099_U319 & new_R2099_U318;
  assign new_R2099_U140 = ~new_R2099_U148 | ~new_R2099_U147;
  assign new_R2099_U141 = ~new_R2099_U167 | ~new_R2099_U56;
  assign new_R2099_U142 = ~new_R2099_U165 | ~new_R2099_U58;
  assign new_R2099_U143 = ~new_R2099_U163 | ~new_R2099_U60;
  assign new_R2099_U144 = ~new_R2099_U161 | ~new_R2099_U62;
  assign new_R2099_U145 = ~new_R2099_U135;
  assign new_R2099_U146 = new_U4178 | new_U4177;
  assign new_R2099_U147 = ~new_R2099_U32 | ~new_R2099_U146;
  assign new_R2099_U148 = ~new_U4177 | ~new_U4178;
  assign new_R2099_U149 = ~new_R2099_U140;
  assign new_R2099_U150 = ~new_R2099_U190 | ~new_R2099_U6;
  assign new_R2099_U151 = ~new_R2099_U150 | ~new_R2099_U140;
  assign new_R2099_U152 = ~new_U2678 | ~new_R2099_U33;
  assign new_R2099_U153 = ~new_R2099_U137;
  assign new_R2099_U154 = ~new_R2099_U112;
  assign new_R2099_U155 = ~new_R2099_U7;
  assign new_R2099_U156 = ~new_R2099_U111;
  assign new_R2099_U157 = ~new_R2099_U8;
  assign new_R2099_U158 = ~new_R2099_U110;
  assign new_R2099_U159 = ~new_R2099_U9;
  assign new_R2099_U160 = ~new_R2099_U109;
  assign new_R2099_U161 = ~new_R2099_U10;
  assign new_R2099_U162 = ~new_R2099_U144;
  assign new_R2099_U163 = ~new_R2099_U11;
  assign new_R2099_U164 = ~new_R2099_U143;
  assign new_R2099_U165 = ~new_R2099_U12;
  assign new_R2099_U166 = ~new_R2099_U142;
  assign new_R2099_U167 = ~new_R2099_U13;
  assign new_R2099_U168 = ~new_R2099_U141;
  assign new_R2099_U169 = ~new_R2099_U14;
  assign new_R2099_U170 = ~new_R2099_U15;
  assign new_R2099_U171 = ~new_R2099_U16;
  assign new_R2099_U172 = ~new_R2099_U17;
  assign new_R2099_U173 = ~new_R2099_U18;
  assign new_R2099_U174 = ~new_R2099_U19;
  assign new_R2099_U175 = ~new_R2099_U20;
  assign new_R2099_U176 = ~new_R2099_U21;
  assign new_R2099_U177 = ~new_R2099_U22;
  assign new_R2099_U178 = ~new_R2099_U23;
  assign new_R2099_U179 = ~new_R2099_U24;
  assign new_R2099_U180 = ~new_R2099_U25;
  assign new_R2099_U181 = ~new_R2099_U136;
  assign new_R2099_U182 = ~new_U4178 | ~new_R2099_U99;
  assign new_R2099_U183 = ~new_U2702 | ~new_R2099_U4;
  assign new_R2099_U184 = ~new_R2099_U27;
  assign new_R2099_U185 = ~new_U4178 | ~new_R2099_U100;
  assign new_R2099_U186 = ~new_U2710 | ~new_R2099_U4;
  assign new_R2099_U187 = ~new_R2099_U32;
  assign new_R2099_U188 = ~new_U4178 | ~new_R2099_U101;
  assign new_R2099_U189 = ~new_U2709 | ~new_R2099_U4;
  assign new_R2099_U190 = ~new_R2099_U33;
  assign new_R2099_U191 = ~new_U4178 | ~new_R2099_U102;
  assign new_R2099_U192 = ~new_U2708 | ~new_R2099_U4;
  assign new_R2099_U193 = ~new_R2099_U35;
  assign new_R2099_U194 = ~new_U4178 | ~new_R2099_U103;
  assign new_R2099_U195 = ~new_U2707 | ~new_R2099_U4;
  assign new_R2099_U196 = ~new_R2099_U34;
  assign new_R2099_U197 = ~new_U4178 | ~new_R2099_U104;
  assign new_R2099_U198 = ~new_U2706 | ~new_R2099_U4;
  assign new_R2099_U199 = ~new_R2099_U30;
  assign new_R2099_U200 = ~new_U4178 | ~new_R2099_U105;
  assign new_R2099_U201 = ~new_U2705 | ~new_R2099_U4;
  assign new_R2099_U202 = ~new_R2099_U31;
  assign new_R2099_U203 = ~new_U4178 | ~new_R2099_U106;
  assign new_R2099_U204 = ~new_U2704 | ~new_R2099_U4;
  assign new_R2099_U205 = ~new_R2099_U28;
  assign new_R2099_U206 = ~new_U4178 | ~new_R2099_U107;
  assign new_R2099_U207 = ~new_U2703 | ~new_R2099_U4;
  assign new_R2099_U208 = ~new_R2099_U29;
  assign new_R2099_U209 = ~new_U4178 | ~new_R2099_U108;
  assign new_R2099_U210 = ~new_U2701 | ~new_R2099_U4;
  assign new_R2099_U211 = ~new_R2099_U26;
  assign new_R2099_U212 = ~new_R2099_U160 | ~new_R2099_U211;
  assign new_R2099_U213 = ~new_R2099_U26 | ~new_R2099_U109;
  assign new_R2099_U214 = ~new_R2099_U184 | ~new_R2099_U159;
  assign new_R2099_U215 = ~new_R2099_U27 | ~new_R2099_U9;
  assign new_R2099_U216 = ~new_R2099_U158 | ~new_R2099_U208;
  assign new_R2099_U217 = ~new_R2099_U29 | ~new_R2099_U110;
  assign new_R2099_U218 = ~new_R2099_U205 | ~new_R2099_U157;
  assign new_R2099_U219 = ~new_R2099_U28 | ~new_R2099_U8;
  assign new_R2099_U220 = ~new_R2099_U156 | ~new_R2099_U202;
  assign new_R2099_U221 = ~new_R2099_U31 | ~new_R2099_U111;
  assign new_R2099_U222 = ~new_R2099_U199 | ~new_R2099_U155;
  assign new_R2099_U223 = ~new_R2099_U30 | ~new_R2099_U7;
  assign new_R2099_U224 = ~new_R2099_U154 | ~new_R2099_U196;
  assign new_R2099_U225 = ~new_R2099_U34 | ~new_R2099_U112;
  assign new_R2099_U226 = ~new_U4178 | ~new_R2099_U113;
  assign new_R2099_U227 = ~new_U2682 | ~new_R2099_U4;
  assign new_R2099_U228 = ~new_R2099_U45;
  assign new_R2099_U229 = ~new_U4178 | ~new_R2099_U114;
  assign new_R2099_U230 = ~new_U2683 | ~new_R2099_U4;
  assign new_R2099_U231 = ~new_R2099_U46;
  assign new_R2099_U232 = ~new_U4178 | ~new_R2099_U115;
  assign new_R2099_U233 = ~new_U2684 | ~new_R2099_U4;
  assign new_R2099_U234 = ~new_R2099_U47;
  assign new_R2099_U235 = ~new_U4178 | ~new_R2099_U116;
  assign new_R2099_U236 = ~new_U2685 | ~new_R2099_U4;
  assign new_R2099_U237 = ~new_R2099_U48;
  assign new_R2099_U238 = ~new_U4178 | ~new_R2099_U117;
  assign new_R2099_U239 = ~new_U2686 | ~new_R2099_U4;
  assign new_R2099_U240 = ~new_R2099_U49;
  assign new_R2099_U241 = ~new_U4178 | ~new_R2099_U118;
  assign new_R2099_U242 = ~new_U2687 | ~new_R2099_U4;
  assign new_R2099_U243 = ~new_R2099_U50;
  assign new_R2099_U244 = ~new_U4178 | ~new_R2099_U119;
  assign new_R2099_U245 = ~new_U2688 | ~new_R2099_U4;
  assign new_R2099_U246 = ~new_R2099_U51;
  assign new_R2099_U247 = ~new_U4178 | ~new_R2099_U120;
  assign new_R2099_U248 = ~new_U2689 | ~new_R2099_U4;
  assign new_R2099_U249 = ~new_R2099_U52;
  assign new_R2099_U250 = ~new_U4178 | ~new_R2099_U121;
  assign new_R2099_U251 = ~new_U2690 | ~new_R2099_U4;
  assign new_R2099_U252 = ~new_R2099_U53;
  assign new_R2099_U253 = ~new_U4178 | ~new_R2099_U122;
  assign new_R2099_U254 = ~new_U2691 | ~new_R2099_U4;
  assign new_R2099_U255 = ~new_R2099_U54;
  assign new_R2099_U256 = ~new_U4178 | ~new_R2099_U123;
  assign new_R2099_U257 = ~new_U2692 | ~new_R2099_U4;
  assign new_R2099_U258 = ~new_R2099_U55;
  assign new_R2099_U259 = ~new_U4178 | ~new_R2099_U124;
  assign new_R2099_U260 = ~new_U2700 | ~new_R2099_U4;
  assign new_R2099_U261 = ~new_R2099_U62;
  assign new_R2099_U262 = ~new_U4178 | ~new_R2099_U125;
  assign new_R2099_U263 = ~new_U2699 | ~new_R2099_U4;
  assign new_R2099_U264 = ~new_R2099_U63;
  assign new_R2099_U265 = ~new_U4178 | ~new_R2099_U126;
  assign new_R2099_U266 = ~new_U2698 | ~new_R2099_U4;
  assign new_R2099_U267 = ~new_R2099_U60;
  assign new_R2099_U268 = ~new_U4178 | ~new_R2099_U127;
  assign new_R2099_U269 = ~new_U2697 | ~new_R2099_U4;
  assign new_R2099_U270 = ~new_R2099_U61;
  assign new_R2099_U271 = ~new_U4178 | ~new_R2099_U128;
  assign new_R2099_U272 = ~new_U2696 | ~new_R2099_U4;
  assign new_R2099_U273 = ~new_R2099_U58;
  assign new_R2099_U274 = ~new_U4178 | ~new_R2099_U129;
  assign new_R2099_U275 = ~new_U2695 | ~new_R2099_U4;
  assign new_R2099_U276 = ~new_R2099_U59;
  assign new_R2099_U277 = ~new_U4178 | ~new_R2099_U130;
  assign new_R2099_U278 = ~new_U2694 | ~new_R2099_U4;
  assign new_R2099_U279 = ~new_R2099_U56;
  assign new_R2099_U280 = ~new_U4178 | ~new_R2099_U131;
  assign new_R2099_U281 = ~new_U2693 | ~new_R2099_U4;
  assign new_R2099_U282 = ~new_R2099_U57;
  assign new_R2099_U283 = ~new_U4178 | ~new_R2099_U132;
  assign new_R2099_U284 = ~new_U2680 | ~new_R2099_U4;
  assign new_R2099_U285 = ~new_R2099_U43;
  assign new_R2099_U286 = ~new_U4178 | ~new_R2099_U133;
  assign new_R2099_U287 = ~new_U2681 | ~new_R2099_U4;
  assign new_R2099_U288 = ~new_R2099_U44;
  assign new_R2099_U289 = ~new_U4178 | ~new_R2099_U134;
  assign new_R2099_U290 = ~new_U2679 | ~new_R2099_U4;
  assign new_R2099_U291 = ~new_R2099_U97;
  assign new_R2099_U292 = ~new_R2099_U145 | ~new_R2099_U291;
  assign new_R2099_U293 = ~new_R2099_U97 | ~new_R2099_U135;
  assign new_R2099_U294 = ~new_R2099_U181 | ~new_R2099_U285;
  assign new_R2099_U295 = ~new_R2099_U43 | ~new_R2099_U136;
  assign new_R2099_U296 = ~new_R2099_U153 | ~new_R2099_U193;
  assign new_R2099_U297 = ~new_R2099_U35 | ~new_R2099_U137;
  assign new_R2099_U298 = ~new_R2099_U288 | ~new_R2099_U180;
  assign new_R2099_U299 = ~new_R2099_U44 | ~new_R2099_U25;
  assign new_R2099_U300 = ~new_R2099_U228 | ~new_R2099_U179;
  assign new_R2099_U301 = ~new_R2099_U45 | ~new_R2099_U24;
  assign new_R2099_U302 = ~new_R2099_U231 | ~new_R2099_U178;
  assign new_R2099_U303 = ~new_R2099_U46 | ~new_R2099_U23;
  assign new_R2099_U304 = ~new_R2099_U234 | ~new_R2099_U177;
  assign new_R2099_U305 = ~new_R2099_U47 | ~new_R2099_U22;
  assign new_R2099_U306 = ~new_R2099_U237 | ~new_R2099_U176;
  assign new_R2099_U307 = ~new_R2099_U48 | ~new_R2099_U21;
  assign new_R2099_U308 = ~new_R2099_U240 | ~new_R2099_U175;
  assign new_R2099_U309 = ~new_R2099_U49 | ~new_R2099_U20;
  assign new_R2099_U310 = ~new_R2099_U243 | ~new_R2099_U174;
  assign new_R2099_U311 = ~new_R2099_U50 | ~new_R2099_U19;
  assign new_R2099_U312 = ~new_R2099_U246 | ~new_R2099_U173;
  assign new_R2099_U313 = ~new_R2099_U51 | ~new_R2099_U18;
  assign new_R2099_U314 = ~new_R2099_U249 | ~new_R2099_U172;
  assign new_R2099_U315 = ~new_R2099_U52 | ~new_R2099_U17;
  assign new_R2099_U316 = ~new_R2099_U252 | ~new_R2099_U171;
  assign new_R2099_U317 = ~new_R2099_U53 | ~new_R2099_U16;
  assign new_R2099_U318 = ~new_R2099_U190 | ~new_U2678;
  assign new_R2099_U319 = ~new_R2099_U33 | ~new_R2099_U6;
  assign new_R2099_U320 = ~new_R2099_U190 | ~new_U2678;
  assign new_R2099_U321 = ~new_R2099_U33 | ~new_R2099_U6;
  assign new_R2099_U322 = ~new_R2099_U321 | ~new_R2099_U320;
  assign new_R2099_U323 = ~new_R2099_U139 | ~new_R2099_U140;
  assign new_R2099_U324 = ~new_R2099_U149 | ~new_R2099_U322;
  assign new_R2099_U325 = ~new_R2099_U255 | ~new_R2099_U170;
  assign new_R2099_U326 = ~new_R2099_U54 | ~new_R2099_U15;
  assign new_R2099_U327 = ~new_R2099_U258 | ~new_R2099_U169;
  assign new_R2099_U328 = ~new_R2099_U55 | ~new_R2099_U14;
  assign new_R2099_U329 = ~new_R2099_U168 | ~new_R2099_U282;
  assign new_R2099_U330 = ~new_R2099_U57 | ~new_R2099_U141;
  assign new_R2099_U331 = ~new_R2099_U279 | ~new_R2099_U167;
  assign new_R2099_U332 = ~new_R2099_U56 | ~new_R2099_U13;
  assign new_R2099_U333 = ~new_R2099_U166 | ~new_R2099_U276;
  assign new_R2099_U334 = ~new_R2099_U59 | ~new_R2099_U142;
  assign new_R2099_U335 = ~new_R2099_U273 | ~new_R2099_U165;
  assign new_R2099_U336 = ~new_R2099_U58 | ~new_R2099_U12;
  assign new_R2099_U337 = ~new_R2099_U164 | ~new_R2099_U270;
  assign new_R2099_U338 = ~new_R2099_U61 | ~new_R2099_U143;
  assign new_R2099_U339 = ~new_R2099_U267 | ~new_R2099_U163;
  assign new_R2099_U340 = ~new_R2099_U60 | ~new_R2099_U11;
  assign new_R2099_U341 = ~new_R2099_U162 | ~new_R2099_U264;
  assign new_R2099_U342 = ~new_R2099_U63 | ~new_R2099_U144;
  assign new_R2099_U343 = ~new_R2099_U261 | ~new_R2099_U161;
  assign new_R2099_U344 = ~new_R2099_U62 | ~new_R2099_U10;
  assign new_R2099_U345 = ~new_U4177 | ~new_R2099_U4;
  assign new_R2099_U346 = ~new_U4178 | ~new_R2099_U5;
  assign new_R2099_U347 = ~new_R2099_U98;
  assign new_R2099_U348 = ~new_R2099_U32 | ~new_R2099_U347;
  assign new_R2099_U349 = ~new_R2099_U98 | ~new_R2099_U187;
  assign new_R2167_U6 = ~new_U2716;
  assign new_R2167_U7 = ~new_U2714;
  assign new_R2167_U8 = ~new_U2720;
  assign new_R2167_U9 = ~new_U2719;
  assign new_R2167_U10 = ~new_U2713;
  assign new_R2167_U11 = ~new_U2712;
  assign new_R2167_U12 = ~new_U2718;
  assign new_R2167_U13 = ~new_U2717;
  assign new_R2167_U14 = ~new_U2711;
  assign new_R2167_U15 = ~new_U2356;
  assign new_R2167_U16 = ~STATE2_REG_0_;
  assign new_R2167_U17 = ~new_R2167_U50 | ~new_R2167_U49;
  assign new_R2167_U18 = new_R2167_U29 & new_R2167_U30;
  assign new_R2167_U19 = new_R2167_U32 & new_R2167_U33;
  assign new_R2167_U20 = new_R2167_U35 & new_R2167_U36;
  assign new_R2167_U21 = new_R2167_U38 & new_R2167_U39;
  assign new_R2167_U22 = ~new_U2721;
  assign new_R2167_U23 = ~new_U2722;
  assign new_R2167_U24 = ~new_U2715 | ~new_R2167_U23;
  assign new_R2167_U25 = ~new_U2715 | ~new_R2167_U22;
  assign new_R2167_U26 = new_U2721 | new_U2722;
  assign new_R2167_U27 = ~new_U2714 | ~new_R2167_U8;
  assign new_R2167_U28 = ~new_R2167_U24 | ~new_R2167_U25 | ~new_R2167_U27 | ~new_R2167_U26;
  assign new_R2167_U29 = ~new_U2720 | ~new_R2167_U7;
  assign new_R2167_U30 = ~new_U2719 | ~new_R2167_U10;
  assign new_R2167_U31 = ~new_R2167_U18 | ~new_R2167_U28;
  assign new_R2167_U32 = ~new_U2713 | ~new_R2167_U9;
  assign new_R2167_U33 = ~new_U2712 | ~new_R2167_U12;
  assign new_R2167_U34 = ~new_R2167_U19 | ~new_R2167_U31;
  assign new_R2167_U35 = ~new_U2718 | ~new_R2167_U11;
  assign new_R2167_U36 = ~new_U2717 | ~new_R2167_U14;
  assign new_R2167_U37 = ~new_R2167_U20 | ~new_R2167_U34;
  assign new_R2167_U38 = ~new_U2711 | ~new_R2167_U13;
  assign new_R2167_U39 = ~new_U2356 | ~new_R2167_U6;
  assign new_R2167_U40 = ~new_R2167_U21 | ~new_R2167_U37;
  assign new_R2167_U41 = ~new_U2716 | ~new_R2167_U15;
  assign new_R2167_U42 = ~new_R2167_U40 | ~new_R2167_U41;
  assign new_R2167_U43 = ~new_U2716 | ~new_R2167_U16;
  assign new_R2167_U44 = ~new_R2167_U42 | ~new_R2167_U6;
  assign new_R2167_U45 = ~new_R2167_U44 | ~new_R2167_U43;
  assign new_R2167_U46 = ~STATE2_REG_0_ | ~new_R2167_U6;
  assign new_R2167_U47 = ~new_U2716 | ~new_R2167_U42;
  assign new_R2167_U48 = ~new_R2167_U47 | ~new_R2167_U46;
  assign new_R2167_U49 = ~new_R2167_U45 | ~new_R2167_U15;
  assign new_R2167_U50 = ~new_U2356 | ~new_R2167_U48;
  assign new_SUB_357_U6 = ~new_U3220;
  assign new_SUB_357_U7 = ~new_U3215;
  assign new_SUB_357_U8 = ~new_U3221;
  assign new_SUB_357_U9 = ~new_U3219;
  assign new_SUB_357_U10 = ~new_U3214;
  assign new_SUB_357_U11 = ~new_U3217;
  assign new_SUB_357_U12 = ~new_U3216;
  assign new_SUB_357_U13 = ~new_U3218;
  assign new_LT_563_1260_U6 = new_LT_563_1260_U9 & new_LT_563_1260_U8;
  assign new_LT_563_1260_U7 = ~new_U2673;
  assign new_LT_563_1260_U8 = ~new_R584_U8 | ~new_LT_563_1260_U7;
  assign new_LT_563_1260_U9 = ~new_R584_U9 | ~new_LT_563_1260_U7;
  assign new_SUB_580_U6 = ~new_SUB_580_U10 | ~new_SUB_580_U9;
  assign new_SUB_580_U7 = ~INSTADDRPOINTER_REG_1_;
  assign new_SUB_580_U8 = ~INSTADDRPOINTER_REG_0_;
  assign new_SUB_580_U9 = ~INSTADDRPOINTER_REG_1_ | ~new_SUB_580_U8;
  assign new_SUB_580_U10 = ~INSTADDRPOINTER_REG_0_ | ~new_SUB_580_U7;
  assign new_R2096_U4 = ~REIP_REG_1_;
  assign new_R2096_U5 = ~REIP_REG_2_;
  assign new_R2096_U6 = ~REIP_REG_2_ | ~REIP_REG_1_;
  assign new_R2096_U7 = ~REIP_REG_3_;
  assign new_R2096_U8 = ~REIP_REG_3_ | ~new_R2096_U94;
  assign new_R2096_U9 = ~REIP_REG_4_;
  assign new_R2096_U10 = ~REIP_REG_4_ | ~new_R2096_U95;
  assign new_R2096_U11 = ~REIP_REG_5_;
  assign new_R2096_U12 = ~REIP_REG_5_ | ~new_R2096_U96;
  assign new_R2096_U13 = ~REIP_REG_6_;
  assign new_R2096_U14 = ~REIP_REG_6_ | ~new_R2096_U97;
  assign new_R2096_U15 = ~REIP_REG_7_;
  assign new_R2096_U16 = ~REIP_REG_7_ | ~new_R2096_U98;
  assign new_R2096_U17 = ~REIP_REG_8_;
  assign new_R2096_U18 = ~REIP_REG_9_;
  assign new_R2096_U19 = ~REIP_REG_8_ | ~new_R2096_U99;
  assign new_R2096_U20 = ~new_R2096_U100 | ~REIP_REG_9_;
  assign new_R2096_U21 = ~REIP_REG_10_;
  assign new_R2096_U22 = ~REIP_REG_10_ | ~new_R2096_U101;
  assign new_R2096_U23 = ~REIP_REG_11_;
  assign new_R2096_U24 = ~REIP_REG_11_ | ~new_R2096_U102;
  assign new_R2096_U25 = ~REIP_REG_12_;
  assign new_R2096_U26 = ~REIP_REG_12_ | ~new_R2096_U103;
  assign new_R2096_U27 = ~REIP_REG_13_;
  assign new_R2096_U28 = ~REIP_REG_13_ | ~new_R2096_U104;
  assign new_R2096_U29 = ~REIP_REG_14_;
  assign new_R2096_U30 = ~REIP_REG_14_ | ~new_R2096_U105;
  assign new_R2096_U31 = ~REIP_REG_15_;
  assign new_R2096_U32 = ~REIP_REG_15_ | ~new_R2096_U106;
  assign new_R2096_U33 = ~REIP_REG_16_;
  assign new_R2096_U34 = ~REIP_REG_16_ | ~new_R2096_U107;
  assign new_R2096_U35 = ~REIP_REG_17_;
  assign new_R2096_U36 = ~REIP_REG_17_ | ~new_R2096_U108;
  assign new_R2096_U37 = ~REIP_REG_18_;
  assign new_R2096_U38 = ~REIP_REG_18_ | ~new_R2096_U109;
  assign new_R2096_U39 = ~REIP_REG_19_;
  assign new_R2096_U40 = ~REIP_REG_19_ | ~new_R2096_U110;
  assign new_R2096_U41 = ~REIP_REG_20_;
  assign new_R2096_U42 = ~REIP_REG_20_ | ~new_R2096_U111;
  assign new_R2096_U43 = ~REIP_REG_21_;
  assign new_R2096_U44 = ~REIP_REG_21_ | ~new_R2096_U112;
  assign new_R2096_U45 = ~REIP_REG_22_;
  assign new_R2096_U46 = ~REIP_REG_22_ | ~new_R2096_U113;
  assign new_R2096_U47 = ~REIP_REG_23_;
  assign new_R2096_U48 = ~REIP_REG_23_ | ~new_R2096_U114;
  assign new_R2096_U49 = ~REIP_REG_24_;
  assign new_R2096_U50 = ~REIP_REG_24_ | ~new_R2096_U115;
  assign new_R2096_U51 = ~REIP_REG_25_;
  assign new_R2096_U52 = ~REIP_REG_25_ | ~new_R2096_U116;
  assign new_R2096_U53 = ~REIP_REG_26_;
  assign new_R2096_U54 = ~REIP_REG_26_ | ~new_R2096_U117;
  assign new_R2096_U55 = ~REIP_REG_27_;
  assign new_R2096_U56 = ~REIP_REG_27_ | ~new_R2096_U118;
  assign new_R2096_U57 = ~REIP_REG_28_;
  assign new_R2096_U58 = ~REIP_REG_28_ | ~new_R2096_U119;
  assign new_R2096_U59 = ~REIP_REG_29_;
  assign new_R2096_U60 = ~REIP_REG_29_ | ~new_R2096_U120;
  assign new_R2096_U61 = ~REIP_REG_30_;
  assign new_R2096_U62 = ~new_R2096_U124 | ~new_R2096_U123;
  assign new_R2096_U63 = ~new_R2096_U126 | ~new_R2096_U125;
  assign new_R2096_U64 = ~new_R2096_U128 | ~new_R2096_U127;
  assign new_R2096_U65 = ~new_R2096_U130 | ~new_R2096_U129;
  assign new_R2096_U66 = ~new_R2096_U132 | ~new_R2096_U131;
  assign new_R2096_U67 = ~new_R2096_U134 | ~new_R2096_U133;
  assign new_R2096_U68 = ~new_R2096_U136 | ~new_R2096_U135;
  assign new_R2096_U69 = ~new_R2096_U138 | ~new_R2096_U137;
  assign new_R2096_U70 = ~new_R2096_U140 | ~new_R2096_U139;
  assign new_R2096_U71 = ~new_R2096_U142 | ~new_R2096_U141;
  assign new_R2096_U72 = ~new_R2096_U144 | ~new_R2096_U143;
  assign new_R2096_U73 = ~new_R2096_U146 | ~new_R2096_U145;
  assign new_R2096_U74 = ~new_R2096_U148 | ~new_R2096_U147;
  assign new_R2096_U75 = ~new_R2096_U150 | ~new_R2096_U149;
  assign new_R2096_U76 = ~new_R2096_U152 | ~new_R2096_U151;
  assign new_R2096_U77 = ~new_R2096_U154 | ~new_R2096_U153;
  assign new_R2096_U78 = ~new_R2096_U156 | ~new_R2096_U155;
  assign new_R2096_U79 = ~new_R2096_U158 | ~new_R2096_U157;
  assign new_R2096_U80 = ~new_R2096_U160 | ~new_R2096_U159;
  assign new_R2096_U81 = ~new_R2096_U162 | ~new_R2096_U161;
  assign new_R2096_U82 = ~new_R2096_U164 | ~new_R2096_U163;
  assign new_R2096_U83 = ~new_R2096_U166 | ~new_R2096_U165;
  assign new_R2096_U84 = ~new_R2096_U168 | ~new_R2096_U167;
  assign new_R2096_U85 = ~new_R2096_U170 | ~new_R2096_U169;
  assign new_R2096_U86 = ~new_R2096_U172 | ~new_R2096_U171;
  assign new_R2096_U87 = ~new_R2096_U174 | ~new_R2096_U173;
  assign new_R2096_U88 = ~new_R2096_U176 | ~new_R2096_U175;
  assign new_R2096_U89 = ~new_R2096_U178 | ~new_R2096_U177;
  assign new_R2096_U90 = ~new_R2096_U180 | ~new_R2096_U179;
  assign new_R2096_U91 = ~new_R2096_U182 | ~new_R2096_U181;
  assign new_R2096_U92 = ~REIP_REG_31_;
  assign new_R2096_U93 = ~REIP_REG_30_ | ~new_R2096_U121;
  assign new_R2096_U94 = ~new_R2096_U6;
  assign new_R2096_U95 = ~new_R2096_U8;
  assign new_R2096_U96 = ~new_R2096_U10;
  assign new_R2096_U97 = ~new_R2096_U12;
  assign new_R2096_U98 = ~new_R2096_U14;
  assign new_R2096_U99 = ~new_R2096_U16;
  assign new_R2096_U100 = ~new_R2096_U19;
  assign new_R2096_U101 = ~new_R2096_U20;
  assign new_R2096_U102 = ~new_R2096_U22;
  assign new_R2096_U103 = ~new_R2096_U24;
  assign new_R2096_U104 = ~new_R2096_U26;
  assign new_R2096_U105 = ~new_R2096_U28;
  assign new_R2096_U106 = ~new_R2096_U30;
  assign new_R2096_U107 = ~new_R2096_U32;
  assign new_R2096_U108 = ~new_R2096_U34;
  assign new_R2096_U109 = ~new_R2096_U36;
  assign new_R2096_U110 = ~new_R2096_U38;
  assign new_R2096_U111 = ~new_R2096_U40;
  assign new_R2096_U112 = ~new_R2096_U42;
  assign new_R2096_U113 = ~new_R2096_U44;
  assign new_R2096_U114 = ~new_R2096_U46;
  assign new_R2096_U115 = ~new_R2096_U48;
  assign new_R2096_U116 = ~new_R2096_U50;
  assign new_R2096_U117 = ~new_R2096_U52;
  assign new_R2096_U118 = ~new_R2096_U54;
  assign new_R2096_U119 = ~new_R2096_U56;
  assign new_R2096_U120 = ~new_R2096_U58;
  assign new_R2096_U121 = ~new_R2096_U60;
  assign new_R2096_U122 = ~new_R2096_U93;
  assign new_R2096_U123 = ~REIP_REG_9_ | ~new_R2096_U19;
  assign new_R2096_U124 = ~new_R2096_U100 | ~new_R2096_U18;
  assign new_R2096_U125 = ~REIP_REG_8_ | ~new_R2096_U16;
  assign new_R2096_U126 = ~new_R2096_U99 | ~new_R2096_U17;
  assign new_R2096_U127 = ~REIP_REG_7_ | ~new_R2096_U14;
  assign new_R2096_U128 = ~new_R2096_U98 | ~new_R2096_U15;
  assign new_R2096_U129 = ~REIP_REG_6_ | ~new_R2096_U12;
  assign new_R2096_U130 = ~new_R2096_U97 | ~new_R2096_U13;
  assign new_R2096_U131 = ~REIP_REG_5_ | ~new_R2096_U10;
  assign new_R2096_U132 = ~new_R2096_U96 | ~new_R2096_U11;
  assign new_R2096_U133 = ~REIP_REG_4_ | ~new_R2096_U8;
  assign new_R2096_U134 = ~new_R2096_U95 | ~new_R2096_U9;
  assign new_R2096_U135 = ~REIP_REG_3_ | ~new_R2096_U6;
  assign new_R2096_U136 = ~new_R2096_U94 | ~new_R2096_U7;
  assign new_R2096_U137 = ~REIP_REG_31_ | ~new_R2096_U93;
  assign new_R2096_U138 = ~new_R2096_U122 | ~new_R2096_U92;
  assign new_R2096_U139 = ~REIP_REG_30_ | ~new_R2096_U60;
  assign new_R2096_U140 = ~new_R2096_U121 | ~new_R2096_U61;
  assign new_R2096_U141 = ~REIP_REG_2_ | ~new_R2096_U4;
  assign new_R2096_U142 = ~REIP_REG_1_ | ~new_R2096_U5;
  assign new_R2096_U143 = ~REIP_REG_29_ | ~new_R2096_U58;
  assign new_R2096_U144 = ~new_R2096_U120 | ~new_R2096_U59;
  assign new_R2096_U145 = ~REIP_REG_28_ | ~new_R2096_U56;
  assign new_R2096_U146 = ~new_R2096_U119 | ~new_R2096_U57;
  assign new_R2096_U147 = ~REIP_REG_27_ | ~new_R2096_U54;
  assign new_R2096_U148 = ~new_R2096_U118 | ~new_R2096_U55;
  assign new_R2096_U149 = ~REIP_REG_26_ | ~new_R2096_U52;
  assign new_R2096_U150 = ~new_R2096_U117 | ~new_R2096_U53;
  assign new_R2096_U151 = ~REIP_REG_25_ | ~new_R2096_U50;
  assign new_R2096_U152 = ~new_R2096_U116 | ~new_R2096_U51;
  assign new_R2096_U153 = ~REIP_REG_24_ | ~new_R2096_U48;
  assign new_R2096_U154 = ~new_R2096_U115 | ~new_R2096_U49;
  assign new_R2096_U155 = ~REIP_REG_23_ | ~new_R2096_U46;
  assign new_R2096_U156 = ~new_R2096_U114 | ~new_R2096_U47;
  assign new_R2096_U157 = ~REIP_REG_22_ | ~new_R2096_U44;
  assign new_R2096_U158 = ~new_R2096_U113 | ~new_R2096_U45;
  assign new_R2096_U159 = ~REIP_REG_21_ | ~new_R2096_U42;
  assign new_R2096_U160 = ~new_R2096_U112 | ~new_R2096_U43;
  assign new_R2096_U161 = ~REIP_REG_20_ | ~new_R2096_U40;
  assign new_R2096_U162 = ~new_R2096_U111 | ~new_R2096_U41;
  assign new_R2096_U163 = ~REIP_REG_19_ | ~new_R2096_U38;
  assign new_R2096_U164 = ~new_R2096_U110 | ~new_R2096_U39;
  assign new_R2096_U165 = ~REIP_REG_18_ | ~new_R2096_U36;
  assign new_R2096_U166 = ~new_R2096_U109 | ~new_R2096_U37;
  assign new_R2096_U167 = ~REIP_REG_17_ | ~new_R2096_U34;
  assign new_R2096_U168 = ~new_R2096_U108 | ~new_R2096_U35;
  assign new_R2096_U169 = ~REIP_REG_16_ | ~new_R2096_U32;
  assign new_R2096_U170 = ~new_R2096_U107 | ~new_R2096_U33;
  assign new_R2096_U171 = ~REIP_REG_15_ | ~new_R2096_U30;
  assign new_R2096_U172 = ~new_R2096_U106 | ~new_R2096_U31;
  assign new_R2096_U173 = ~REIP_REG_14_ | ~new_R2096_U28;
  assign new_R2096_U174 = ~new_R2096_U105 | ~new_R2096_U29;
  assign new_R2096_U175 = ~REIP_REG_13_ | ~new_R2096_U26;
  assign new_R2096_U176 = ~new_R2096_U104 | ~new_R2096_U27;
  assign new_R2096_U177 = ~REIP_REG_12_ | ~new_R2096_U24;
  assign new_R2096_U178 = ~new_R2096_U103 | ~new_R2096_U25;
  assign new_R2096_U179 = ~REIP_REG_11_ | ~new_R2096_U22;
  assign new_R2096_U180 = ~new_R2096_U102 | ~new_R2096_U23;
  assign new_R2096_U181 = ~REIP_REG_10_ | ~new_R2096_U20;
  assign new_R2096_U182 = ~new_R2096_U101 | ~new_R2096_U21;
  assign new_LT_563_U6 = new_LT_563_U27 & new_LT_563_U26;
  assign new_LT_563_U7 = ~INSTQUEUEWR_ADDR_REG_2_;
  assign new_LT_563_U8 = ~new_U3478;
  assign new_LT_563_U9 = ~new_U3477;
  assign new_LT_563_U10 = ~INSTQUEUEWR_ADDR_REG_3_;
  assign new_LT_563_U11 = ~INSTQUEUEWR_ADDR_REG_4_;
  assign new_LT_563_U12 = ~new_U3476;
  assign new_LT_563_U13 = new_LT_563_U21 & new_LT_563_U22;
  assign new_LT_563_U14 = new_LT_563_U24 & new_LT_563_U25;
  assign new_LT_563_U15 = ~new_U3479;
  assign new_LT_563_U16 = ~new_U3480;
  assign new_LT_563_U17 = ~INSTQUEUEWR_ADDR_REG_0_ | ~new_LT_563_U16 | ~new_LT_563_U15;
  assign new_LT_563_U18 = ~INSTQUEUEWR_ADDR_REG_1_ | ~new_LT_563_U15;
  assign new_LT_563_U19 = ~INSTQUEUEWR_ADDR_REG_2_ | ~new_LT_563_U8;
  assign new_LT_563_U20 = ~new_LT_563_U17 | ~new_LT_563_U18 | ~new_LT_563_U28 | ~new_LT_563_U19;
  assign new_LT_563_U21 = ~new_U3478 | ~new_LT_563_U7;
  assign new_LT_563_U22 = ~new_U3477 | ~new_LT_563_U10;
  assign new_LT_563_U23 = ~new_LT_563_U13 | ~new_LT_563_U20;
  assign new_LT_563_U24 = ~INSTQUEUEWR_ADDR_REG_3_ | ~new_LT_563_U9;
  assign new_LT_563_U25 = ~INSTQUEUEWR_ADDR_REG_4_ | ~new_LT_563_U12;
  assign new_LT_563_U26 = ~new_LT_563_U14 | ~new_LT_563_U23;
  assign new_LT_563_U27 = ~new_U3476 | ~new_LT_563_U11;
  assign new_LT_563_U28 = ~new_LT_563_U16 | ~INSTQUEUEWR_ADDR_REG_0_ | ~INSTQUEUEWR_ADDR_REG_1_;
  assign new_R2238_U6 = ~new_R2238_U45 | ~new_R2238_U44;
  assign new_R2238_U7 = ~new_R2238_U9 | ~new_R2238_U46;
  assign new_R2238_U8 = ~INSTQUEUERD_ADDR_REG_0_;
  assign new_R2238_U9 = ~INSTQUEUERD_ADDR_REG_0_ | ~new_R2238_U18;
  assign new_R2238_U10 = ~INSTQUEUEWR_ADDR_REG_1_;
  assign new_R2238_U11 = ~INSTQUEUERD_ADDR_REG_2_;
  assign new_R2238_U12 = ~INSTQUEUEWR_ADDR_REG_2_;
  assign new_R2238_U13 = ~INSTQUEUERD_ADDR_REG_3_;
  assign new_R2238_U14 = ~INSTQUEUEWR_ADDR_REG_3_;
  assign new_R2238_U15 = ~INSTQUEUEWR_ADDR_REG_4_;
  assign new_R2238_U16 = ~new_R2238_U41 | ~new_R2238_U40;
  assign new_R2238_U17 = ~INSTQUEUERD_ADDR_REG_4_;
  assign new_R2238_U18 = ~INSTQUEUEWR_ADDR_REG_0_;
  assign new_R2238_U19 = ~new_R2238_U51 | ~new_R2238_U50;
  assign new_R2238_U20 = ~new_R2238_U56 | ~new_R2238_U55;
  assign new_R2238_U21 = ~new_R2238_U61 | ~new_R2238_U60;
  assign new_R2238_U22 = ~new_R2238_U66 | ~new_R2238_U65;
  assign new_R2238_U23 = ~new_R2238_U48 | ~new_R2238_U47;
  assign new_R2238_U24 = ~new_R2238_U53 | ~new_R2238_U52;
  assign new_R2238_U25 = ~new_R2238_U58 | ~new_R2238_U57;
  assign new_R2238_U26 = ~new_R2238_U63 | ~new_R2238_U62;
  assign new_R2238_U27 = ~new_R2238_U37 | ~new_R2238_U36;
  assign new_R2238_U28 = ~new_R2238_U33 | ~new_R2238_U32;
  assign new_R2238_U29 = ~INSTQUEUERD_ADDR_REG_1_;
  assign new_R2238_U30 = ~new_R2238_U9;
  assign new_R2238_U31 = ~new_R2238_U30 | ~new_R2238_U10;
  assign new_R2238_U32 = ~new_R2238_U31 | ~new_R2238_U29;
  assign new_R2238_U33 = ~INSTQUEUEWR_ADDR_REG_1_ | ~new_R2238_U9;
  assign new_R2238_U34 = ~new_R2238_U28;
  assign new_R2238_U35 = ~INSTQUEUERD_ADDR_REG_2_ | ~new_R2238_U12;
  assign new_R2238_U36 = ~new_R2238_U35 | ~new_R2238_U28;
  assign new_R2238_U37 = ~INSTQUEUEWR_ADDR_REG_2_ | ~new_R2238_U11;
  assign new_R2238_U38 = ~new_R2238_U27;
  assign new_R2238_U39 = ~INSTQUEUERD_ADDR_REG_3_ | ~new_R2238_U14;
  assign new_R2238_U40 = ~new_R2238_U39 | ~new_R2238_U27;
  assign new_R2238_U41 = ~INSTQUEUEWR_ADDR_REG_3_ | ~new_R2238_U13;
  assign new_R2238_U42 = ~new_R2238_U16;
  assign new_R2238_U43 = ~INSTQUEUEWR_ADDR_REG_4_ | ~new_R2238_U17;
  assign new_R2238_U44 = ~new_R2238_U42 | ~new_R2238_U43;
  assign new_R2238_U45 = ~INSTQUEUERD_ADDR_REG_4_ | ~new_R2238_U15;
  assign new_R2238_U46 = ~INSTQUEUEWR_ADDR_REG_0_ | ~new_R2238_U8;
  assign new_R2238_U47 = ~INSTQUEUERD_ADDR_REG_4_ | ~new_R2238_U15;
  assign new_R2238_U48 = ~INSTQUEUEWR_ADDR_REG_4_ | ~new_R2238_U17;
  assign new_R2238_U49 = ~new_R2238_U23;
  assign new_R2238_U50 = ~new_R2238_U49 | ~new_R2238_U42;
  assign new_R2238_U51 = ~new_R2238_U23 | ~new_R2238_U16;
  assign new_R2238_U52 = ~INSTQUEUERD_ADDR_REG_3_ | ~new_R2238_U14;
  assign new_R2238_U53 = ~INSTQUEUEWR_ADDR_REG_3_ | ~new_R2238_U13;
  assign new_R2238_U54 = ~new_R2238_U24;
  assign new_R2238_U55 = ~new_R2238_U38 | ~new_R2238_U54;
  assign new_R2238_U56 = ~new_R2238_U24 | ~new_R2238_U27;
  assign new_R2238_U57 = ~INSTQUEUERD_ADDR_REG_2_ | ~new_R2238_U12;
  assign new_R2238_U58 = ~INSTQUEUEWR_ADDR_REG_2_ | ~new_R2238_U11;
  assign new_R2238_U59 = ~new_R2238_U25;
  assign new_R2238_U60 = ~new_R2238_U34 | ~new_R2238_U59;
  assign new_R2238_U61 = ~new_R2238_U25 | ~new_R2238_U28;
  assign new_R2238_U62 = ~INSTQUEUERD_ADDR_REG_1_ | ~new_R2238_U10;
  assign new_R2238_U63 = ~INSTQUEUEWR_ADDR_REG_1_ | ~new_R2238_U29;
  assign new_R2238_U64 = ~new_R2238_U26;
  assign new_R2238_U65 = ~new_R2238_U64 | ~new_R2238_U30;
  assign new_R2238_U66 = ~new_R2238_U26 | ~new_R2238_U9;
  assign new_SUB_450_U6 = ~new_SUB_450_U45 | ~new_SUB_450_U44;
  assign new_SUB_450_U7 = ~new_SUB_450_U9 | ~new_SUB_450_U46;
  assign new_SUB_450_U8 = ~INSTQUEUERD_ADDR_REG_0_;
  assign new_SUB_450_U9 = ~INSTQUEUERD_ADDR_REG_0_ | ~new_SUB_450_U18;
  assign new_SUB_450_U10 = ~INSTQUEUEWR_ADDR_REG_1_;
  assign new_SUB_450_U11 = ~INSTQUEUERD_ADDR_REG_2_;
  assign new_SUB_450_U12 = ~INSTQUEUEWR_ADDR_REG_2_;
  assign new_SUB_450_U13 = ~INSTQUEUERD_ADDR_REG_3_;
  assign new_SUB_450_U14 = ~INSTQUEUEWR_ADDR_REG_3_;
  assign new_SUB_450_U15 = ~INSTQUEUEWR_ADDR_REG_4_;
  assign new_SUB_450_U16 = ~new_SUB_450_U41 | ~new_SUB_450_U40;
  assign new_SUB_450_U17 = ~INSTQUEUERD_ADDR_REG_4_;
  assign new_SUB_450_U18 = ~INSTQUEUEWR_ADDR_REG_0_;
  assign new_SUB_450_U19 = ~new_SUB_450_U51 | ~new_SUB_450_U50;
  assign new_SUB_450_U20 = ~new_SUB_450_U56 | ~new_SUB_450_U55;
  assign new_SUB_450_U21 = ~new_SUB_450_U61 | ~new_SUB_450_U60;
  assign new_SUB_450_U22 = ~new_SUB_450_U66 | ~new_SUB_450_U65;
  assign new_SUB_450_U23 = ~new_SUB_450_U48 | ~new_SUB_450_U47;
  assign new_SUB_450_U24 = ~new_SUB_450_U53 | ~new_SUB_450_U52;
  assign new_SUB_450_U25 = ~new_SUB_450_U58 | ~new_SUB_450_U57;
  assign new_SUB_450_U26 = ~new_SUB_450_U63 | ~new_SUB_450_U62;
  assign new_SUB_450_U27 = ~new_SUB_450_U37 | ~new_SUB_450_U36;
  assign new_SUB_450_U28 = ~new_SUB_450_U33 | ~new_SUB_450_U32;
  assign new_SUB_450_U29 = ~INSTQUEUERD_ADDR_REG_1_;
  assign new_SUB_450_U30 = ~new_SUB_450_U9;
  assign new_SUB_450_U31 = ~new_SUB_450_U30 | ~new_SUB_450_U10;
  assign new_SUB_450_U32 = ~new_SUB_450_U31 | ~new_SUB_450_U29;
  assign new_SUB_450_U33 = ~INSTQUEUEWR_ADDR_REG_1_ | ~new_SUB_450_U9;
  assign new_SUB_450_U34 = ~new_SUB_450_U28;
  assign new_SUB_450_U35 = ~INSTQUEUERD_ADDR_REG_2_ | ~new_SUB_450_U12;
  assign new_SUB_450_U36 = ~new_SUB_450_U35 | ~new_SUB_450_U28;
  assign new_SUB_450_U37 = ~INSTQUEUEWR_ADDR_REG_2_ | ~new_SUB_450_U11;
  assign new_SUB_450_U38 = ~new_SUB_450_U27;
  assign new_SUB_450_U39 = ~INSTQUEUERD_ADDR_REG_3_ | ~new_SUB_450_U14;
  assign new_SUB_450_U40 = ~new_SUB_450_U39 | ~new_SUB_450_U27;
  assign new_SUB_450_U41 = ~INSTQUEUEWR_ADDR_REG_3_ | ~new_SUB_450_U13;
  assign new_SUB_450_U42 = ~new_SUB_450_U16;
  assign new_SUB_450_U43 = ~INSTQUEUEWR_ADDR_REG_4_ | ~new_SUB_450_U17;
  assign new_SUB_450_U44 = ~new_SUB_450_U42 | ~new_SUB_450_U43;
  assign new_SUB_450_U45 = ~INSTQUEUERD_ADDR_REG_4_ | ~new_SUB_450_U15;
  assign new_SUB_450_U46 = ~INSTQUEUEWR_ADDR_REG_0_ | ~new_SUB_450_U8;
  assign new_SUB_450_U47 = ~INSTQUEUERD_ADDR_REG_4_ | ~new_SUB_450_U15;
  assign new_SUB_450_U48 = ~INSTQUEUEWR_ADDR_REG_4_ | ~new_SUB_450_U17;
  assign new_SUB_450_U49 = ~new_SUB_450_U23;
  assign new_SUB_450_U50 = ~new_SUB_450_U49 | ~new_SUB_450_U42;
  assign new_SUB_450_U51 = ~new_SUB_450_U23 | ~new_SUB_450_U16;
  assign new_SUB_450_U52 = ~INSTQUEUERD_ADDR_REG_3_ | ~new_SUB_450_U14;
  assign new_SUB_450_U53 = ~INSTQUEUEWR_ADDR_REG_3_ | ~new_SUB_450_U13;
  assign new_SUB_450_U54 = ~new_SUB_450_U24;
  assign new_SUB_450_U55 = ~new_SUB_450_U38 | ~new_SUB_450_U54;
  assign new_SUB_450_U56 = ~new_SUB_450_U24 | ~new_SUB_450_U27;
  assign new_SUB_450_U57 = ~INSTQUEUERD_ADDR_REG_2_ | ~new_SUB_450_U12;
  assign new_SUB_450_U58 = ~INSTQUEUEWR_ADDR_REG_2_ | ~new_SUB_450_U11;
  assign new_SUB_450_U59 = ~new_SUB_450_U25;
  assign new_SUB_450_U60 = ~new_SUB_450_U34 | ~new_SUB_450_U59;
  assign new_SUB_450_U61 = ~new_SUB_450_U25 | ~new_SUB_450_U28;
  assign new_SUB_450_U62 = ~INSTQUEUERD_ADDR_REG_1_ | ~new_SUB_450_U10;
  assign new_SUB_450_U63 = ~INSTQUEUEWR_ADDR_REG_1_ | ~new_SUB_450_U29;
  assign new_SUB_450_U64 = ~new_SUB_450_U26;
  assign new_SUB_450_U65 = ~new_SUB_450_U64 | ~new_SUB_450_U30;
  assign new_SUB_450_U66 = ~new_SUB_450_U26 | ~new_SUB_450_U9;
  assign new_ADD_371_U4 = ~new_U3214;
  assign new_ADD_371_U5 = ~new_ADD_371_U24 | ~new_ADD_371_U32;
  assign new_ADD_371_U6 = new_ADD_371_U22 & new_ADD_371_U30;
  assign new_ADD_371_U7 = ~new_U3215;
  assign new_ADD_371_U8 = ~new_U3217;
  assign new_ADD_371_U9 = ~new_U3217 | ~new_ADD_371_U24;
  assign new_ADD_371_U10 = ~new_U3218;
  assign new_ADD_371_U11 = ~new_U3218 | ~new_ADD_371_U28;
  assign new_ADD_371_U12 = ~new_U3219;
  assign new_ADD_371_U13 = ~new_U3219 | ~new_ADD_371_U29;
  assign new_ADD_371_U14 = ~new_U3221;
  assign new_ADD_371_U15 = ~new_U3220;
  assign new_ADD_371_U16 = ~new_U3216;
  assign new_ADD_371_U17 = ~new_ADD_371_U34 | ~new_ADD_371_U33;
  assign new_ADD_371_U18 = ~new_ADD_371_U36 | ~new_ADD_371_U35;
  assign new_ADD_371_U19 = ~new_ADD_371_U38 | ~new_ADD_371_U37;
  assign new_ADD_371_U20 = ~new_ADD_371_U40 | ~new_ADD_371_U39;
  assign new_ADD_371_U21 = ~new_ADD_371_U44 | ~new_ADD_371_U43;
  assign new_ADD_371_U22 = new_U3221 & new_U3220;
  assign new_ADD_371_U23 = ~new_U3220 | ~new_ADD_371_U30;
  assign new_ADD_371_U24 = ~new_ADD_371_U16 | ~new_ADD_371_U26;
  assign new_ADD_371_U25 = new_ADD_371_U42 & new_ADD_371_U41;
  assign new_ADD_371_U26 = ~new_U3215 | ~new_U3214;
  assign new_ADD_371_U27 = ~new_ADD_371_U24;
  assign new_ADD_371_U28 = ~new_ADD_371_U9;
  assign new_ADD_371_U29 = ~new_ADD_371_U11;
  assign new_ADD_371_U30 = ~new_ADD_371_U13;
  assign new_ADD_371_U31 = ~new_ADD_371_U23;
  assign new_ADD_371_U32 = ~new_U3216 | ~new_U3215 | ~new_U3214;
  assign new_ADD_371_U33 = ~new_U3221 | ~new_ADD_371_U23;
  assign new_ADD_371_U34 = ~new_ADD_371_U31 | ~new_ADD_371_U14;
  assign new_ADD_371_U35 = ~new_U3220 | ~new_ADD_371_U13;
  assign new_ADD_371_U36 = ~new_ADD_371_U30 | ~new_ADD_371_U15;
  assign new_ADD_371_U37 = ~new_U3219 | ~new_ADD_371_U11;
  assign new_ADD_371_U38 = ~new_ADD_371_U29 | ~new_ADD_371_U12;
  assign new_ADD_371_U39 = ~new_U3218 | ~new_ADD_371_U9;
  assign new_ADD_371_U40 = ~new_ADD_371_U28 | ~new_ADD_371_U10;
  assign new_ADD_371_U41 = ~new_U3217 | ~new_ADD_371_U24;
  assign new_ADD_371_U42 = ~new_ADD_371_U27 | ~new_ADD_371_U8;
  assign new_ADD_371_U43 = ~new_U3215 | ~new_ADD_371_U4;
  assign new_ADD_371_U44 = ~new_U3214 | ~new_ADD_371_U7;
  assign new_ADD_405_U4 = ~INSTADDRPOINTER_REG_0_;
  assign new_ADD_405_U5 = ~new_ADD_405_U92 | ~new_ADD_405_U126;
  assign new_ADD_405_U6 = ~INSTADDRPOINTER_REG_1_;
  assign new_ADD_405_U7 = ~INSTADDRPOINTER_REG_3_;
  assign new_ADD_405_U8 = ~INSTADDRPOINTER_REG_3_ | ~new_ADD_405_U92;
  assign new_ADD_405_U9 = ~INSTADDRPOINTER_REG_4_;
  assign new_ADD_405_U10 = ~INSTADDRPOINTER_REG_4_ | ~new_ADD_405_U98;
  assign new_ADD_405_U11 = ~INSTADDRPOINTER_REG_5_;
  assign new_ADD_405_U12 = ~INSTADDRPOINTER_REG_5_ | ~new_ADD_405_U99;
  assign new_ADD_405_U13 = ~INSTADDRPOINTER_REG_6_;
  assign new_ADD_405_U14 = ~INSTADDRPOINTER_REG_6_ | ~new_ADD_405_U100;
  assign new_ADD_405_U15 = ~INSTADDRPOINTER_REG_7_;
  assign new_ADD_405_U16 = ~INSTADDRPOINTER_REG_7_ | ~new_ADD_405_U101;
  assign new_ADD_405_U17 = ~INSTADDRPOINTER_REG_8_;
  assign new_ADD_405_U18 = ~INSTADDRPOINTER_REG_9_;
  assign new_ADD_405_U19 = ~INSTADDRPOINTER_REG_8_ | ~new_ADD_405_U102;
  assign new_ADD_405_U20 = ~new_ADD_405_U103 | ~INSTADDRPOINTER_REG_9_;
  assign new_ADD_405_U21 = ~INSTADDRPOINTER_REG_10_;
  assign new_ADD_405_U22 = ~INSTADDRPOINTER_REG_10_ | ~new_ADD_405_U104;
  assign new_ADD_405_U23 = ~INSTADDRPOINTER_REG_11_;
  assign new_ADD_405_U24 = ~INSTADDRPOINTER_REG_11_ | ~new_ADD_405_U105;
  assign new_ADD_405_U25 = ~INSTADDRPOINTER_REG_12_;
  assign new_ADD_405_U26 = ~INSTADDRPOINTER_REG_12_ | ~new_ADD_405_U106;
  assign new_ADD_405_U27 = ~INSTADDRPOINTER_REG_13_;
  assign new_ADD_405_U28 = ~INSTADDRPOINTER_REG_13_ | ~new_ADD_405_U107;
  assign new_ADD_405_U29 = ~INSTADDRPOINTER_REG_14_;
  assign new_ADD_405_U30 = ~INSTADDRPOINTER_REG_14_ | ~new_ADD_405_U108;
  assign new_ADD_405_U31 = ~INSTADDRPOINTER_REG_15_;
  assign new_ADD_405_U32 = ~INSTADDRPOINTER_REG_15_ | ~new_ADD_405_U109;
  assign new_ADD_405_U33 = ~INSTADDRPOINTER_REG_16_;
  assign new_ADD_405_U34 = ~INSTADDRPOINTER_REG_16_ | ~new_ADD_405_U110;
  assign new_ADD_405_U35 = ~INSTADDRPOINTER_REG_17_;
  assign new_ADD_405_U36 = ~INSTADDRPOINTER_REG_17_ | ~new_ADD_405_U111;
  assign new_ADD_405_U37 = ~INSTADDRPOINTER_REG_18_;
  assign new_ADD_405_U38 = ~INSTADDRPOINTER_REG_18_ | ~new_ADD_405_U112;
  assign new_ADD_405_U39 = ~INSTADDRPOINTER_REG_19_;
  assign new_ADD_405_U40 = ~INSTADDRPOINTER_REG_19_ | ~new_ADD_405_U113;
  assign new_ADD_405_U41 = ~INSTADDRPOINTER_REG_20_;
  assign new_ADD_405_U42 = ~INSTADDRPOINTER_REG_20_ | ~new_ADD_405_U114;
  assign new_ADD_405_U43 = ~INSTADDRPOINTER_REG_21_;
  assign new_ADD_405_U44 = ~INSTADDRPOINTER_REG_21_ | ~new_ADD_405_U115;
  assign new_ADD_405_U45 = ~INSTADDRPOINTER_REG_22_;
  assign new_ADD_405_U46 = ~INSTADDRPOINTER_REG_22_ | ~new_ADD_405_U116;
  assign new_ADD_405_U47 = ~INSTADDRPOINTER_REG_23_;
  assign new_ADD_405_U48 = ~INSTADDRPOINTER_REG_23_ | ~new_ADD_405_U117;
  assign new_ADD_405_U49 = ~INSTADDRPOINTER_REG_24_;
  assign new_ADD_405_U50 = ~INSTADDRPOINTER_REG_24_ | ~new_ADD_405_U118;
  assign new_ADD_405_U51 = ~INSTADDRPOINTER_REG_25_;
  assign new_ADD_405_U52 = ~INSTADDRPOINTER_REG_25_ | ~new_ADD_405_U119;
  assign new_ADD_405_U53 = ~INSTADDRPOINTER_REG_26_;
  assign new_ADD_405_U54 = ~INSTADDRPOINTER_REG_26_ | ~new_ADD_405_U120;
  assign new_ADD_405_U55 = ~INSTADDRPOINTER_REG_27_;
  assign new_ADD_405_U56 = ~INSTADDRPOINTER_REG_27_ | ~new_ADD_405_U121;
  assign new_ADD_405_U57 = ~INSTADDRPOINTER_REG_28_;
  assign new_ADD_405_U58 = ~INSTADDRPOINTER_REG_28_ | ~new_ADD_405_U122;
  assign new_ADD_405_U59 = ~INSTADDRPOINTER_REG_29_;
  assign new_ADD_405_U60 = ~INSTADDRPOINTER_REG_29_ | ~new_ADD_405_U123;
  assign new_ADD_405_U61 = ~INSTADDRPOINTER_REG_30_;
  assign new_ADD_405_U62 = ~INSTADDRPOINTER_REG_2_;
  assign new_ADD_405_U63 = ~new_ADD_405_U128 | ~new_ADD_405_U127;
  assign new_ADD_405_U64 = ~new_ADD_405_U130 | ~new_ADD_405_U129;
  assign new_ADD_405_U65 = ~new_ADD_405_U132 | ~new_ADD_405_U131;
  assign new_ADD_405_U66 = ~new_ADD_405_U134 | ~new_ADD_405_U133;
  assign new_ADD_405_U67 = ~new_ADD_405_U136 | ~new_ADD_405_U135;
  assign new_ADD_405_U68 = ~new_ADD_405_U138 | ~new_ADD_405_U137;
  assign new_ADD_405_U69 = ~new_ADD_405_U142 | ~new_ADD_405_U141;
  assign new_ADD_405_U70 = ~new_ADD_405_U144 | ~new_ADD_405_U143;
  assign new_ADD_405_U71 = ~new_ADD_405_U146 | ~new_ADD_405_U145;
  assign new_ADD_405_U72 = ~new_ADD_405_U148 | ~new_ADD_405_U147;
  assign new_ADD_405_U73 = ~new_ADD_405_U150 | ~new_ADD_405_U149;
  assign new_ADD_405_U74 = ~new_ADD_405_U152 | ~new_ADD_405_U151;
  assign new_ADD_405_U75 = ~new_ADD_405_U154 | ~new_ADD_405_U153;
  assign new_ADD_405_U76 = ~new_ADD_405_U156 | ~new_ADD_405_U155;
  assign new_ADD_405_U77 = ~new_ADD_405_U158 | ~new_ADD_405_U157;
  assign new_ADD_405_U78 = ~new_ADD_405_U160 | ~new_ADD_405_U159;
  assign new_ADD_405_U79 = ~new_ADD_405_U162 | ~new_ADD_405_U161;
  assign new_ADD_405_U80 = ~new_ADD_405_U164 | ~new_ADD_405_U163;
  assign new_ADD_405_U81 = ~new_ADD_405_U166 | ~new_ADD_405_U165;
  assign new_ADD_405_U82 = ~new_ADD_405_U168 | ~new_ADD_405_U167;
  assign new_ADD_405_U83 = ~new_ADD_405_U170 | ~new_ADD_405_U169;
  assign new_ADD_405_U84 = ~new_ADD_405_U172 | ~new_ADD_405_U171;
  assign new_ADD_405_U85 = ~new_ADD_405_U174 | ~new_ADD_405_U173;
  assign new_ADD_405_U86 = ~new_ADD_405_U176 | ~new_ADD_405_U175;
  assign new_ADD_405_U87 = ~new_ADD_405_U178 | ~new_ADD_405_U177;
  assign new_ADD_405_U88 = ~new_ADD_405_U180 | ~new_ADD_405_U179;
  assign new_ADD_405_U89 = ~new_ADD_405_U182 | ~new_ADD_405_U181;
  assign new_ADD_405_U90 = ~new_ADD_405_U184 | ~new_ADD_405_U183;
  assign new_ADD_405_U91 = ~new_ADD_405_U186 | ~new_ADD_405_U185;
  assign new_ADD_405_U92 = ~new_ADD_405_U62 | ~new_ADD_405_U96;
  assign new_ADD_405_U93 = new_ADD_405_U140 & new_ADD_405_U139;
  assign new_ADD_405_U94 = ~INSTADDRPOINTER_REG_31_;
  assign new_ADD_405_U95 = ~INSTADDRPOINTER_REG_30_ | ~new_ADD_405_U124;
  assign new_ADD_405_U96 = ~INSTADDRPOINTER_REG_1_ | ~INSTADDRPOINTER_REG_0_;
  assign new_ADD_405_U97 = ~new_ADD_405_U92;
  assign new_ADD_405_U98 = ~new_ADD_405_U8;
  assign new_ADD_405_U99 = ~new_ADD_405_U10;
  assign new_ADD_405_U100 = ~new_ADD_405_U12;
  assign new_ADD_405_U101 = ~new_ADD_405_U14;
  assign new_ADD_405_U102 = ~new_ADD_405_U16;
  assign new_ADD_405_U103 = ~new_ADD_405_U19;
  assign new_ADD_405_U104 = ~new_ADD_405_U20;
  assign new_ADD_405_U105 = ~new_ADD_405_U22;
  assign new_ADD_405_U106 = ~new_ADD_405_U24;
  assign new_ADD_405_U107 = ~new_ADD_405_U26;
  assign new_ADD_405_U108 = ~new_ADD_405_U28;
  assign new_ADD_405_U109 = ~new_ADD_405_U30;
  assign new_ADD_405_U110 = ~new_ADD_405_U32;
  assign new_ADD_405_U111 = ~new_ADD_405_U34;
  assign new_ADD_405_U112 = ~new_ADD_405_U36;
  assign new_ADD_405_U113 = ~new_ADD_405_U38;
  assign new_ADD_405_U114 = ~new_ADD_405_U40;
  assign new_ADD_405_U115 = ~new_ADD_405_U42;
  assign new_ADD_405_U116 = ~new_ADD_405_U44;
  assign new_ADD_405_U117 = ~new_ADD_405_U46;
  assign new_ADD_405_U118 = ~new_ADD_405_U48;
  assign new_ADD_405_U119 = ~new_ADD_405_U50;
  assign new_ADD_405_U120 = ~new_ADD_405_U52;
  assign new_ADD_405_U121 = ~new_ADD_405_U54;
  assign new_ADD_405_U122 = ~new_ADD_405_U56;
  assign new_ADD_405_U123 = ~new_ADD_405_U58;
  assign new_ADD_405_U124 = ~new_ADD_405_U60;
  assign new_ADD_405_U125 = ~new_ADD_405_U95;
  assign new_ADD_405_U126 = ~INSTADDRPOINTER_REG_2_ | ~INSTADDRPOINTER_REG_1_ | ~INSTADDRPOINTER_REG_0_;
  assign new_ADD_405_U127 = ~INSTADDRPOINTER_REG_9_ | ~new_ADD_405_U19;
  assign new_ADD_405_U128 = ~new_ADD_405_U103 | ~new_ADD_405_U18;
  assign new_ADD_405_U129 = ~INSTADDRPOINTER_REG_8_ | ~new_ADD_405_U16;
  assign new_ADD_405_U130 = ~new_ADD_405_U102 | ~new_ADD_405_U17;
  assign new_ADD_405_U131 = ~INSTADDRPOINTER_REG_7_ | ~new_ADD_405_U14;
  assign new_ADD_405_U132 = ~new_ADD_405_U101 | ~new_ADD_405_U15;
  assign new_ADD_405_U133 = ~INSTADDRPOINTER_REG_6_ | ~new_ADD_405_U12;
  assign new_ADD_405_U134 = ~new_ADD_405_U100 | ~new_ADD_405_U13;
  assign new_ADD_405_U135 = ~INSTADDRPOINTER_REG_5_ | ~new_ADD_405_U10;
  assign new_ADD_405_U136 = ~new_ADD_405_U99 | ~new_ADD_405_U11;
  assign new_ADD_405_U137 = ~INSTADDRPOINTER_REG_4_ | ~new_ADD_405_U8;
  assign new_ADD_405_U138 = ~new_ADD_405_U98 | ~new_ADD_405_U9;
  assign new_ADD_405_U139 = ~INSTADDRPOINTER_REG_3_ | ~new_ADD_405_U92;
  assign new_ADD_405_U140 = ~new_ADD_405_U97 | ~new_ADD_405_U7;
  assign new_ADD_405_U141 = ~INSTADDRPOINTER_REG_31_ | ~new_ADD_405_U95;
  assign new_ADD_405_U142 = ~new_ADD_405_U125 | ~new_ADD_405_U94;
  assign new_ADD_405_U143 = ~INSTADDRPOINTER_REG_30_ | ~new_ADD_405_U60;
  assign new_ADD_405_U144 = ~new_ADD_405_U124 | ~new_ADD_405_U61;
  assign new_ADD_405_U145 = ~INSTADDRPOINTER_REG_29_ | ~new_ADD_405_U58;
  assign new_ADD_405_U146 = ~new_ADD_405_U123 | ~new_ADD_405_U59;
  assign new_ADD_405_U147 = ~INSTADDRPOINTER_REG_28_ | ~new_ADD_405_U56;
  assign new_ADD_405_U148 = ~new_ADD_405_U122 | ~new_ADD_405_U57;
  assign new_ADD_405_U149 = ~INSTADDRPOINTER_REG_27_ | ~new_ADD_405_U54;
  assign new_ADD_405_U150 = ~new_ADD_405_U121 | ~new_ADD_405_U55;
  assign new_ADD_405_U151 = ~INSTADDRPOINTER_REG_26_ | ~new_ADD_405_U52;
  assign new_ADD_405_U152 = ~new_ADD_405_U120 | ~new_ADD_405_U53;
  assign new_ADD_405_U153 = ~INSTADDRPOINTER_REG_25_ | ~new_ADD_405_U50;
  assign new_ADD_405_U154 = ~new_ADD_405_U119 | ~new_ADD_405_U51;
  assign new_ADD_405_U155 = ~INSTADDRPOINTER_REG_24_ | ~new_ADD_405_U48;
  assign new_ADD_405_U156 = ~new_ADD_405_U118 | ~new_ADD_405_U49;
  assign new_ADD_405_U157 = ~INSTADDRPOINTER_REG_23_ | ~new_ADD_405_U46;
  assign new_ADD_405_U158 = ~new_ADD_405_U117 | ~new_ADD_405_U47;
  assign new_ADD_405_U159 = ~INSTADDRPOINTER_REG_22_ | ~new_ADD_405_U44;
  assign new_ADD_405_U160 = ~new_ADD_405_U116 | ~new_ADD_405_U45;
  assign new_ADD_405_U161 = ~INSTADDRPOINTER_REG_21_ | ~new_ADD_405_U42;
  assign new_ADD_405_U162 = ~new_ADD_405_U115 | ~new_ADD_405_U43;
  assign new_ADD_405_U163 = ~INSTADDRPOINTER_REG_20_ | ~new_ADD_405_U40;
  assign new_ADD_405_U164 = ~new_ADD_405_U114 | ~new_ADD_405_U41;
  assign new_ADD_405_U165 = ~INSTADDRPOINTER_REG_1_ | ~new_ADD_405_U4;
  assign new_ADD_405_U166 = ~INSTADDRPOINTER_REG_0_ | ~new_ADD_405_U6;
  assign new_ADD_405_U167 = ~INSTADDRPOINTER_REG_19_ | ~new_ADD_405_U38;
  assign new_ADD_405_U168 = ~new_ADD_405_U113 | ~new_ADD_405_U39;
  assign new_ADD_405_U169 = ~INSTADDRPOINTER_REG_18_ | ~new_ADD_405_U36;
  assign new_ADD_405_U170 = ~new_ADD_405_U112 | ~new_ADD_405_U37;
  assign new_ADD_405_U171 = ~INSTADDRPOINTER_REG_17_ | ~new_ADD_405_U34;
  assign new_ADD_405_U172 = ~new_ADD_405_U111 | ~new_ADD_405_U35;
  assign new_ADD_405_U173 = ~INSTADDRPOINTER_REG_16_ | ~new_ADD_405_U32;
  assign new_ADD_405_U174 = ~new_ADD_405_U110 | ~new_ADD_405_U33;
  assign new_ADD_405_U175 = ~INSTADDRPOINTER_REG_15_ | ~new_ADD_405_U30;
  assign new_ADD_405_U176 = ~new_ADD_405_U109 | ~new_ADD_405_U31;
  assign new_ADD_405_U177 = ~INSTADDRPOINTER_REG_14_ | ~new_ADD_405_U28;
  assign new_ADD_405_U178 = ~new_ADD_405_U108 | ~new_ADD_405_U29;
  assign new_ADD_405_U179 = ~INSTADDRPOINTER_REG_13_ | ~new_ADD_405_U26;
  assign new_ADD_405_U180 = ~new_ADD_405_U107 | ~new_ADD_405_U27;
  assign new_ADD_405_U181 = ~INSTADDRPOINTER_REG_12_ | ~new_ADD_405_U24;
  assign new_ADD_405_U182 = ~new_ADD_405_U106 | ~new_ADD_405_U25;
  assign new_ADD_405_U183 = ~INSTADDRPOINTER_REG_11_ | ~new_ADD_405_U22;
  assign new_ADD_405_U184 = ~new_ADD_405_U105 | ~new_ADD_405_U23;
  assign new_ADD_405_U185 = ~INSTADDRPOINTER_REG_10_ | ~new_ADD_405_U20;
  assign new_ADD_405_U186 = ~new_ADD_405_U104 | ~new_ADD_405_U21;
  assign new_GTE_485_U6 = ~new_R2238_U6 & ~new_GTE_485_U7;
  assign new_GTE_485_U7 = ~new_R2238_U21 & ~new_R2238_U22 & ~new_R2238_U19 & ~new_R2238_U20;
  assign new_ADD_515_U4 = ~INSTADDRPOINTER_REG_1_;
  assign new_ADD_515_U5 = ~INSTADDRPOINTER_REG_2_;
  assign new_ADD_515_U6 = ~INSTADDRPOINTER_REG_2_ | ~INSTADDRPOINTER_REG_1_;
  assign new_ADD_515_U7 = ~INSTADDRPOINTER_REG_3_;
  assign new_ADD_515_U8 = ~INSTADDRPOINTER_REG_3_ | ~new_ADD_515_U94;
  assign new_ADD_515_U9 = ~INSTADDRPOINTER_REG_4_;
  assign new_ADD_515_U10 = ~INSTADDRPOINTER_REG_4_ | ~new_ADD_515_U95;
  assign new_ADD_515_U11 = ~INSTADDRPOINTER_REG_5_;
  assign new_ADD_515_U12 = ~INSTADDRPOINTER_REG_5_ | ~new_ADD_515_U96;
  assign new_ADD_515_U13 = ~INSTADDRPOINTER_REG_6_;
  assign new_ADD_515_U14 = ~INSTADDRPOINTER_REG_6_ | ~new_ADD_515_U97;
  assign new_ADD_515_U15 = ~INSTADDRPOINTER_REG_7_;
  assign new_ADD_515_U16 = ~INSTADDRPOINTER_REG_7_ | ~new_ADD_515_U98;
  assign new_ADD_515_U17 = ~INSTADDRPOINTER_REG_8_;
  assign new_ADD_515_U18 = ~INSTADDRPOINTER_REG_9_;
  assign new_ADD_515_U19 = ~INSTADDRPOINTER_REG_8_ | ~new_ADD_515_U99;
  assign new_ADD_515_U20 = ~new_ADD_515_U100 | ~INSTADDRPOINTER_REG_9_;
  assign new_ADD_515_U21 = ~INSTADDRPOINTER_REG_10_;
  assign new_ADD_515_U22 = ~INSTADDRPOINTER_REG_10_ | ~new_ADD_515_U101;
  assign new_ADD_515_U23 = ~INSTADDRPOINTER_REG_11_;
  assign new_ADD_515_U24 = ~INSTADDRPOINTER_REG_11_ | ~new_ADD_515_U102;
  assign new_ADD_515_U25 = ~INSTADDRPOINTER_REG_12_;
  assign new_ADD_515_U26 = ~INSTADDRPOINTER_REG_12_ | ~new_ADD_515_U103;
  assign new_ADD_515_U27 = ~INSTADDRPOINTER_REG_13_;
  assign new_ADD_515_U28 = ~INSTADDRPOINTER_REG_13_ | ~new_ADD_515_U104;
  assign new_ADD_515_U29 = ~INSTADDRPOINTER_REG_14_;
  assign new_ADD_515_U30 = ~INSTADDRPOINTER_REG_14_ | ~new_ADD_515_U105;
  assign new_ADD_515_U31 = ~INSTADDRPOINTER_REG_15_;
  assign new_ADD_515_U32 = ~INSTADDRPOINTER_REG_15_ | ~new_ADD_515_U106;
  assign new_ADD_515_U33 = ~INSTADDRPOINTER_REG_16_;
  assign new_ADD_515_U34 = ~INSTADDRPOINTER_REG_16_ | ~new_ADD_515_U107;
  assign new_ADD_515_U35 = ~INSTADDRPOINTER_REG_17_;
  assign new_ADD_515_U36 = ~INSTADDRPOINTER_REG_17_ | ~new_ADD_515_U108;
  assign new_ADD_515_U37 = ~INSTADDRPOINTER_REG_18_;
  assign new_ADD_515_U38 = ~INSTADDRPOINTER_REG_18_ | ~new_ADD_515_U109;
  assign new_ADD_515_U39 = ~INSTADDRPOINTER_REG_19_;
  assign new_ADD_515_U40 = ~INSTADDRPOINTER_REG_19_ | ~new_ADD_515_U110;
  assign new_ADD_515_U41 = ~INSTADDRPOINTER_REG_20_;
  assign new_ADD_515_U42 = ~INSTADDRPOINTER_REG_20_ | ~new_ADD_515_U111;
  assign new_ADD_515_U43 = ~INSTADDRPOINTER_REG_21_;
  assign new_ADD_515_U44 = ~INSTADDRPOINTER_REG_21_ | ~new_ADD_515_U112;
  assign new_ADD_515_U45 = ~INSTADDRPOINTER_REG_22_;
  assign new_ADD_515_U46 = ~INSTADDRPOINTER_REG_22_ | ~new_ADD_515_U113;
  assign new_ADD_515_U47 = ~INSTADDRPOINTER_REG_23_;
  assign new_ADD_515_U48 = ~INSTADDRPOINTER_REG_23_ | ~new_ADD_515_U114;
  assign new_ADD_515_U49 = ~INSTADDRPOINTER_REG_24_;
  assign new_ADD_515_U50 = ~INSTADDRPOINTER_REG_24_ | ~new_ADD_515_U115;
  assign new_ADD_515_U51 = ~INSTADDRPOINTER_REG_25_;
  assign new_ADD_515_U52 = ~INSTADDRPOINTER_REG_25_ | ~new_ADD_515_U116;
  assign new_ADD_515_U53 = ~INSTADDRPOINTER_REG_26_;
  assign new_ADD_515_U54 = ~INSTADDRPOINTER_REG_26_ | ~new_ADD_515_U117;
  assign new_ADD_515_U55 = ~INSTADDRPOINTER_REG_27_;
  assign new_ADD_515_U56 = ~INSTADDRPOINTER_REG_27_ | ~new_ADD_515_U118;
  assign new_ADD_515_U57 = ~INSTADDRPOINTER_REG_28_;
  assign new_ADD_515_U58 = ~INSTADDRPOINTER_REG_28_ | ~new_ADD_515_U119;
  assign new_ADD_515_U59 = ~INSTADDRPOINTER_REG_29_;
  assign new_ADD_515_U60 = ~INSTADDRPOINTER_REG_29_ | ~new_ADD_515_U120;
  assign new_ADD_515_U61 = ~INSTADDRPOINTER_REG_30_;
  assign new_ADD_515_U62 = ~new_ADD_515_U124 | ~new_ADD_515_U123;
  assign new_ADD_515_U63 = ~new_ADD_515_U126 | ~new_ADD_515_U125;
  assign new_ADD_515_U64 = ~new_ADD_515_U128 | ~new_ADD_515_U127;
  assign new_ADD_515_U65 = ~new_ADD_515_U130 | ~new_ADD_515_U129;
  assign new_ADD_515_U66 = ~new_ADD_515_U132 | ~new_ADD_515_U131;
  assign new_ADD_515_U67 = ~new_ADD_515_U134 | ~new_ADD_515_U133;
  assign new_ADD_515_U68 = ~new_ADD_515_U136 | ~new_ADD_515_U135;
  assign new_ADD_515_U69 = ~new_ADD_515_U138 | ~new_ADD_515_U137;
  assign new_ADD_515_U70 = ~new_ADD_515_U140 | ~new_ADD_515_U139;
  assign new_ADD_515_U71 = ~new_ADD_515_U142 | ~new_ADD_515_U141;
  assign new_ADD_515_U72 = ~new_ADD_515_U144 | ~new_ADD_515_U143;
  assign new_ADD_515_U73 = ~new_ADD_515_U146 | ~new_ADD_515_U145;
  assign new_ADD_515_U74 = ~new_ADD_515_U148 | ~new_ADD_515_U147;
  assign new_ADD_515_U75 = ~new_ADD_515_U150 | ~new_ADD_515_U149;
  assign new_ADD_515_U76 = ~new_ADD_515_U152 | ~new_ADD_515_U151;
  assign new_ADD_515_U77 = ~new_ADD_515_U154 | ~new_ADD_515_U153;
  assign new_ADD_515_U78 = ~new_ADD_515_U156 | ~new_ADD_515_U155;
  assign new_ADD_515_U79 = ~new_ADD_515_U158 | ~new_ADD_515_U157;
  assign new_ADD_515_U80 = ~new_ADD_515_U160 | ~new_ADD_515_U159;
  assign new_ADD_515_U81 = ~new_ADD_515_U162 | ~new_ADD_515_U161;
  assign new_ADD_515_U82 = ~new_ADD_515_U164 | ~new_ADD_515_U163;
  assign new_ADD_515_U83 = ~new_ADD_515_U166 | ~new_ADD_515_U165;
  assign new_ADD_515_U84 = ~new_ADD_515_U168 | ~new_ADD_515_U167;
  assign new_ADD_515_U85 = ~new_ADD_515_U170 | ~new_ADD_515_U169;
  assign new_ADD_515_U86 = ~new_ADD_515_U172 | ~new_ADD_515_U171;
  assign new_ADD_515_U87 = ~new_ADD_515_U174 | ~new_ADD_515_U173;
  assign new_ADD_515_U88 = ~new_ADD_515_U176 | ~new_ADD_515_U175;
  assign new_ADD_515_U89 = ~new_ADD_515_U178 | ~new_ADD_515_U177;
  assign new_ADD_515_U90 = ~new_ADD_515_U180 | ~new_ADD_515_U179;
  assign new_ADD_515_U91 = ~new_ADD_515_U182 | ~new_ADD_515_U181;
  assign new_ADD_515_U92 = ~INSTADDRPOINTER_REG_31_;
  assign new_ADD_515_U93 = ~INSTADDRPOINTER_REG_30_ | ~new_ADD_515_U121;
  assign new_ADD_515_U94 = ~new_ADD_515_U6;
  assign new_ADD_515_U95 = ~new_ADD_515_U8;
  assign new_ADD_515_U96 = ~new_ADD_515_U10;
  assign new_ADD_515_U97 = ~new_ADD_515_U12;
  assign new_ADD_515_U98 = ~new_ADD_515_U14;
  assign new_ADD_515_U99 = ~new_ADD_515_U16;
  assign new_ADD_515_U100 = ~new_ADD_515_U19;
  assign new_ADD_515_U101 = ~new_ADD_515_U20;
  assign new_ADD_515_U102 = ~new_ADD_515_U22;
  assign new_ADD_515_U103 = ~new_ADD_515_U24;
  assign new_ADD_515_U104 = ~new_ADD_515_U26;
  assign new_ADD_515_U105 = ~new_ADD_515_U28;
  assign new_ADD_515_U106 = ~new_ADD_515_U30;
  assign new_ADD_515_U107 = ~new_ADD_515_U32;
  assign new_ADD_515_U108 = ~new_ADD_515_U34;
  assign new_ADD_515_U109 = ~new_ADD_515_U36;
  assign new_ADD_515_U110 = ~new_ADD_515_U38;
  assign new_ADD_515_U111 = ~new_ADD_515_U40;
  assign new_ADD_515_U112 = ~new_ADD_515_U42;
  assign new_ADD_515_U113 = ~new_ADD_515_U44;
  assign new_ADD_515_U114 = ~new_ADD_515_U46;
  assign new_ADD_515_U115 = ~new_ADD_515_U48;
  assign new_ADD_515_U116 = ~new_ADD_515_U50;
  assign new_ADD_515_U117 = ~new_ADD_515_U52;
  assign new_ADD_515_U118 = ~new_ADD_515_U54;
  assign new_ADD_515_U119 = ~new_ADD_515_U56;
  assign new_ADD_515_U120 = ~new_ADD_515_U58;
  assign new_ADD_515_U121 = ~new_ADD_515_U60;
  assign new_ADD_515_U122 = ~new_ADD_515_U93;
  assign new_ADD_515_U123 = ~INSTADDRPOINTER_REG_9_ | ~new_ADD_515_U19;
  assign new_ADD_515_U124 = ~new_ADD_515_U100 | ~new_ADD_515_U18;
  assign new_ADD_515_U125 = ~INSTADDRPOINTER_REG_8_ | ~new_ADD_515_U16;
  assign new_ADD_515_U126 = ~new_ADD_515_U99 | ~new_ADD_515_U17;
  assign new_ADD_515_U127 = ~INSTADDRPOINTER_REG_7_ | ~new_ADD_515_U14;
  assign new_ADD_515_U128 = ~new_ADD_515_U98 | ~new_ADD_515_U15;
  assign new_ADD_515_U129 = ~INSTADDRPOINTER_REG_6_ | ~new_ADD_515_U12;
  assign new_ADD_515_U130 = ~new_ADD_515_U97 | ~new_ADD_515_U13;
  assign new_ADD_515_U131 = ~INSTADDRPOINTER_REG_5_ | ~new_ADD_515_U10;
  assign new_ADD_515_U132 = ~new_ADD_515_U96 | ~new_ADD_515_U11;
  assign new_ADD_515_U133 = ~INSTADDRPOINTER_REG_4_ | ~new_ADD_515_U8;
  assign new_ADD_515_U134 = ~new_ADD_515_U95 | ~new_ADD_515_U9;
  assign new_ADD_515_U135 = ~INSTADDRPOINTER_REG_3_ | ~new_ADD_515_U6;
  assign new_ADD_515_U136 = ~new_ADD_515_U94 | ~new_ADD_515_U7;
  assign new_ADD_515_U137 = ~INSTADDRPOINTER_REG_31_ | ~new_ADD_515_U93;
  assign new_ADD_515_U138 = ~new_ADD_515_U122 | ~new_ADD_515_U92;
  assign new_ADD_515_U139 = ~INSTADDRPOINTER_REG_30_ | ~new_ADD_515_U60;
  assign new_ADD_515_U140 = ~new_ADD_515_U121 | ~new_ADD_515_U61;
  assign new_ADD_515_U141 = ~INSTADDRPOINTER_REG_2_ | ~new_ADD_515_U4;
  assign new_ADD_515_U142 = ~INSTADDRPOINTER_REG_1_ | ~new_ADD_515_U5;
  assign new_ADD_515_U143 = ~INSTADDRPOINTER_REG_29_ | ~new_ADD_515_U58;
  assign new_ADD_515_U144 = ~new_ADD_515_U120 | ~new_ADD_515_U59;
  assign new_ADD_515_U145 = ~INSTADDRPOINTER_REG_28_ | ~new_ADD_515_U56;
  assign new_ADD_515_U146 = ~new_ADD_515_U119 | ~new_ADD_515_U57;
  assign new_ADD_515_U147 = ~INSTADDRPOINTER_REG_27_ | ~new_ADD_515_U54;
  assign new_ADD_515_U148 = ~new_ADD_515_U118 | ~new_ADD_515_U55;
  assign new_ADD_515_U149 = ~INSTADDRPOINTER_REG_26_ | ~new_ADD_515_U52;
  assign new_ADD_515_U150 = ~new_ADD_515_U117 | ~new_ADD_515_U53;
  assign new_ADD_515_U151 = ~INSTADDRPOINTER_REG_25_ | ~new_ADD_515_U50;
  assign new_not_keyinput0 = ~keyinput0;
  assign new_not_keyinput1 = ~keyinput1;
  assign new_not_keyinput2 = ~keyinput2;
  assign new_not_0 = ~Q_0;
  assign new_and_1 = new_not_0 & Q_1;
  assign new_not_2 = ~Q_1;
  assign new_and_3 = Q_0 & new_not_2;
  assign n18703 = new_and_1 | new_and_3;
  assign n18700 = ~Q_0;
  assign new_not_Q_0 = ~Q_0;
  assign new_not_Q_1 = ~Q_1;
  assign new_count_state_1 = new_not_Q_1 & Q_0;
  assign new_count_state_2 = Q_1 & new_not_Q_0;
  assign new_count_state_3 = Q_1 & Q_0;
  assign new_y_mux_key0_and_0 = n228 & new_not_keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key0_and_1 = new_U3445 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key0 = new_y_mux_key0_and_0 | new_y_mux_key0_and_1;
  assign new_y_mux_key1_and_0 = n228 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key1_and_1 = new_U3445 & keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key1 = new_y_mux_key1_and_0 | new_y_mux_key1_and_1;
  assign new_y_mux_key2_and_0 = n228 & keyinput2 & new_not_keyinput0 & new_not_keyinput1;
  assign new_y_mux_key2_and_1 = new_U3445 & new_not_keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key2 = new_y_mux_key2_and_0 | new_y_mux_key2_and_1;
  assign new_y_mux_key3_and_0 = n228 & new_not_keyinput2 & new_not_keyinput0 & keyinput1;
  assign new_y_mux_key3_and_1 = new_U3445 & keyinput2 & keyinput0 & new_not_keyinput1;
  assign new_y_mux_key3 = new_y_mux_key3_and_0 | new_y_mux_key3_and_1;
  assign new__state_1 = new_count_state_1;
  assign new__state_2 = new_count_state_2;
  assign new__state_3 = new_count_state_3;
  assign new__state_5 = new__state_2 | new__state_3;
  assign new_s__state_1 = new__state_1;
  assign new_not_s__state_1 = ~new_s__state_1;
  assign new_I0__state_1 = new_y_mux_key0;
  assign new_I1__state_1 = new_y_mux_key1;
  assign new_and_mux__state_1 = new_not_s__state_1 & new_I0__state_1;
  assign new_and_mux__state_1_2 = new_s__state_1 & new_I1__state_1;
  assign new_y_mux_4 = new_and_mux__state_1 | new_and_mux__state_1_2;
  assign new_s__state_3 = new__state_3;
  assign new_not_s__state_3 = ~new_s__state_3;
  assign new_I0__state_3 = new_y_mux_key2;
  assign new_I1__state_3 = new_y_mux_key3;
  assign new_and_mux__state_3 = new_not_s__state_3 & new_I0__state_3;
  assign new_and_mux__state_3_2 = new_s__state_3 & new_I1__state_3;
  assign new_y_mux_5 = new_and_mux__state_3 | new_and_mux__state_3_2;
  assign new_s__state_5 = new__state_5;
  assign new_not_s__state_5 = ~new_s__state_5;
  assign new_I0__state_5 = new_y_mux_4;
  assign new_I1__state_5 = new_y_mux_5;
  assign new_and_mux__state_5 = new_not_s__state_5 & new_I0__state_5;
  assign new_and_mux__state_5_2 = new_s__state_5 & new_I1__state_5;
  assign n220 = new_and_mux__state_5 | new_and_mux__state_5_2;
  always @ (posedge clock) begin
    BE_N_REG_3_ <= n220;
    BE_N_REG_2_ <= n224;
    BE_N_REG_1_ <= n228;
    BE_N_REG_0_ <= n232;
    ADDRESS_REG_29_ <= n236;
    ADDRESS_REG_28_ <= n240;
    ADDRESS_REG_27_ <= n244;
    ADDRESS_REG_26_ <= n248;
    ADDRESS_REG_25_ <= n252;
    ADDRESS_REG_24_ <= n256;
    ADDRESS_REG_23_ <= n260;
    ADDRESS_REG_22_ <= n264;
    ADDRESS_REG_21_ <= n268;
    ADDRESS_REG_20_ <= n272;
    ADDRESS_REG_19_ <= n276;
    ADDRESS_REG_18_ <= n280;
    ADDRESS_REG_17_ <= n284;
    ADDRESS_REG_16_ <= n288;
    ADDRESS_REG_15_ <= n292;
    ADDRESS_REG_14_ <= n296;
    ADDRESS_REG_13_ <= n300;
    ADDRESS_REG_12_ <= n304;
    ADDRESS_REG_11_ <= n308;
    ADDRESS_REG_10_ <= n312;
    ADDRESS_REG_9_ <= n316;
    ADDRESS_REG_8_ <= n320;
    ADDRESS_REG_7_ <= n324;
    ADDRESS_REG_6_ <= n328;
    ADDRESS_REG_5_ <= n332;
    ADDRESS_REG_4_ <= n336;
    ADDRESS_REG_3_ <= n340;
    ADDRESS_REG_2_ <= n344;
    ADDRESS_REG_1_ <= n348;
    ADDRESS_REG_0_ <= n352;
    STATE_REG_2_ <= n356;
    STATE_REG_1_ <= n361;
    STATE_REG_0_ <= n366;
    DATAWIDTH_REG_0_ <= n371;
    DATAWIDTH_REG_1_ <= n376;
    DATAWIDTH_REG_2_ <= n381;
    DATAWIDTH_REG_3_ <= n386;
    DATAWIDTH_REG_4_ <= n391;
    DATAWIDTH_REG_5_ <= n396;
    DATAWIDTH_REG_6_ <= n401;
    DATAWIDTH_REG_7_ <= n406;
    DATAWIDTH_REG_8_ <= n411;
    DATAWIDTH_REG_9_ <= n416;
    DATAWIDTH_REG_10_ <= n421;
    DATAWIDTH_REG_11_ <= n426;
    DATAWIDTH_REG_12_ <= n431;
    DATAWIDTH_REG_13_ <= n436;
    DATAWIDTH_REG_14_ <= n441;
    DATAWIDTH_REG_15_ <= n446;
    DATAWIDTH_REG_16_ <= n451;
    DATAWIDTH_REG_17_ <= n456;
    DATAWIDTH_REG_18_ <= n461;
    DATAWIDTH_REG_19_ <= n466;
    DATAWIDTH_REG_20_ <= n471;
    DATAWIDTH_REG_21_ <= n476;
    DATAWIDTH_REG_22_ <= n481;
    DATAWIDTH_REG_23_ <= n486;
    DATAWIDTH_REG_24_ <= n491;
    DATAWIDTH_REG_25_ <= n496;
    DATAWIDTH_REG_26_ <= n501;
    DATAWIDTH_REG_27_ <= n506;
    DATAWIDTH_REG_28_ <= n511;
    DATAWIDTH_REG_29_ <= n516;
    DATAWIDTH_REG_30_ <= n521;
    DATAWIDTH_REG_31_ <= n526;
    STATE2_REG_3_ <= n531;
    STATE2_REG_2_ <= n536;
    STATE2_REG_1_ <= n541;
    STATE2_REG_0_ <= n546;
    INSTQUEUE_REG_15__7_ <= n551;
    INSTQUEUE_REG_15__6_ <= n556;
    INSTQUEUE_REG_15__5_ <= n561;
    INSTQUEUE_REG_15__4_ <= n566;
    INSTQUEUE_REG_15__3_ <= n571;
    INSTQUEUE_REG_15__2_ <= n576;
    INSTQUEUE_REG_15__1_ <= n581;
    INSTQUEUE_REG_15__0_ <= n586;
    INSTQUEUE_REG_14__7_ <= n591;
    INSTQUEUE_REG_14__6_ <= n596;
    INSTQUEUE_REG_14__5_ <= n601;
    INSTQUEUE_REG_14__4_ <= n606;
    INSTQUEUE_REG_14__3_ <= n611;
    INSTQUEUE_REG_14__2_ <= n616;
    INSTQUEUE_REG_14__1_ <= n621;
    INSTQUEUE_REG_14__0_ <= n626;
    INSTQUEUE_REG_13__7_ <= n631;
    INSTQUEUE_REG_13__6_ <= n636;
    INSTQUEUE_REG_13__5_ <= n641;
    INSTQUEUE_REG_13__4_ <= n646;
    INSTQUEUE_REG_13__3_ <= n651;
    INSTQUEUE_REG_13__2_ <= n656;
    INSTQUEUE_REG_13__1_ <= n661;
    INSTQUEUE_REG_13__0_ <= n666;
    INSTQUEUE_REG_12__7_ <= n671;
    INSTQUEUE_REG_12__6_ <= n676;
    INSTQUEUE_REG_12__5_ <= n681;
    INSTQUEUE_REG_12__4_ <= n686;
    INSTQUEUE_REG_12__3_ <= n691;
    INSTQUEUE_REG_12__2_ <= n696;
    INSTQUEUE_REG_12__1_ <= n701;
    INSTQUEUE_REG_12__0_ <= n706;
    INSTQUEUE_REG_11__7_ <= n711;
    INSTQUEUE_REG_11__6_ <= n716;
    INSTQUEUE_REG_11__5_ <= n721;
    INSTQUEUE_REG_11__4_ <= n726;
    INSTQUEUE_REG_11__3_ <= n731;
    INSTQUEUE_REG_11__2_ <= n736;
    INSTQUEUE_REG_11__1_ <= n741;
    INSTQUEUE_REG_11__0_ <= n746;
    INSTQUEUE_REG_10__7_ <= n751;
    INSTQUEUE_REG_10__6_ <= n756;
    INSTQUEUE_REG_10__5_ <= n761;
    INSTQUEUE_REG_10__4_ <= n766;
    INSTQUEUE_REG_10__3_ <= n771;
    INSTQUEUE_REG_10__2_ <= n776;
    INSTQUEUE_REG_10__1_ <= n781;
    INSTQUEUE_REG_10__0_ <= n786;
    INSTQUEUE_REG_9__7_ <= n791;
    INSTQUEUE_REG_9__6_ <= n796;
    INSTQUEUE_REG_9__5_ <= n801;
    INSTQUEUE_REG_9__4_ <= n806;
    INSTQUEUE_REG_9__3_ <= n811;
    INSTQUEUE_REG_9__2_ <= n816;
    INSTQUEUE_REG_9__1_ <= n821;
    INSTQUEUE_REG_9__0_ <= n826;
    INSTQUEUE_REG_8__7_ <= n831;
    INSTQUEUE_REG_8__6_ <= n836;
    INSTQUEUE_REG_8__5_ <= n841;
    INSTQUEUE_REG_8__4_ <= n846;
    INSTQUEUE_REG_8__3_ <= n851;
    INSTQUEUE_REG_8__2_ <= n856;
    INSTQUEUE_REG_8__1_ <= n861;
    INSTQUEUE_REG_8__0_ <= n866;
    INSTQUEUE_REG_7__7_ <= n871;
    INSTQUEUE_REG_7__6_ <= n876;
    INSTQUEUE_REG_7__5_ <= n881;
    INSTQUEUE_REG_7__4_ <= n886;
    INSTQUEUE_REG_7__3_ <= n891;
    INSTQUEUE_REG_7__2_ <= n896;
    INSTQUEUE_REG_7__1_ <= n901;
    INSTQUEUE_REG_7__0_ <= n906;
    INSTQUEUE_REG_6__7_ <= n911;
    INSTQUEUE_REG_6__6_ <= n916;
    INSTQUEUE_REG_6__5_ <= n921;
    INSTQUEUE_REG_6__4_ <= n926;
    INSTQUEUE_REG_6__3_ <= n931;
    INSTQUEUE_REG_6__2_ <= n936;
    INSTQUEUE_REG_6__1_ <= n941;
    INSTQUEUE_REG_6__0_ <= n946;
    INSTQUEUE_REG_5__7_ <= n951;
    INSTQUEUE_REG_5__6_ <= n956;
    INSTQUEUE_REG_5__5_ <= n961;
    INSTQUEUE_REG_5__4_ <= n966;
    INSTQUEUE_REG_5__3_ <= n971;
    INSTQUEUE_REG_5__2_ <= n976;
    INSTQUEUE_REG_5__1_ <= n981;
    INSTQUEUE_REG_5__0_ <= n986;
    INSTQUEUE_REG_4__7_ <= n991;
    INSTQUEUE_REG_4__6_ <= n996;
    INSTQUEUE_REG_4__5_ <= n1001;
    INSTQUEUE_REG_4__4_ <= n1006;
    INSTQUEUE_REG_4__3_ <= n1011;
    INSTQUEUE_REG_4__2_ <= n1016;
    INSTQUEUE_REG_4__1_ <= n1021;
    INSTQUEUE_REG_4__0_ <= n1026;
    INSTQUEUE_REG_3__7_ <= n1031;
    INSTQUEUE_REG_3__6_ <= n1036;
    INSTQUEUE_REG_3__5_ <= n1041;
    INSTQUEUE_REG_3__4_ <= n1046;
    INSTQUEUE_REG_3__3_ <= n1051;
    INSTQUEUE_REG_3__2_ <= n1056;
    INSTQUEUE_REG_3__1_ <= n1061;
    INSTQUEUE_REG_3__0_ <= n1066;
    INSTQUEUE_REG_2__7_ <= n1071;
    INSTQUEUE_REG_2__6_ <= n1076;
    INSTQUEUE_REG_2__5_ <= n1081;
    INSTQUEUE_REG_2__4_ <= n1086;
    INSTQUEUE_REG_2__3_ <= n1091;
    INSTQUEUE_REG_2__2_ <= n1096;
    INSTQUEUE_REG_2__1_ <= n1101;
    INSTQUEUE_REG_2__0_ <= n1106;
    INSTQUEUE_REG_1__7_ <= n1111;
    INSTQUEUE_REG_1__6_ <= n1116;
    INSTQUEUE_REG_1__5_ <= n1121;
    INSTQUEUE_REG_1__4_ <= n1126;
    INSTQUEUE_REG_1__3_ <= n1131;
    INSTQUEUE_REG_1__2_ <= n1136;
    INSTQUEUE_REG_1__1_ <= n1141;
    INSTQUEUE_REG_1__0_ <= n1146;
    INSTQUEUE_REG_0__7_ <= n1151;
    INSTQUEUE_REG_0__6_ <= n1156;
    INSTQUEUE_REG_0__5_ <= n1161;
    INSTQUEUE_REG_0__4_ <= n1166;
    INSTQUEUE_REG_0__3_ <= n1171;
    INSTQUEUE_REG_0__2_ <= n1176;
    INSTQUEUE_REG_0__1_ <= n1181;
    INSTQUEUE_REG_0__0_ <= n1186;
    INSTQUEUERD_ADDR_REG_4_ <= n1191;
    INSTQUEUERD_ADDR_REG_3_ <= n1196;
    INSTQUEUERD_ADDR_REG_2_ <= n1201;
    INSTQUEUERD_ADDR_REG_1_ <= n1206;
    INSTQUEUERD_ADDR_REG_0_ <= n1211;
    INSTQUEUEWR_ADDR_REG_4_ <= n1216;
    INSTQUEUEWR_ADDR_REG_3_ <= n1221;
    INSTQUEUEWR_ADDR_REG_2_ <= n1226;
    INSTQUEUEWR_ADDR_REG_1_ <= n1231;
    INSTQUEUEWR_ADDR_REG_0_ <= n1236;
    INSTADDRPOINTER_REG_0_ <= n1241;
    INSTADDRPOINTER_REG_1_ <= n1246;
    INSTADDRPOINTER_REG_2_ <= n1251;
    INSTADDRPOINTER_REG_3_ <= n1256;
    INSTADDRPOINTER_REG_4_ <= n1261;
    INSTADDRPOINTER_REG_5_ <= n1266;
    INSTADDRPOINTER_REG_6_ <= n1271;
    INSTADDRPOINTER_REG_7_ <= n1276;
    INSTADDRPOINTER_REG_8_ <= n1281;
    INSTADDRPOINTER_REG_9_ <= n1286;
    INSTADDRPOINTER_REG_10_ <= n1291;
    INSTADDRPOINTER_REG_11_ <= n1296;
    INSTADDRPOINTER_REG_12_ <= n1301;
    INSTADDRPOINTER_REG_13_ <= n1306;
    INSTADDRPOINTER_REG_14_ <= n1311;
    INSTADDRPOINTER_REG_15_ <= n1316;
    INSTADDRPOINTER_REG_16_ <= n1321;
    INSTADDRPOINTER_REG_17_ <= n1326;
    INSTADDRPOINTER_REG_18_ <= n1331;
    INSTADDRPOINTER_REG_19_ <= n1336;
    INSTADDRPOINTER_REG_20_ <= n1341;
    INSTADDRPOINTER_REG_21_ <= n1346;
    INSTADDRPOINTER_REG_22_ <= n1351;
    INSTADDRPOINTER_REG_23_ <= n1356;
    INSTADDRPOINTER_REG_24_ <= n1361;
    INSTADDRPOINTER_REG_25_ <= n1366;
    INSTADDRPOINTER_REG_26_ <= n1371;
    INSTADDRPOINTER_REG_27_ <= n1376;
    INSTADDRPOINTER_REG_28_ <= n1381;
    INSTADDRPOINTER_REG_29_ <= n1386;
    INSTADDRPOINTER_REG_30_ <= n1391;
    INSTADDRPOINTER_REG_31_ <= n1396;
    PHYADDRPOINTER_REG_0_ <= n1401;
    PHYADDRPOINTER_REG_1_ <= n1406;
    PHYADDRPOINTER_REG_2_ <= n1411;
    PHYADDRPOINTER_REG_3_ <= n1416;
    PHYADDRPOINTER_REG_4_ <= n1421;
    PHYADDRPOINTER_REG_5_ <= n1426;
    PHYADDRPOINTER_REG_6_ <= n1431;
    PHYADDRPOINTER_REG_7_ <= n1436;
    PHYADDRPOINTER_REG_8_ <= n1441;
    PHYADDRPOINTER_REG_9_ <= n1446;
    PHYADDRPOINTER_REG_10_ <= n1451;
    PHYADDRPOINTER_REG_11_ <= n1456;
    PHYADDRPOINTER_REG_12_ <= n1461;
    PHYADDRPOINTER_REG_13_ <= n1466;
    PHYADDRPOINTER_REG_14_ <= n1471;
    PHYADDRPOINTER_REG_15_ <= n1476;
    PHYADDRPOINTER_REG_16_ <= n1481;
    PHYADDRPOINTER_REG_17_ <= n1486;
    PHYADDRPOINTER_REG_18_ <= n1491;
    PHYADDRPOINTER_REG_19_ <= n1496;
    PHYADDRPOINTER_REG_20_ <= n1501;
    PHYADDRPOINTER_REG_21_ <= n1506;
    PHYADDRPOINTER_REG_22_ <= n1511;
    PHYADDRPOINTER_REG_23_ <= n1516;
    PHYADDRPOINTER_REG_24_ <= n1521;
    PHYADDRPOINTER_REG_25_ <= n1526;
    PHYADDRPOINTER_REG_26_ <= n1531;
    PHYADDRPOINTER_REG_27_ <= n1536;
    PHYADDRPOINTER_REG_28_ <= n1541;
    PHYADDRPOINTER_REG_29_ <= n1546;
    PHYADDRPOINTER_REG_30_ <= n1551;
    PHYADDRPOINTER_REG_31_ <= n1556;
    LWORD_REG_15_ <= n1561;
    LWORD_REG_14_ <= n1566;
    LWORD_REG_13_ <= n1571;
    LWORD_REG_12_ <= n1576;
    LWORD_REG_11_ <= n1581;
    LWORD_REG_10_ <= n1586;
    LWORD_REG_9_ <= n1591;
    LWORD_REG_8_ <= n1596;
    LWORD_REG_7_ <= n1601;
    LWORD_REG_6_ <= n1606;
    LWORD_REG_5_ <= n1611;
    LWORD_REG_4_ <= n1616;
    LWORD_REG_3_ <= n1621;
    LWORD_REG_2_ <= n1626;
    LWORD_REG_1_ <= n1631;
    LWORD_REG_0_ <= n1636;
    UWORD_REG_14_ <= n1641;
    UWORD_REG_13_ <= n1646;
    UWORD_REG_12_ <= n1651;
    UWORD_REG_11_ <= n1656;
    UWORD_REG_10_ <= n1661;
    UWORD_REG_9_ <= n1666;
    UWORD_REG_8_ <= n1671;
    UWORD_REG_7_ <= n1676;
    UWORD_REG_6_ <= n1681;
    UWORD_REG_5_ <= n1686;
    UWORD_REG_4_ <= n1691;
    UWORD_REG_3_ <= n1696;
    UWORD_REG_2_ <= n1701;
    UWORD_REG_1_ <= n1706;
    UWORD_REG_0_ <= n1711;
    DATAO_REG_0_ <= n1716;
    DATAO_REG_1_ <= n1720;
    DATAO_REG_2_ <= n1724;
    DATAO_REG_3_ <= n1728;
    DATAO_REG_4_ <= n1732;
    DATAO_REG_5_ <= n1736;
    DATAO_REG_6_ <= n1740;
    DATAO_REG_7_ <= n1744;
    DATAO_REG_8_ <= n1748;
    DATAO_REG_9_ <= n1752;
    DATAO_REG_10_ <= n1756;
    DATAO_REG_11_ <= n1760;
    DATAO_REG_12_ <= n1764;
    DATAO_REG_13_ <= n1768;
    DATAO_REG_14_ <= n1772;
    DATAO_REG_15_ <= n1776;
    DATAO_REG_16_ <= n1780;
    DATAO_REG_17_ <= n1784;
    DATAO_REG_18_ <= n1788;
    DATAO_REG_19_ <= n1792;
    DATAO_REG_20_ <= n1796;
    DATAO_REG_21_ <= n1800;
    DATAO_REG_22_ <= n1804;
    DATAO_REG_23_ <= n1808;
    DATAO_REG_24_ <= n1812;
    DATAO_REG_25_ <= n1816;
    DATAO_REG_26_ <= n1820;
    DATAO_REG_27_ <= n1824;
    DATAO_REG_28_ <= n1828;
    DATAO_REG_29_ <= n1832;
    DATAO_REG_30_ <= n1836;
    DATAO_REG_31_ <= n1840;
    EAX_REG_0_ <= n1844;
    EAX_REG_1_ <= n1849;
    EAX_REG_2_ <= n1854;
    EAX_REG_3_ <= n1859;
    EAX_REG_4_ <= n1864;
    EAX_REG_5_ <= n1869;
    EAX_REG_6_ <= n1874;
    EAX_REG_7_ <= n1879;
    EAX_REG_8_ <= n1884;
    EAX_REG_9_ <= n1889;
    EAX_REG_10_ <= n1894;
    EAX_REG_11_ <= n1899;
    EAX_REG_12_ <= n1904;
    EAX_REG_13_ <= n1909;
    EAX_REG_14_ <= n1914;
    EAX_REG_15_ <= n1919;
    EAX_REG_16_ <= n1924;
    EAX_REG_17_ <= n1929;
    EAX_REG_18_ <= n1934;
    EAX_REG_19_ <= n1939;
    EAX_REG_20_ <= n1944;
    EAX_REG_21_ <= n1949;
    EAX_REG_22_ <= n1954;
    EAX_REG_23_ <= n1959;
    EAX_REG_24_ <= n1964;
    EAX_REG_25_ <= n1969;
    EAX_REG_26_ <= n1974;
    EAX_REG_27_ <= n1979;
    EAX_REG_28_ <= n1984;
    EAX_REG_29_ <= n1989;
    EAX_REG_30_ <= n1994;
    EAX_REG_31_ <= n1999;
    EBX_REG_0_ <= n2004;
    EBX_REG_1_ <= n2009;
    EBX_REG_2_ <= n2014;
    EBX_REG_3_ <= n2019;
    EBX_REG_4_ <= n2024;
    EBX_REG_5_ <= n2029;
    EBX_REG_6_ <= n2034;
    EBX_REG_7_ <= n2039;
    EBX_REG_8_ <= n2044;
    EBX_REG_9_ <= n2049;
    EBX_REG_10_ <= n2054;
    EBX_REG_11_ <= n2059;
    EBX_REG_12_ <= n2064;
    EBX_REG_13_ <= n2069;
    EBX_REG_14_ <= n2074;
    EBX_REG_15_ <= n2079;
    EBX_REG_16_ <= n2084;
    EBX_REG_17_ <= n2089;
    EBX_REG_18_ <= n2094;
    EBX_REG_19_ <= n2099;
    EBX_REG_20_ <= n2104;
    EBX_REG_21_ <= n2109;
    EBX_REG_22_ <= n2114;
    EBX_REG_23_ <= n2119;
    EBX_REG_24_ <= n2124;
    EBX_REG_25_ <= n2129;
    EBX_REG_26_ <= n2134;
    EBX_REG_27_ <= n2139;
    EBX_REG_28_ <= n2144;
    EBX_REG_29_ <= n2149;
    EBX_REG_30_ <= n2154;
    EBX_REG_31_ <= n2159;
    REIP_REG_0_ <= n2164;
    REIP_REG_1_ <= n2169;
    REIP_REG_2_ <= n2174;
    REIP_REG_3_ <= n2179;
    REIP_REG_4_ <= n2184;
    REIP_REG_5_ <= n2189;
    REIP_REG_6_ <= n2194;
    REIP_REG_7_ <= n2199;
    REIP_REG_8_ <= n2204;
    REIP_REG_9_ <= n2209;
    REIP_REG_10_ <= n2214;
    REIP_REG_11_ <= n2219;
    REIP_REG_12_ <= n2224;
    REIP_REG_13_ <= n2229;
    REIP_REG_14_ <= n2234;
    REIP_REG_15_ <= n2239;
    REIP_REG_16_ <= n2244;
    REIP_REG_17_ <= n2249;
    REIP_REG_18_ <= n2254;
    REIP_REG_19_ <= n2259;
    REIP_REG_20_ <= n2264;
    REIP_REG_21_ <= n2269;
    REIP_REG_22_ <= n2274;
    REIP_REG_23_ <= n2279;
    REIP_REG_24_ <= n2284;
    REIP_REG_25_ <= n2289;
    REIP_REG_26_ <= n2294;
    REIP_REG_27_ <= n2299;
    REIP_REG_28_ <= n2304;
    REIP_REG_29_ <= n2309;
    REIP_REG_30_ <= n2314;
    REIP_REG_31_ <= n2319;
    BYTEENABLE_REG_3_ <= n2324;
    BYTEENABLE_REG_2_ <= n2329;
    BYTEENABLE_REG_1_ <= n2334;
    BYTEENABLE_REG_0_ <= n2339;
    W_R_N_REG <= n2344;
    FLUSH_REG <= n2348;
    MORE_REG <= n2353;
    STATEBS16_REG <= n2358;
    REQUESTPENDING_REG <= n2363;
    D_C_N_REG <= n2368;
    M_IO_N_REG <= n2372;
    CODEFETCH_REG <= n2376;
    ADS_N_REG <= n2381;
    READREQUEST_REG <= n2385;
    MEMORYFETCH_REG <= n2390;
    Q_0 <= n18700;
    Q_1 <= n18703;
  end
endmodule
