library ieee;
use ieee.std_logic_1164.all;

entity cyr is
   port ( clk,rst,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,
	x16,x17,x18,x19,x20 : in std_logic;
        y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,
	y16,y17,y18,y19,y20,y21,y22,y23,y24,y25,y26,y27,y28,y29,y30,
	y31,y32,y33,y34,y35,y36,y37,y38,y39,y40,y41,y42,y43,y44,y45,
	y46,y47,y48,y49,y50,y51,y52,y53,y54,y55,y56,y57,y58,y59,y60,
	y61,y62,y63,y64,y65,y66,y67,y68,y69,y70,y71,y72,y73,y74,y75
	 : out std_logic );
end cyr;

architecture ARC of cyr is

   type states_cyr is ( s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,
	s16,s17,s18,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29,s30,
	s31,s32,s33,s34,s35,s36,s37,s38,s39,s40,s41,s42 );
   signal current_cyr : states_cyr;

begin
   process (clk , rst)
   procedure proc_cyr is
   begin

	y1   <= '0' ;	y2   <= '0' ;	y3   <= '0' ;	y4   <= '0' ;
	y5   <= '0' ;	y6   <= '0' ;	y7   <= '0' ;	y8   <= '0' ;
	y9   <= '0' ;	y10  <= '0' ;	y11  <= '0' ;	y12  <= '0' ;
	y13  <= '0' ;	y14  <= '0' ;	y15  <= '0' ;	y16  <= '0' ;
	y17  <= '0' ;	y18  <= '0' ;	y19  <= '0' ;	y20  <= '0' ;
	y21  <= '0' ;	y22  <= '0' ;	y23  <= '0' ;	y24  <= '0' ;
	y25  <= '0' ;	y26  <= '0' ;	y27  <= '0' ;	y28  <= '0' ;
	y29  <= '0' ;	y30  <= '0' ;	y31  <= '0' ;	y32  <= '0' ;
	y33  <= '0' ;	y34  <= '0' ;	y35  <= '0' ;	y36  <= '0' ;
	y37  <= '0' ;	y38  <= '0' ;	y39  <= '0' ;	y40  <= '0' ;
	y41  <= '0' ;	y42  <= '0' ;	y43  <= '0' ;	y44  <= '0' ;
	y45  <= '0' ;	y46  <= '0' ;	y47  <= '0' ;	y48  <= '0' ;
	y49  <= '0' ;	y50  <= '0' ;	y51  <= '0' ;	y52  <= '0' ;
	y53  <= '0' ;	y54  <= '0' ;	y55  <= '0' ;	y56  <= '0' ;
	y57  <= '0' ;	y58  <= '0' ;	y59  <= '0' ;	y60  <= '0' ;
	y61  <= '0' ;	y62  <= '0' ;	y63  <= '0' ;	y64  <= '0' ;
	y65  <= '0' ;	y66  <= '0' ;	y67  <= '0' ;	y68  <= '0' ;
	y69  <= '0' ;	y70  <= '0' ;	y71  <= '0' ;	y72  <= '0' ;
	y73  <= '0' ;	y74  <= '0' ;	y75  <= '0' ;

   case current_cyr is
   when s1 =>
      if ( x1 and x2 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_cyr <= s2;

      elsif ( x1 and not x2 ) = '1' then
         y1 <= '1' ;
         current_cyr <= s3;

      else
         current_cyr <= s1;

      end if;

   when s2 =>
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_cyr <= s4;

   when s3 =>
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_cyr <= s5;

   when s4 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y69 <= '1' ;
         y70 <= '1' ;
         y71 <= '1' ;
         current_cyr <= s6;

   when s5 =>
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         y68 <= '1' ;
         current_cyr <= s7;

   when s6 =>
         y58 <= '1' ;
         current_cyr <= s8;

   when s7 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_cyr <= s9;

   when s8 =>
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_cyr <= s10;

   when s9 =>
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_cyr <= s11;

   when s10 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_cyr <= s12;

   when s11 =>
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         y68 <= '1' ;
         current_cyr <= s13;

   when s12 =>
         y23 <= '1' ;
         y72 <= '1' ;
         y73 <= '1' ;
         current_cyr <= s1;

   when s13 =>
         y9 <= '1' ;
         current_cyr <= s14;

   when s14 =>
      if ( x3 and x5 and x6 and x7 and x9 ) = '1' then
         y21 <= '1' ;
         current_cyr <= s15;

      elsif ( x3 and x5 and x6 and x7 and not x9 ) = '1' then
         y75 <= '1' ;
         current_cyr <= s15;

      elsif ( x3 and x5 and x6 and not x7 and x8 and x9 and x12 ) = '1' then
         y23 <= '1' ;
         current_cyr <= s15;

      elsif ( x3 and x5 and x6 and not x7 and x8 and x9 and not x12 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( x3 and x5 and x6 and not x7 and x8 and x9 and not x12 and x20 and not x13 ) = '1' then
         current_cyr <= s1;

      elsif ( x3 and x5 and x6 and not x7 and x8 and x9 and not x12 and not x20 ) = '1' then
         current_cyr <= s1;

      elsif ( x3 and x5 and x6 and not x7 and x8 and not x9 and x13 ) = '1' then
         y23 <= '1' ;
         current_cyr <= s15;

      elsif ( x3 and x5 and x6 and not x7 and x8 and not x9 and not x13 and x20 and x12 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( x3 and x5 and x6 and not x7 and x8 and not x9 and not x13 and x20 and not x12 ) = '1' then
         current_cyr <= s1;

      elsif ( x3 and x5 and x6 and not x7 and x8 and not x9 and not x13 and not x20 ) = '1' then
         current_cyr <= s1;

      elsif ( x3 and x5 and x6 and not x7 and not x8 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         y26 <= '1' ;
         current_cyr <= s15;

      elsif ( x3 and x5 and x6 and not x7 and not x8 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         y29 <= '1' ;
         current_cyr <= s15;

      elsif ( x3 and x5 and not x6 and x11 and x7 and x8 and x9 ) = '1' then
         y47 <= '1' ;
         current_cyr <= s15;

      elsif ( x3 and x5 and not x6 and x11 and x7 and x8 and not x9 ) = '1' then
         y48 <= '1' ;
         current_cyr <= s15;

      elsif ( x3 and x5 and not x6 and x11 and x7 and not x8 and x9 ) = '1' then
         y49 <= '1' ;
         current_cyr <= s15;

      elsif ( x3 and x5 and not x6 and x11 and x7 and not x8 and not x9 ) = '1' then
         y50 <= '1' ;
         current_cyr <= s15;

      elsif ( x3 and x5 and not x6 and x11 and not x7 and x8 and x9 ) = '1' then
         y51 <= '1' ;
         current_cyr <= s16;

      elsif ( x3 and x5 and not x6 and x11 and not x7 and x8 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y28 <= '1' ;
         current_cyr <= s17;

      elsif ( x3 and x5 and not x6 and x11 and not x7 and not x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y55 <= '1' ;
         current_cyr <= s15;

      elsif ( x3 and x5 and not x6 and not x11 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y41 <= '1' ;
         current_cyr <= s19;

      elsif ( x3 and not x5 and x6 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y41 <= '1' ;
         current_cyr <= s19;

      elsif ( x3 and not x5 and not x6 and x11 and x8 and x9 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_cyr <= s15;

      elsif ( x3 and not x5 and not x6 and x11 and x8 and not x9 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_cyr <= s15;

      elsif ( x3 and not x5 and not x6 and x11 and not x8 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_cyr <= s15;

      elsif ( x3 and not x5 and not x6 and not x11 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y41 <= '1' ;
         current_cyr <= s19;

      else
         y5 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_cyr <= s21;

      end if;

   when s15 =>
      if ( x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( x20 and not x13 and not x12 ) = '1' then
         current_cyr <= s1;

      else
         current_cyr <= s1;

      end if;

   when s16 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y24 <= '1' ;
         current_cyr <= s22;

   when s17 =>
         y57 <= '1' ;
         current_cyr <= s23;

   when s18 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y54 <= '1' ;
         current_cyr <= s24;

   when s19 =>
      if ( x10 ) = '1' then
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_cyr <= s25;

      elsif ( not x10 and x14 and x6 and x7 and x8 ) = '1' then
         y63 <= '1' ;
         current_cyr <= s26;

      elsif ( not x10 and x14 and x6 and x7 and not x8 and x9 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y74 <= '1' ;
         current_cyr <= s27;

      elsif ( not x10 and x14 and x6 and x7 and not x8 and not x9 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_cyr <= s15;

      elsif ( not x10 and x14 and x6 and x7 and not x8 and not x9 and not x17 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( not x10 and x14 and x6 and x7 and not x8 and not x9 and not x17 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( not x10 and x14 and x6 and x7 and not x8 and not x9 and not x17 and x20 and not x13 and not x12 ) = '1' then
         current_cyr <= s1;

      elsif ( not x10 and x14 and x6 and x7 and not x8 and not x9 and not x17 and not x20 ) = '1' then
         current_cyr <= s1;

      elsif ( not x10 and x14 and x6 and not x7 and x8 and x9 and x18 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_cyr <= s15;

      elsif ( not x10 and x14 and x6 and not x7 and x8 and x9 and not x18 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( not x10 and x14 and x6 and not x7 and x8 and x9 and not x18 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( not x10 and x14 and x6 and not x7 and x8 and x9 and not x18 and x20 and not x13 and not x12 ) = '1' then
         current_cyr <= s1;

      elsif ( not x10 and x14 and x6 and not x7 and x8 and x9 and not x18 and not x20 ) = '1' then
         current_cyr <= s1;

      elsif ( not x10 and x14 and x6 and not x7 and x8 and not x9 and x19 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_cyr <= s15;

      elsif ( not x10 and x14 and x6 and not x7 and x8 and not x9 and not x19 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( not x10 and x14 and x6 and not x7 and x8 and not x9 and not x19 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( not x10 and x14 and x6 and not x7 and x8 and not x9 and not x19 and x20 and not x13 and not x12 ) = '1' then
         current_cyr <= s1;

      elsif ( not x10 and x14 and x6 and not x7 and x8 and not x9 and not x19 and not x20 ) = '1' then
         current_cyr <= s1;

      elsif ( not x10 and x14 and x6 and not x7 and not x8 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_cyr <= s15;

      elsif ( not x10 and x14 and x6 and not x7 and not x8 and not x9 ) = '1' then
         y65 <= '1' ;
         current_cyr <= s15;

      elsif ( not x10 and x14 and not x6 ) = '1' then
         y57 <= '1' ;
         current_cyr <= s28;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y40 <= '1' ;
         y45 <= '1' ;
         current_cyr <= s20;

      end if;

   when s20 =>
      if ( x6 and x7 and x8 ) = '1' then
         y63 <= '1' ;
         current_cyr <= s26;

      elsif ( x6 and x7 and not x8 and x9 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y74 <= '1' ;
         current_cyr <= s27;

      elsif ( x6 and x7 and not x8 and not x9 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_cyr <= s15;

      elsif ( x6 and x7 and not x8 and not x9 and not x17 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( x6 and x7 and not x8 and not x9 and not x17 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( x6 and x7 and not x8 and not x9 and not x17 and x20 and not x13 and not x12 ) = '1' then
         current_cyr <= s1;

      elsif ( x6 and x7 and not x8 and not x9 and not x17 and not x20 ) = '1' then
         current_cyr <= s1;

      elsif ( x6 and not x7 and x8 and x9 and x18 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_cyr <= s15;

      elsif ( x6 and not x7 and x8 and x9 and not x18 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( x6 and not x7 and x8 and x9 and not x18 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( x6 and not x7 and x8 and x9 and not x18 and x20 and not x13 and not x12 ) = '1' then
         current_cyr <= s1;

      elsif ( x6 and not x7 and x8 and x9 and not x18 and not x20 ) = '1' then
         current_cyr <= s1;

      elsif ( x6 and not x7 and x8 and not x9 and x19 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_cyr <= s15;

      elsif ( x6 and not x7 and x8 and not x9 and not x19 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( x6 and not x7 and x8 and not x9 and not x19 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( x6 and not x7 and x8 and not x9 and not x19 and x20 and not x13 and not x12 ) = '1' then
         current_cyr <= s1;

      elsif ( x6 and not x7 and x8 and not x9 and not x19 and not x20 ) = '1' then
         current_cyr <= s1;

      elsif ( x6 and not x7 and not x8 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_cyr <= s15;

      elsif ( x6 and not x7 and not x8 and not x9 ) = '1' then
         y65 <= '1' ;
         current_cyr <= s15;

      else
         y57 <= '1' ;
         current_cyr <= s28;

      end if;

   when s21 =>
      if ( x4 ) = '1' then
         y67 <= '1' ;
         current_cyr <= s3;

      elsif ( not x4 and x5 and x6 and x7 and x9 ) = '1' then
         y21 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and x5 and x6 and x7 and not x9 ) = '1' then
         y75 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and x5 and x6 and not x7 and x8 and x9 and x12 ) = '1' then
         y23 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and x5 and x6 and not x7 and x8 and x9 and not x12 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( not x4 and x5 and x6 and not x7 and x8 and x9 and not x12 and x20 and not x13 ) = '1' then
         current_cyr <= s1;

      elsif ( not x4 and x5 and x6 and not x7 and x8 and x9 and not x12 and not x20 ) = '1' then
         current_cyr <= s1;

      elsif ( not x4 and x5 and x6 and not x7 and x8 and not x9 and x13 ) = '1' then
         y23 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and x5 and x6 and not x7 and x8 and not x9 and not x13 and x20 and x12 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( not x4 and x5 and x6 and not x7 and x8 and not x9 and not x13 and x20 and not x12 ) = '1' then
         current_cyr <= s1;

      elsif ( not x4 and x5 and x6 and not x7 and x8 and not x9 and not x13 and not x20 ) = '1' then
         current_cyr <= s1;

      elsif ( not x4 and x5 and x6 and not x7 and not x8 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y24 <= '1' ;
         y25 <= '1' ;
         y26 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and x5 and x6 and not x7 and not x8 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y27 <= '1' ;
         y28 <= '1' ;
         y29 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and x5 and not x6 and x3 and x11 and x7 and x8 and x9 ) = '1' then
         y47 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and x5 and not x6 and x3 and x11 and x7 and x8 and not x9 ) = '1' then
         y48 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and x5 and not x6 and x3 and x11 and x7 and not x8 and x9 ) = '1' then
         y49 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and x5 and not x6 and x3 and x11 and x7 and not x8 and not x9 ) = '1' then
         y50 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and x5 and not x6 and x3 and x11 and not x7 and x8 and x9 ) = '1' then
         y51 <= '1' ;
         current_cyr <= s16;

      elsif ( not x4 and x5 and not x6 and x3 and x11 and not x7 and x8 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y28 <= '1' ;
         current_cyr <= s17;

      elsif ( not x4 and x5 and not x6 and x3 and x11 and not x7 and not x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y55 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and x5 and not x6 and x3 and not x11 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y41 <= '1' ;
         current_cyr <= s19;

      elsif ( not x4 and x5 and not x6 and not x3 and x10 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y46 <= '1' ;
         current_cyr <= s20;

      elsif ( not x4 and x5 and not x6 and not x3 and not x10 and x7 and x8 and x9 ) = '1' then
         y47 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and x5 and not x6 and not x3 and not x10 and x7 and x8 and not x9 ) = '1' then
         y48 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and x5 and not x6 and not x3 and not x10 and x7 and not x8 and x9 ) = '1' then
         y49 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and x5 and not x6 and not x3 and not x10 and x7 and not x8 and not x9 ) = '1' then
         y50 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and x5 and not x6 and not x3 and not x10 and not x7 and x8 and x9 ) = '1' then
         y51 <= '1' ;
         current_cyr <= s18;

      elsif ( not x4 and x5 and not x6 and not x3 and not x10 and not x7 and x8 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y53 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and x5 and not x6 and not x3 and not x10 and not x7 and not x8 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y54 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and x5 and not x6 and not x3 and not x10 and not x7 and not x8 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and not x5 and x6 and x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y41 <= '1' ;
         current_cyr <= s19;

      elsif ( not x4 and not x5 and x6 and not x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y46 <= '1' ;
         current_cyr <= s20;

      elsif ( not x4 and not x5 and not x6 and x3 and x11 and x8 and x9 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and not x5 and not x6 and x3 and x11 and x8 and not x9 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and not x5 and not x6 and x3 and x11 and not x8 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and not x5 and not x6 and x3 and not x11 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y41 <= '1' ;
         current_cyr <= s19;

      elsif ( not x4 and not x5 and not x6 and not x3 and x10 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y46 <= '1' ;
         current_cyr <= s20;

      elsif ( not x4 and not x5 and not x6 and not x3 and not x10 and x7 and x8 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and not x5 and not x6 and not x3 and not x10 and x7 and x8 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and not x5 and not x6 and not x3 and not x10 and x7 and not x8 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y30 <= '1' ;
         y31 <= '1' ;
         y38 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and not x5 and not x6 and not x3 and not x10 and x7 and not x8 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         y39 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and not x5 and not x6 and not x3 and not x10 and not x7 and x8 and x9 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y40 <= '1' ;
         current_cyr <= s15;

      elsif ( not x4 and not x5 and not x6 and not x3 and not x10 and not x7 and x8 and not x9 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y40 <= '1' ;
         current_cyr <= s15;

      else
         y5 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         y40 <= '1' ;
         current_cyr <= s15;

      end if;

   when s22 =>
         y56 <= '1' ;
         current_cyr <= s17;

   when s23 =>
         y58 <= '1' ;
         current_cyr <= s29;

   when s24 =>
         y52 <= '1' ;
         current_cyr <= s15;

   when s25 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         y60 <= '1' ;
         y61 <= '1' ;
         y62 <= '1' ;
         current_cyr <= s30;

   when s26 =>
      if ( x16 ) = '1' then
         y23 <= '1' ;
         current_cyr <= s15;

      elsif ( not x16 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( not x16 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( not x16 and x20 and not x13 and not x12 ) = '1' then
         current_cyr <= s1;

      else
         current_cyr <= s1;

      end if;

   when s27 =>
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_cyr <= s31;

   when s28 =>
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_cyr <= s32;

   when s29 =>
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_cyr <= s33;

   when s30 =>
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_cyr <= s34;

   when s31 =>
         y33 <= '1' ;
         current_cyr <= s35;

   when s32 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y33 <= '1' ;
         y59 <= '1' ;
         y60 <= '1' ;
         y61 <= '1' ;
         y62 <= '1' ;
         current_cyr <= s36;

   when s33 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y59 <= '1' ;
         y69 <= '1' ;
         y70 <= '1' ;
         y71 <= '1' ;
         current_cyr <= s37;

   when s34 =>
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y74 <= '1' ;
         current_cyr <= s38;

   when s35 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y69 <= '1' ;
         y70 <= '1' ;
         y71 <= '1' ;
         current_cyr <= s39;

   when s36 =>
      if ( x15 ) = '1' then
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_cyr <= s40;

      else
         y5 <= '1' ;
         y42 <= '1' ;
         y43 <= '1' ;
         y44 <= '1' ;
         current_cyr <= s32;

      end if;

   when s37 =>
      if ( x15 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_cyr <= s15;

      else
         y58 <= '1' ;
         current_cyr <= s29;

      end if;

   when s38 =>
      if ( x14 and x6 and x7 and x8 ) = '1' then
         y63 <= '1' ;
         current_cyr <= s26;

      elsif ( x14 and x6 and x7 and not x8 and x9 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         y74 <= '1' ;
         current_cyr <= s27;

      elsif ( x14 and x6 and x7 and not x8 and not x9 and x17 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_cyr <= s15;

      elsif ( x14 and x6 and x7 and not x8 and not x9 and not x17 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( x14 and x6 and x7 and not x8 and not x9 and not x17 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( x14 and x6 and x7 and not x8 and not x9 and not x17 and x20 and not x13 and not x12 ) = '1' then
         current_cyr <= s1;

      elsif ( x14 and x6 and x7 and not x8 and not x9 and not x17 and not x20 ) = '1' then
         current_cyr <= s1;

      elsif ( x14 and x6 and not x7 and x8 and x9 and x18 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_cyr <= s15;

      elsif ( x14 and x6 and not x7 and x8 and x9 and not x18 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( x14 and x6 and not x7 and x8 and x9 and not x18 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( x14 and x6 and not x7 and x8 and x9 and not x18 and x20 and not x13 and not x12 ) = '1' then
         current_cyr <= s1;

      elsif ( x14 and x6 and not x7 and x8 and x9 and not x18 and not x20 ) = '1' then
         current_cyr <= s1;

      elsif ( x14 and x6 and not x7 and x8 and not x9 and x19 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_cyr <= s15;

      elsif ( x14 and x6 and not x7 and x8 and not x9 and not x19 and x20 and x13 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( x14 and x6 and not x7 and x8 and not x9 and not x19 and x20 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_cyr <= s1;

      elsif ( x14 and x6 and not x7 and x8 and not x9 and not x19 and x20 and not x13 and not x12 ) = '1' then
         current_cyr <= s1;

      elsif ( x14 and x6 and not x7 and x8 and not x9 and not x19 and not x20 ) = '1' then
         current_cyr <= s1;

      elsif ( x14 and x6 and not x7 and not x8 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_cyr <= s15;

      elsif ( x14 and x6 and not x7 and not x8 and not x9 ) = '1' then
         y65 <= '1' ;
         current_cyr <= s15;

      elsif ( x14 and not x6 ) = '1' then
         y57 <= '1' ;
         current_cyr <= s28;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y20 <= '1' ;
         y40 <= '1' ;
         y45 <= '1' ;
         current_cyr <= s20;

      end if;

   when s39 =>
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_cyr <= s41;

   when s40 =>
      if ( x5 and x7 and x8 and x9 ) = '1' then
         y47 <= '1' ;
         current_cyr <= s15;

      elsif ( x5 and x7 and x8 and not x9 ) = '1' then
         y48 <= '1' ;
         current_cyr <= s15;

      elsif ( x5 and x7 and not x8 and x9 ) = '1' then
         y49 <= '1' ;
         current_cyr <= s15;

      elsif ( x5 and x7 and not x8 and not x9 ) = '1' then
         y50 <= '1' ;
         current_cyr <= s15;

      elsif ( x5 and not x7 and x3 and x8 and x9 ) = '1' then
         y51 <= '1' ;
         current_cyr <= s16;

      elsif ( x5 and not x7 and x3 and x8 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y28 <= '1' ;
         current_cyr <= s17;

      elsif ( x5 and not x7 and x3 and not x8 and x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y55 <= '1' ;
         current_cyr <= s15;

      elsif ( x5 and not x7 and x3 and not x8 and not x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y24 <= '1' ;
         current_cyr <= s15;

      elsif ( x5 and not x7 and not x3 and x8 and x10 and x9 ) = '1' then
         y51 <= '1' ;
         current_cyr <= s16;

      elsif ( x5 and not x7 and not x3 and x8 and x10 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y28 <= '1' ;
         current_cyr <= s17;

      elsif ( x5 and not x7 and not x3 and x8 and not x10 and x9 ) = '1' then
         y51 <= '1' ;
         current_cyr <= s18;

      elsif ( x5 and not x7 and not x3 and x8 and not x10 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y16 <= '1' ;
         y53 <= '1' ;
         current_cyr <= s15;

      elsif ( x5 and not x7 and not x3 and not x8 and x9 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y24 <= '1' ;
         current_cyr <= s15;

      elsif ( x5 and not x7 and not x3 and not x8 and x9 and not x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         y54 <= '1' ;
         current_cyr <= s15;

      elsif ( x5 and not x7 and not x3 and not x8 and not x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         current_cyr <= s15;

      elsif ( not x5 and x8 and x9 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y66 <= '1' ;
         current_cyr <= s15;

      elsif ( not x5 and x8 and not x9 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y66 <= '1' ;
         current_cyr <= s15;

      else
         y5 <= '1' ;
         y16 <= '1' ;
         y18 <= '1' ;
         y20 <= '1' ;
         y66 <= '1' ;
         current_cyr <= s15;

      end if;

   when s41 =>
         y33 <= '1' ;
         current_cyr <= s42;

   when s42 =>
         y3 <= '1' ;
         y5 <= '1' ;
         y45 <= '1' ;
         y64 <= '1' ;
         current_cyr <= s15;

   end case;
   end proc_cyr;

   begin
      if ( rst = '1' ) then
	y1   <= '0' ;	y2   <= '0' ;	y3   <= '0' ;	y4   <= '0' ;
	y5   <= '0' ;	y6   <= '0' ;	y7   <= '0' ;	y8   <= '0' ;
	y9   <= '0' ;	y10  <= '0' ;	y11  <= '0' ;	y12  <= '0' ;
	y13  <= '0' ;	y14  <= '0' ;	y15  <= '0' ;	y16  <= '0' ;
	y17  <= '0' ;	y18  <= '0' ;	y19  <= '0' ;	y20  <= '0' ;
	y21  <= '0' ;	y22  <= '0' ;	y23  <= '0' ;	y24  <= '0' ;
	y25  <= '0' ;	y26  <= '0' ;	y27  <= '0' ;	y28  <= '0' ;
	y29  <= '0' ;	y30  <= '0' ;	y31  <= '0' ;	y32  <= '0' ;
	y33  <= '0' ;	y34  <= '0' ;	y35  <= '0' ;	y36  <= '0' ;
	y37  <= '0' ;	y38  <= '0' ;	y39  <= '0' ;	y40  <= '0' ;
	y41  <= '0' ;	y42  <= '0' ;	y43  <= '0' ;	y44  <= '0' ;
	y45  <= '0' ;	y46  <= '0' ;	y47  <= '0' ;	y48  <= '0' ;
	y49  <= '0' ;	y50  <= '0' ;	y51  <= '0' ;	y52  <= '0' ;
	y53  <= '0' ;	y54  <= '0' ;	y55  <= '0' ;	y56  <= '0' ;
	y57  <= '0' ;	y58  <= '0' ;	y59  <= '0' ;	y60  <= '0' ;
	y61  <= '0' ;	y62  <= '0' ;	y63  <= '0' ;	y64  <= '0' ;
	y65  <= '0' ;	y66  <= '0' ;	y67  <= '0' ;	y68  <= '0' ;
	y69  <= '0' ;	y70  <= '0' ;	y71  <= '0' ;	y72  <= '0' ;
	y73  <= '0' ;	y74  <= '0' ;	y75  <= '0' ;
	current_cyr <= s1;
      elsif (clk'event and clk ='1') then
        proc_cyr;
      end if;
   end process;
end ARC;
