library ieee;
use ieee.std_logic_1164.all;

entity pp is
   port ( clk,rst,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,
	x16,x17,x18,x19,x20 : in std_logic;
        y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,
	y16,y17,y18,y19,y20,y21,y22,y23,y24,y25,y26,y27,y28 : out std_logic );
end pp;

architecture ARC of pp is

   type states_pp is ( s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,
	s16,s17 );
   signal current_pp : states_pp;

begin
   process (clk , rst)
   procedure proc_pp is
   begin

	y1   <= '0' ;	y2   <= '0' ;	y3   <= '0' ;	y4   <= '0' ;
	y5   <= '0' ;	y6   <= '0' ;	y7   <= '0' ;	y8   <= '0' ;
	y9   <= '0' ;	y10  <= '0' ;	y11  <= '0' ;	y12  <= '0' ;
	y13  <= '0' ;	y14  <= '0' ;	y15  <= '0' ;	y16  <= '0' ;
	y17  <= '0' ;	y18  <= '0' ;	y19  <= '0' ;	y20  <= '0' ;
	y21  <= '0' ;	y22  <= '0' ;	y23  <= '0' ;	y24  <= '0' ;
	y25  <= '0' ;	y26  <= '0' ;	y27  <= '0' ;	y28  <= '0' ;


   case current_pp is
   when s1 =>
      if ( x13 and x1 and x10 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_pp <= s2;

      elsif ( x13 and x1 and not x10 and x2 and x3 and x15 ) = '1' then
         current_pp <= s1;

      elsif ( x13 and x1 and not x10 and x2 and x3 and not x15 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_pp <= s3;

      elsif ( x13 and x1 and not x10 and x2 and not x3 and x4 and x5 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_pp <= s4;

      elsif ( x13 and x1 and not x10 and x2 and not x3 and x4 and not x5 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_pp <= s5;

      elsif ( x13 and x1 and not x10 and x2 and not x3 and not x4 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_pp <= s2;

      elsif ( x13 and x1 and not x10 and not x2 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_pp <= s6;

      elsif ( x13 and not x1 and x10 and x2 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s7;

      elsif ( x13 and not x1 and x10 and not x2 and x15 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s7;

      elsif ( x13 and not x1 and x10 and not x2 and not x15 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_pp <= s3;

      elsif ( x13 and not x1 and not x10 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s7;

      elsif ( not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_pp <= s6;

      elsif ( not x13 and not x12 and x10 and x1 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_pp <= s2;

      elsif ( not x13 and not x12 and x10 and not x1 and x4 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s7;

      elsif ( not x13 and not x12 and x10 and not x1 and not x4 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_pp <= s3;

      else
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_pp <= s6;

      end if;

   when s2 =>
      if ( x13 and x10 and x3 and x5 ) = '1' then
         y2 <= '1' ;
         y20 <= '1' ;
         y25 <= '1' ;
         current_pp <= s8;

      elsif ( x13 and x10 and x3 and not x5 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_pp <= s9;

      elsif ( x13 and x10 and not x3 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_pp <= s4;

      elsif ( x13 and not x10 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_pp <= s5;

      elsif ( not x13 and x12 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_pp <= s3;

      elsif ( not x13 and not x12 and x5 and x10 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s7;

      elsif ( not x13 and not x12 and x5 and not x10 and x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_pp <= s10;

      elsif ( not x13 and not x12 and x5 and not x10 and not x3 and x4 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s11;

      elsif ( not x13 and not x12 and x5 and not x10 and not x3 and not x4 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_pp <= s9;

      elsif ( not x13 and not x12 and not x5 and x10 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_pp <= s9;

      else
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_pp <= s5;

      end if;

   when s3 =>
      if ( x13 and x10 and x9 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_pp <= s5;

      elsif ( x13 and x10 and not x9 and x17 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s7;

      elsif ( x13 and x10 and not x9 and not x17 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_pp <= s3;

      elsif ( x13 and not x10 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_pp <= s4;

      elsif ( not x13 and x12 and x4 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_pp <= s4;

      elsif ( not x13 and x12 and not x4 ) = '1' then
         current_pp <= s1;

      elsif ( not x13 and not x12 and x10 and x2 and x16 ) = '1' then
         y2 <= '1' ;
         y20 <= '1' ;
         y25 <= '1' ;
         current_pp <= s8;

      elsif ( not x13 and not x12 and x10 and x2 and not x16 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_pp <= s9;

      elsif ( not x13 and not x12 and x10 and not x2 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_pp <= s4;

      elsif ( not x13 and not x12 and not x10 and x18 and x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_pp <= s10;

      elsif ( not x13 and not x12 and not x10 and x18 and not x3 and x4 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s11;

      elsif ( not x13 and not x12 and not x10 and x18 and not x3 and not x4 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_pp <= s9;

      else
         y11 <= '1' ;
         y18 <= '1' ;
         current_pp <= s4;

      end if;

   when s4 =>
      if ( x13 and x10 and x6 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_pp <= s2;

      elsif ( x13 and x10 and not x6 and x4 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s7;

      elsif ( x13 and x10 and not x6 and not x4 ) = '1' then
         current_pp <= s1;

      elsif ( x13 and not x10 ) = '1' then
         current_pp <= s1;

      elsif ( not x13 and x12 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_pp <= s9;

      elsif ( not x13 and not x12 and x10 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_pp <= s12;

      else
         y11 <= '1' ;
         y23 <= '1' ;
         current_pp <= s9;

      end if;

   when s5 =>
      if ( x13 and x10 and x7 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_pp <= s2;

      elsif ( x13 and x10 and not x7 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_pp <= s9;

      elsif ( x13 and not x10 ) = '1' then
         current_pp <= s1;

      elsif ( not x13 and x12 and x15 and x9 ) = '1' then
         current_pp <= s5;

      elsif ( not x13 and x12 and x15 and not x9 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_pp <= s9;

      elsif ( not x13 and x12 and not x15 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_pp <= s3;

      else
         y11 <= '1' ;
         y18 <= '1' ;
         current_pp <= s4;

      end if;

   when s6 =>
      if ( x13 and x10 and x9 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_pp <= s5;

      elsif ( x13 and x10 and not x9 and x17 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s7;

      elsif ( x13 and x10 and not x9 and not x17 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_pp <= s3;

      elsif ( x13 and not x10 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_pp <= s2;

      elsif ( not x13 and x1 and x12 and x2 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_pp <= s2;

      elsif ( not x13 and x1 and x12 and not x2 and x3 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s7;

      elsif ( not x13 and x1 and x12 and not x2 and not x3 ) = '1' then
         current_pp <= s6;

      elsif ( not x13 and x1 and not x12 and x5 and x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_pp <= s10;

      elsif ( not x13 and x1 and not x12 and x5 and not x3 and x4 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s11;

      elsif ( not x13 and x1 and not x12 and x5 and not x3 and not x4 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_pp <= s9;

      elsif ( not x13 and x1 and not x12 and not x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_pp <= s3;

      elsif ( not x13 and not x1 and x12 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_pp <= s5;

      elsif ( not x13 and not x1 and not x12 and x2 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_pp <= s2;

      else
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s7;

      end if;

   when s7 =>
      if ( x13 and x10 and x17 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s11;

      elsif ( x13 and x10 and not x17 and x15 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s7;

      elsif ( x13 and x10 and not x17 and not x15 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_pp <= s3;

      elsif ( x13 and not x10 and x3 and x15 ) = '1' then
         current_pp <= s7;

      elsif ( x13 and not x10 and x3 and not x15 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_pp <= s3;

      elsif ( x13 and not x10 and not x3 and x4 and x5 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_pp <= s4;

      elsif ( x13 and not x10 and not x3 and x4 and not x5 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_pp <= s5;

      elsif ( x13 and not x10 and not x3 and not x4 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_pp <= s2;

      elsif ( not x13 and x12 and x4 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_pp <= s4;

      elsif ( not x13 and x12 and not x4 ) = '1' then
         current_pp <= s1;

      elsif ( not x13 and not x12 and x10 and x11 ) = '1' then
         current_pp <= s1;

      elsif ( not x13 and not x12 and x10 and not x11 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         current_pp <= s13;

      else
         y11 <= '1' ;
         y18 <= '1' ;
         current_pp <= s4;

      end if;

   when s8 =>
      if ( x13 ) = '1' then
         y4 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_pp <= s6;

      elsif ( not x13 and x10 and x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y9 <= '1' ;
         current_pp <= s14;

      elsif ( not x13 and x10 and not x5 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         y26 <= '1' ;
         current_pp <= s15;

      else
         y11 <= '1' ;
         y23 <= '1' ;
         current_pp <= s9;

      end if;

   when s9 =>
      if ( x13 and x20 ) = '1' then
         current_pp <= s1;

      elsif ( x13 and not x20 ) = '1' then
         y11 <= '1' ;
         y18 <= '1' ;
         current_pp <= s4;

      elsif ( not x13 and x12 ) = '1' then
         current_pp <= s1;

      elsif ( not x13 and not x12 and x10 and x3 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_pp <= s2;

      elsif ( not x13 and not x12 and x10 and not x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_pp <= s10;

      elsif ( not x13 and not x12 and not x10 and x19 and x16 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_pp <= s16;

      elsif ( not x13 and not x12 and not x10 and x19 and not x16 ) = '1' then
         current_pp <= s1;

      else
         y2 <= '1' ;
         y20 <= '1' ;
         y25 <= '1' ;
         current_pp <= s8;

      end if;

   when s10 =>
      if ( x10 and x7 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s11;

      elsif ( x10 and not x7 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_pp <= s16;

      else
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_pp <= s3;

      end if;

   when s11 =>
      if ( x13 and x8 and x1 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_pp <= s2;

      elsif ( x13 and x8 and not x1 and x14 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_pp <= s5;

      elsif ( x13 and x8 and not x1 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_pp <= s3;

      elsif ( x13 and not x8 ) = '1' then
         y2 <= '1' ;
         y20 <= '1' ;
         y25 <= '1' ;
         current_pp <= s8;

      elsif ( not x13 and x10 ) = '1' then
         current_pp <= s1;

      elsif ( not x13 and not x10 and x6 and x7 and x5 and x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_pp <= s10;

      elsif ( not x13 and not x10 and x6 and x7 and x5 and not x3 and x4 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s11;

      elsif ( not x13 and not x10 and x6 and x7 and x5 and not x3 and not x4 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_pp <= s9;

      elsif ( not x13 and not x10 and x6 and x7 and not x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_pp <= s3;

      elsif ( not x13 and not x10 and x6 and not x7 and x8 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_pp <= s16;

      elsif ( not x13 and not x10 and x6 and not x7 and not x8 and x5 and x3 ) = '1' then
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_pp <= s10;

      elsif ( not x13 and not x10 and x6 and not x7 and not x8 and x5 and not x3 and x4 ) = '1' then
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s11;

      elsif ( not x13 and not x10 and x6 and not x7 and not x8 and x5 and not x3 and not x4 ) = '1' then
         y11 <= '1' ;
         y23 <= '1' ;
         current_pp <= s9;

      elsif ( not x13 and not x10 and x6 and not x7 and not x8 and not x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_pp <= s3;

      elsif ( not x13 and not x10 and not x6 and x16 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_pp <= s16;

      else
         current_pp <= s1;

      end if;

   when s12 =>
      if ( x6 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y20 <= '1' ;
         current_pp <= s17;

      else
         y19 <= '1' ;
         y20 <= '1' ;
         y22 <= '1' ;
         y26 <= '1' ;
         current_pp <= s15;

      end if;

   when s13 =>
      if ( x9 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s7;

      else
         y15 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s11;

      end if;

   when s14 =>
         y7 <= '1' ;
         y13 <= '1' ;
         y28 <= '1' ;
         current_pp <= s5;

   when s15 =>
      if ( x8 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_pp <= s3;

      else
         y6 <= '1' ;
         y7 <= '1' ;
         y20 <= '1' ;
         current_pp <= s17;

      end if;

   when s16 =>
      if ( x10 and x15 ) = '1' then
         current_pp <= s1;

      elsif ( x10 and not x15 ) = '1' then
         y16 <= '1' ;
         y22 <= '1' ;
         y24 <= '1' ;
         current_pp <= s7;

      else
         current_pp <= s1;

      end if;

   when s17 =>
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y5 <= '1' ;
         current_pp <= s3;

   end case;
   end proc_pp;

   begin
      if ( rst = '1' ) then
	y1   <= '0' ;	y2   <= '0' ;	y3   <= '0' ;	y4   <= '0' ;
	y5   <= '0' ;	y6   <= '0' ;	y7   <= '0' ;	y8   <= '0' ;
	y9   <= '0' ;	y10  <= '0' ;	y11  <= '0' ;	y12  <= '0' ;
	y13  <= '0' ;	y14  <= '0' ;	y15  <= '0' ;	y16  <= '0' ;
	y17  <= '0' ;	y18  <= '0' ;	y19  <= '0' ;	y20  <= '0' ;
	y21  <= '0' ;	y22  <= '0' ;	y23  <= '0' ;	y24  <= '0' ;
	y25  <= '0' ;	y26  <= '0' ;	y27  <= '0' ;	y28  <= '0' ;

	current_pp <= s1;
      elsif (clk'event and clk ='1') then
        proc_pp;
      end if;
   end process;
end ARC;
