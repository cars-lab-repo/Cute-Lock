library ieee;
use ieee.std_logic_1164.all;

entity proc888 is
   port ( clk,rst,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,
	x16,x17,x18,x19,x20 : in std_logic;
        y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,
	y16,y17,y18,y19,y20,y21,y22,y23,y24,y25,y26,y27,y28,y29,y30,
	y31,y32,y33,y34,y35,y36,y37,y38,y39,y40,y41,y42,y43,y44,y45
	 : out std_logic );
end proc888;

architecture ARC of proc888 is

   type states_proc888 is ( s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,
	s16,s17,s18,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29,s30,
	s31,s32,s33,s34,s35,s36,s37,s38,s39,s40,s41,s42,s43,s44,s45,
	s46,s47,s48,s49,s50,s51,s52,s53,s54,s55,s56,s57,s58,s59,s60,
	s61,s62,s63,s64,s65,s66,s67,s68,s69,s70,s71,s72,s73,s74 );
   signal current_proc888 : states_proc888;

begin
   process (clk , rst)
   procedure proc_proc888 is
   begin

	y1   <= '0' ;	y2   <= '0' ;	y3   <= '0' ;	y4   <= '0' ;
	y5   <= '0' ;	y6   <= '0' ;	y7   <= '0' ;	y8   <= '0' ;
	y9   <= '0' ;	y10  <= '0' ;	y11  <= '0' ;	y12  <= '0' ;
	y13  <= '0' ;	y14  <= '0' ;	y15  <= '0' ;	y16  <= '0' ;
	y17  <= '0' ;	y18  <= '0' ;	y19  <= '0' ;	y20  <= '0' ;
	y21  <= '0' ;	y22  <= '0' ;	y23  <= '0' ;	y24  <= '0' ;
	y25  <= '0' ;	y26  <= '0' ;	y27  <= '0' ;	y28  <= '0' ;
	y29  <= '0' ;	y30  <= '0' ;	y31  <= '0' ;	y32  <= '0' ;
	y33  <= '0' ;	y34  <= '0' ;	y35  <= '0' ;	y36  <= '0' ;
	y37  <= '0' ;	y38  <= '0' ;	y39  <= '0' ;	y40  <= '0' ;
	y41  <= '0' ;	y42  <= '0' ;	y43  <= '0' ;	y44  <= '0' ;
	y45  <= '0' ;

   case current_proc888 is
   when s1 =>
      if ( x6 and x5 and x20 and x19 ) = '1' then
         y40 <= '1' ;
         y18 <= '1' ;
         y9 <= '1' ;
         y8 <= '1' ;
         y25 <= '1' ;
         current_proc888 <= s2;

      elsif ( x6 and x5 and x20 and not x19 ) = '1' then
         y40 <= '1' ;
         y8 <= '1' ;
         y43 <= '1' ;
         current_proc888 <= s3;

      elsif ( x6 and x5 and not x20 and x19 ) = '1' then
         y40 <= '1' ;
         y8 <= '1' ;
         y18 <= '1' ;
         y9 <= '1' ;
         y45 <= '1' ;
         current_proc888 <= s4;

      elsif ( x6 and x5 and not x20 and not x19 ) = '1' then
         y40 <= '1' ;
         y9 <= '1' ;
         y2 <= '1' ;
         y43 <= '1' ;
         current_proc888 <= s5;

      elsif ( x6 and not x5 and x4 ) = '1' then
         y6 <= '1' ;
         y40 <= '1' ;
         y18 <= '1' ;
         y1 <= '1' ;
         y8 <= '1' ;
         current_proc888 <= s6;

      elsif ( x6 and not x5 and not x4 ) = '1' then
         y11 <= '1' ;
         y40 <= '1' ;
         y2 <= '1' ;
         y20 <= '1' ;
         current_proc888 <= s7;

      else
         current_proc888 <= s1;

      end if;

   when s2 =>
         y17 <= '1' ;
         current_proc888 <= s8;

   when s3 =>
         y17 <= '1' ;
         current_proc888 <= s9;

   when s4 =>
         y17 <= '1' ;
         current_proc888 <= s10;

   when s5 =>
         y17 <= '1' ;
         current_proc888 <= s11;

   when s6 =>
         y17 <= '1' ;
         current_proc888 <= s12;

   when s7 =>
         y28 <= '1' ;
         current_proc888 <= s13;

   when s8 =>
         y18 <= '1' ;
         y9 <= '1' ;
         y1 <= '1' ;
         y25 <= '1' ;
         current_proc888 <= s1;

   when s9 =>
         y44 <= '1' ;
         current_proc888 <= s1;

   when s10 =>
         y18 <= '1' ;
         y9 <= '1' ;
         y1 <= '1' ;
         y45 <= '1' ;
         current_proc888 <= s1;

   when s11 =>
         y2 <= '1' ;
         y44 <= '1' ;
         current_proc888 <= s1;

   when s12 =>
         y18 <= '1' ;
         y1 <= '1' ;
         y2 <= '1' ;
         y45 <= '1' ;
         current_proc888 <= s14;

   when s13 =>
         y11 <= '1' ;
         y40 <= '1' ;
         y34 <= '1' ;
         y35 <= '1' ;
         current_proc888 <= s15;

   when s14 =>
         y17 <= '1' ;
         current_proc888 <= s16;

   when s15 =>
         y28 <= '1' ;
         current_proc888 <= s17;

   when s16 =>
         y18 <= '1' ;
         y1 <= '1' ;
         y25 <= '1' ;
         current_proc888 <= s18;

   when s17 =>
      if ( x12 and x14 and x13 and x16 ) = '1' then
         y33 <= '1' ;
         current_proc888 <= s19;

      elsif ( x12 and x14 and x13 and not x16 ) = '1' then
         y32 <= '1' ;
         current_proc888 <= s19;

      elsif ( x12 and x14 and not x13 ) = '1' then
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s20;

      elsif ( x12 and not x14 and x15 and x13 and x16 ) = '1' then
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s20;

      elsif ( x12 and not x14 and x15 and x13 and not x16 ) = '1' then
         y18 <= '1' ;
         y9 <= '1' ;
         y2 <= '1' ;
         y16 <= '1' ;
         y10 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y29 <= '1' ;
         current_proc888 <= s21;

      elsif ( x12 and not x14 and x15 and not x13 ) = '1' then
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s20;

      elsif ( x12 and not x14 and not x15 and x13 and x16 and x11 ) = '1' then
         y28 <= '1' ;
         current_proc888 <= s22;

      elsif ( x12 and not x14 and not x15 and x13 and x16 and not x11 and x18 and x10 ) = '1' then
         y42 <= '1' ;
         current_proc888 <= s1;

      elsif ( x12 and not x14 and not x15 and x13 and x16 and not x11 and x18 and not x10 ) = '1' then
         current_proc888 <= s1;

      elsif ( x12 and not x14 and not x15 and x13 and x16 and not x11 and not x18 ) = '1' then
         current_proc888 <= s1;

      elsif ( x12 and not x14 and not x15 and x13 and not x16 and x10 ) = '1' then
         y28 <= '1' ;
         current_proc888 <= s22;

      elsif ( x12 and not x14 and not x15 and x13 and not x16 and not x10 and x18 and x11 ) = '1' then
         y42 <= '1' ;
         current_proc888 <= s1;

      elsif ( x12 and not x14 and not x15 and x13 and not x16 and not x10 and x18 and not x11 ) = '1' then
         current_proc888 <= s1;

      elsif ( x12 and not x14 and not x15 and x13 and not x16 and not x10 and not x18 ) = '1' then
         current_proc888 <= s1;

      elsif ( x12 and not x14 and not x15 and not x13 and x3 ) = '1' then
         y11 <= '1' ;
         y40 <= '1' ;
         y2 <= '1' ;
         y36 <= '1' ;
         current_proc888 <= s23;

      elsif ( x12 and not x14 and not x15 and not x13 and not x3 and x16 and x2 ) = '1' then
         y41 <= '1' ;
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s24;

      elsif ( x12 and not x14 and not x15 and not x13 and not x3 and x16 and not x2 ) = '1' then
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s20;

      elsif ( x12 and not x14 and not x15 and not x13 and not x3 and not x16 ) = '1' then
         y41 <= '1' ;
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s24;

      elsif ( not x12 and x3 ) = '1' then
         y11 <= '1' ;
         y40 <= '1' ;
         y2 <= '1' ;
         y36 <= '1' ;
         current_proc888 <= s23;

      elsif ( not x12 and not x3 and x13 and x15 and x16 ) = '1' then
         y41 <= '1' ;
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s24;

      elsif ( not x12 and not x3 and x13 and x15 and not x16 and x9 ) = '1' then
         y41 <= '1' ;
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s24;

      elsif ( not x12 and not x3 and x13 and x15 and not x16 and not x9 and x18 and x10 ) = '1' then
         y42 <= '1' ;
         current_proc888 <= s1;

      elsif ( not x12 and not x3 and x13 and x15 and not x16 and not x9 and x18 and not x10 and x11 ) = '1' then
         y42 <= '1' ;
         current_proc888 <= s1;

      elsif ( not x12 and not x3 and x13 and x15 and not x16 and not x9 and x18 and not x10 and not x11 ) = '1' then
         current_proc888 <= s1;

      elsif ( not x12 and not x3 and x13 and x15 and not x16 and not x9 and not x18 ) = '1' then
         current_proc888 <= s1;

      elsif ( not x12 and not x3 and x13 and not x15 and x16 and x8 ) = '1' then
         y41 <= '1' ;
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s24;

      elsif ( not x12 and not x3 and x13 and not x15 and x16 and not x8 and x18 and x10 ) = '1' then
         y42 <= '1' ;
         current_proc888 <= s1;

      elsif ( not x12 and not x3 and x13 and not x15 and x16 and not x8 and x18 and not x10 and x11 ) = '1' then
         y42 <= '1' ;
         current_proc888 <= s1;

      elsif ( not x12 and not x3 and x13 and not x15 and x16 and not x8 and x18 and not x10 and not x11 ) = '1' then
         current_proc888 <= s1;

      elsif ( not x12 and not x3 and x13 and not x15 and x16 and not x8 and not x18 ) = '1' then
         current_proc888 <= s1;

      elsif ( not x12 and not x3 and x13 and not x15 and not x16 and x7 ) = '1' then
         y41 <= '1' ;
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s24;

      elsif ( not x12 and not x3 and x13 and not x15 and not x16 and not x7 and x18 and x10 ) = '1' then
         y42 <= '1' ;
         current_proc888 <= s1;

      elsif ( not x12 and not x3 and x13 and not x15 and not x16 and not x7 and x18 and not x10 and x11 ) = '1' then
         y42 <= '1' ;
         current_proc888 <= s1;

      elsif ( not x12 and not x3 and x13 and not x15 and not x16 and not x7 and x18 and not x10 and not x11 ) = '1' then
         current_proc888 <= s1;

      elsif ( not x12 and not x3 and x13 and not x15 and not x16 and not x7 and not x18 ) = '1' then
         current_proc888 <= s1;

      else
         y41 <= '1' ;
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s24;

      end if;

   when s18 =>
         y17 <= '1' ;
         current_proc888 <= s25;

   when s19 =>
      if ( x18 and x10 ) = '1' then
         y42 <= '1' ;
         current_proc888 <= s1;

      elsif ( x18 and not x10 and x11 ) = '1' then
         y42 <= '1' ;
         current_proc888 <= s1;

      elsif ( x18 and not x10 and not x11 ) = '1' then
         current_proc888 <= s1;

      else
         current_proc888 <= s1;

      end if;

   when s20 =>
         y23 <= '1' ;
         current_proc888 <= s26;

   when s21 =>
         y21 <= '1' ;
         y22 <= '1' ;
         y9 <= '1' ;
         current_proc888 <= s27;

   when s22 =>
         y28 <= '1' ;
         current_proc888 <= s28;

   when s23 =>
         y28 <= '1' ;
         current_proc888 <= s29;

   when s24 =>
         y23 <= '1' ;
         current_proc888 <= s30;

   when s25 =>
         y18 <= '1' ;
         y1 <= '1' ;
         y2 <= '1' ;
         y25 <= '1' ;
         current_proc888 <= s31;

   when s26 =>
         y24 <= '1' ;
         y10 <= '1' ;
         y34 <= '1' ;
         y8 <= '1' ;
         current_proc888 <= s32;

   when s27 =>
         y23 <= '1' ;
         current_proc888 <= s33;

   when s28 =>
         y28 <= '1' ;
         current_proc888 <= s34;

   when s29 =>
         y11 <= '1' ;
         y40 <= '1' ;
         y34 <= '1' ;
         y37 <= '1' ;
         current_proc888 <= s35;

   when s30 =>
         y24 <= '1' ;
         y10 <= '1' ;
         y34 <= '1' ;
         y8 <= '1' ;
         current_proc888 <= s36;

   when s31 =>
         y18 <= '1' ;
         y9 <= '1' ;
         y1 <= '1' ;
         y2 <= '1' ;
         y16 <= '1' ;
         y34 <= '1' ;
         y33 <= '1' ;
         y19 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_proc888 <= s1;

   when s32 =>
      if ( x13 ) = '1' then
         y30 <= '1' ;
         y31 <= '1' ;
         current_proc888 <= s19;

      elsif ( not x13 and x15 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_proc888 <= s37;

      elsif ( not x13 and not x15 and x14 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_proc888 <= s37;

      else
         y41 <= '1' ;
         y9 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_proc888 <= s38;

      end if;

   when s33 =>
         y24 <= '1' ;
         y18 <= '1' ;
         y22 <= '1' ;
         current_proc888 <= s19;

   when s34 =>
         y28 <= '1' ;
         current_proc888 <= s19;

   when s35 =>
         y28 <= '1' ;
         current_proc888 <= s39;

   when s36 =>
      if ( x12 and x16 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_proc888 <= s40;

      elsif ( x12 and not x16 and x2 ) = '1' then
         y6 <= '1' ;
         y9 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_proc888 <= s41;

      elsif ( x12 and not x16 and not x2 ) = '1' then
         y21 <= '1' ;
         y22 <= '1' ;
         y9 <= '1' ;
         current_proc888 <= s27;

      elsif ( not x12 and x13 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_proc888 <= s19;

      elsif ( not x12 and not x13 and x2 and x14 ) = '1' then
         y6 <= '1' ;
         y8 <= '1' ;
         y4 <= '1' ;
         current_proc888 <= s42;

      elsif ( not x12 and not x13 and x2 and not x14 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_proc888 <= s40;

      elsif ( not x12 and not x13 and not x2 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_proc888 <= s43;

      else
         y1 <= '1' ;
         y10 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_proc888 <= s44;

      end if;

   when s37 =>
         y9 <= '1' ;
         y2 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_proc888 <= s45;

   when s38 =>
         y23 <= '1' ;
         current_proc888 <= s46;

   when s39 =>
      if ( x12 and x1 and x16 and x2 ) = '1' then
         y11 <= '1' ;
         y8 <= '1' ;
         y4 <= '1' ;
         current_proc888 <= s48;

      elsif ( x12 and x1 and x16 and not x2 and x17 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y8 <= '1' ;
         y21 <= '1' ;
         y25 <= '1' ;
         current_proc888 <= s41;

      elsif ( x12 and x1 and x16 and not x2 and not x17 ) = '1' then
         y41 <= '1' ;
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s52;

      elsif ( x12 and x1 and not x16 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_proc888 <= s47;

      elsif ( x12 and not x1 and x2 ) = '1' then
         y11 <= '1' ;
         y8 <= '1' ;
         y4 <= '1' ;
         current_proc888 <= s48;

      elsif ( x12 and not x1 and not x2 and x17 and x16 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y8 <= '1' ;
         y21 <= '1' ;
         y25 <= '1' ;
         current_proc888 <= s41;

      elsif ( x12 and not x1 and not x2 and x17 and not x16 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_proc888 <= s49;

      elsif ( x12 and not x1 and not x2 and not x17 ) = '1' then
         y41 <= '1' ;
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s52;

      elsif ( not x12 and x13 and x15 and x16 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_proc888 <= s19;

      elsif ( not x12 and x13 and x15 and x16 and not x1 and x2 ) = '1' then
         y11 <= '1' ;
         y8 <= '1' ;
         y4 <= '1' ;
         current_proc888 <= s48;

      elsif ( not x12 and x13 and x15 and x16 and not x1 and not x2 and x17 ) = '1' then
         y11 <= '1' ;
         y8 <= '1' ;
         y26 <= '1' ;
         current_proc888 <= s50;

      elsif ( not x12 and x13 and x15 and x16 and not x1 and not x2 and not x17 ) = '1' then
         y41 <= '1' ;
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s52;

      elsif ( not x12 and x13 and x15 and not x16 and x9 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_proc888 <= s19;

      elsif ( not x12 and x13 and x15 and not x16 and x9 and not x1 and x2 ) = '1' then
         y11 <= '1' ;
         y8 <= '1' ;
         y4 <= '1' ;
         current_proc888 <= s48;

      elsif ( not x12 and x13 and x15 and not x16 and x9 and not x1 and not x2 and x17 ) = '1' then
         y11 <= '1' ;
         y8 <= '1' ;
         y26 <= '1' ;
         current_proc888 <= s50;

      elsif ( not x12 and x13 and x15 and not x16 and x9 and not x1 and not x2 and not x17 ) = '1' then
         y41 <= '1' ;
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s52;

      elsif ( not x12 and x13 and x15 and not x16 and not x9 and x18 and x10 ) = '1' then
         y42 <= '1' ;
         current_proc888 <= s1;

      elsif ( not x12 and x13 and x15 and not x16 and not x9 and x18 and not x10 and x11 ) = '1' then
         y42 <= '1' ;
         current_proc888 <= s1;

      elsif ( not x12 and x13 and x15 and not x16 and not x9 and x18 and not x10 and not x11 ) = '1' then
         current_proc888 <= s1;

      elsif ( not x12 and x13 and x15 and not x16 and not x9 and not x18 ) = '1' then
         current_proc888 <= s1;

      elsif ( not x12 and x13 and not x15 and x16 and x8 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_proc888 <= s19;

      elsif ( not x12 and x13 and not x15 and x16 and x8 and not x1 and x2 ) = '1' then
         y11 <= '1' ;
         y8 <= '1' ;
         y4 <= '1' ;
         current_proc888 <= s48;

      elsif ( not x12 and x13 and not x15 and x16 and x8 and not x1 and not x2 and x17 ) = '1' then
         y11 <= '1' ;
         y8 <= '1' ;
         y26 <= '1' ;
         current_proc888 <= s50;

      elsif ( not x12 and x13 and not x15 and x16 and x8 and not x1 and not x2 and not x17 ) = '1' then
         y41 <= '1' ;
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s52;

      elsif ( not x12 and x13 and not x15 and x16 and not x8 and x18 and x10 ) = '1' then
         y42 <= '1' ;
         current_proc888 <= s1;

      elsif ( not x12 and x13 and not x15 and x16 and not x8 and x18 and not x10 and x11 ) = '1' then
         y42 <= '1' ;
         current_proc888 <= s1;

      elsif ( not x12 and x13 and not x15 and x16 and not x8 and x18 and not x10 and not x11 ) = '1' then
         current_proc888 <= s1;

      elsif ( not x12 and x13 and not x15 and x16 and not x8 and not x18 ) = '1' then
         current_proc888 <= s1;

      elsif ( not x12 and x13 and not x15 and not x16 and x7 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_proc888 <= s19;

      elsif ( not x12 and x13 and not x15 and not x16 and x7 and not x1 and x2 ) = '1' then
         y11 <= '1' ;
         y8 <= '1' ;
         y4 <= '1' ;
         current_proc888 <= s48;

      elsif ( not x12 and x13 and not x15 and not x16 and x7 and not x1 and not x2 and x17 ) = '1' then
         y11 <= '1' ;
         y8 <= '1' ;
         y26 <= '1' ;
         current_proc888 <= s50;

      elsif ( not x12 and x13 and not x15 and not x16 and x7 and not x1 and not x2 and not x17 ) = '1' then
         y41 <= '1' ;
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s52;

      elsif ( not x12 and x13 and not x15 and not x16 and not x7 and x18 and x10 ) = '1' then
         y42 <= '1' ;
         current_proc888 <= s1;

      elsif ( not x12 and x13 and not x15 and not x16 and not x7 and x18 and not x10 and x11 ) = '1' then
         y42 <= '1' ;
         current_proc888 <= s1;

      elsif ( not x12 and x13 and not x15 and not x16 and not x7 and x18 and not x10 and not x11 ) = '1' then
         current_proc888 <= s1;

      elsif ( not x12 and x13 and not x15 and not x16 and not x7 and not x18 ) = '1' then
         current_proc888 <= s1;

      elsif ( not x12 and not x13 and x1 and x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_proc888 <= s47;

      elsif ( not x12 and not x13 and x1 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_proc888 <= s44;

      elsif ( not x12 and not x13 and not x1 and x2 ) = '1' then
         y11 <= '1' ;
         y8 <= '1' ;
         y4 <= '1' ;
         current_proc888 <= s48;

      elsif ( not x12 and not x13 and not x1 and not x2 and x17 and x14 ) = '1' then
         y11 <= '1' ;
         y9 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s50;

      elsif ( not x12 and not x13 and not x1 and not x2 and x17 and not x14 ) = '1' then
         y11 <= '1' ;
         y8 <= '1' ;
         y4 <= '1' ;
         current_proc888 <= s51;

      else
         y41 <= '1' ;
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s52;

      end if;

   when s40 =>
      if ( x12 ) = '1' then
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s53;

      else
         y4 <= '1' ;
         current_proc888 <= s42;

      end if;

   when s41 =>
         y17 <= '1' ;
         y23 <= '1' ;
         current_proc888 <= s54;

   when s42 =>
         y17 <= '1' ;
         current_proc888 <= s55;

   when s43 =>
         y9 <= '1' ;
         y2 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y16 <= '1' ;
         current_proc888 <= s56;

   when s44 =>
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s53;

   when s45 =>
         y23 <= '1' ;
         current_proc888 <= s57;

   when s46 =>
         y24 <= '1' ;
         y18 <= '1' ;
         y22 <= '1' ;
         current_proc888 <= s19;

   when s47 =>
      if ( x12 ) = '1' then
         y21 <= '1' ;
         y22 <= '1' ;
         y9 <= '1' ;
         current_proc888 <= s58;

      else
         y6 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_proc888 <= s43;

      end if;

   when s48 =>
         y17 <= '1' ;
         current_proc888 <= s59;

   when s49 =>
         y6 <= '1' ;
         y9 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_proc888 <= s41;

   when s50 =>
         y17 <= '1' ;
         current_proc888 <= s60;

   when s51 =>
         y17 <= '1' ;
         current_proc888 <= s61;

   when s52 =>
         y23 <= '1' ;
         current_proc888 <= s62;

   when s53 =>
         y23 <= '1' ;
         current_proc888 <= s63;

   when s54 =>
      if ( x16 ) = '1' then
         y24 <= '1' ;
         y1 <= '1' ;
         y25 <= '1' ;
         current_proc888 <= s19;

      else
         y24 <= '1' ;
         y22 <= '1' ;
         current_proc888 <= s19;

      end if;

   when s55 =>
         y5 <= '1' ;
         current_proc888 <= s64;

   when s56 =>
         y21 <= '1' ;
         y22 <= '1' ;
         y9 <= '1' ;
         current_proc888 <= s58;

   when s57 =>
         y24 <= '1' ;
         y16 <= '1' ;
         y22 <= '1' ;
         current_proc888 <= s19;

   when s58 =>
         y23 <= '1' ;
         current_proc888 <= s65;

   when s59 =>
         y5 <= '1' ;
         current_proc888 <= s66;

   when s60 =>
      if ( x13 ) = '1' then
         y27 <= '1' ;
         current_proc888 <= s19;

      else
         y8 <= '1' ;
         current_proc888 <= s67;

      end if;

   when s61 =>
         y5 <= '1' ;
         current_proc888 <= s44;

   when s62 =>
         y24 <= '1' ;
         y10 <= '1' ;
         y34 <= '1' ;
         y8 <= '1' ;
         current_proc888 <= s68;

   when s63 =>
         y24 <= '1' ;
         y10 <= '1' ;
         y34 <= '1' ;
         y8 <= '1' ;
         current_proc888 <= s69;

   when s64 =>
      if ( x14 ) = '1' then
         y18 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y10 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_proc888 <= s67;

      else
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s53;

      end if;

   when s65 =>
         y24 <= '1' ;
         y18 <= '1' ;
         y22 <= '1' ;
         current_proc888 <= s19;

   when s66 =>
         y18 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y10 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_proc888 <= s70;

   when s67 =>
         y6 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_proc888 <= s43;

   when s68 =>
         y38 <= '1' ;
         y39 <= '1' ;
         current_proc888 <= s71;

   when s69 =>
      if ( x12 ) = '1' then
         y9 <= '1' ;
         y25 <= '1' ;
         current_proc888 <= s72;

      else
         y6 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_proc888 <= s43;

      end if;

   when s70 =>
      if ( x17 and x12 and x16 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y8 <= '1' ;
         y21 <= '1' ;
         y25 <= '1' ;
         current_proc888 <= s41;

      elsif ( x17 and x12 and not x16 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_proc888 <= s49;

      elsif ( x17 and not x12 and x13 ) = '1' then
         y11 <= '1' ;
         y8 <= '1' ;
         y26 <= '1' ;
         current_proc888 <= s50;

      elsif ( x17 and not x12 and not x13 and x14 ) = '1' then
         y11 <= '1' ;
         y9 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s50;

      elsif ( x17 and not x12 and not x13 and not x14 ) = '1' then
         y11 <= '1' ;
         y8 <= '1' ;
         y4 <= '1' ;
         current_proc888 <= s51;

      else
         y41 <= '1' ;
         y1 <= '1' ;
         y21 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s52;

      end if;

   when s71 =>
         y9 <= '1' ;
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y10 <= '1' ;
         y34 <= '1' ;
         y36 <= '1' ;
         y37 <= '1' ;
         current_proc888 <= s73;

   when s72 =>
         y17 <= '1' ;
         current_proc888 <= s74;

   when s73 =>
      if ( x12 and x16 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y8 <= '1' ;
         y21 <= '1' ;
         y25 <= '1' ;
         current_proc888 <= s41;

      elsif ( x12 and not x16 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_proc888 <= s49;

      elsif ( not x12 and x13 ) = '1' then
         y11 <= '1' ;
         y8 <= '1' ;
         y26 <= '1' ;
         current_proc888 <= s50;

      elsif ( not x12 and not x13 and x14 ) = '1' then
         y11 <= '1' ;
         y9 <= '1' ;
         y7 <= '1' ;
         current_proc888 <= s50;

      else
         y11 <= '1' ;
         y8 <= '1' ;
         y4 <= '1' ;
         current_proc888 <= s51;

      end if;

   when s74 =>
         y25 <= '1' ;
         y18 <= '1' ;
         current_proc888 <= s19;

   end case;
   end proc_proc888;

   begin
      if ( rst = '1' ) then
	y1   <= '0' ;	y2   <= '0' ;	y3   <= '0' ;	y4   <= '0' ;
	y5   <= '0' ;	y6   <= '0' ;	y7   <= '0' ;	y8   <= '0' ;
	y9   <= '0' ;	y10  <= '0' ;	y11  <= '0' ;	y12  <= '0' ;
	y13  <= '0' ;	y14  <= '0' ;	y15  <= '0' ;	y16  <= '0' ;
	y17  <= '0' ;	y18  <= '0' ;	y19  <= '0' ;	y20  <= '0' ;
	y21  <= '0' ;	y22  <= '0' ;	y23  <= '0' ;	y24  <= '0' ;
	y25  <= '0' ;	y26  <= '0' ;	y27  <= '0' ;	y28  <= '0' ;
	y29  <= '0' ;	y30  <= '0' ;	y31  <= '0' ;	y32  <= '0' ;
	y33  <= '0' ;	y34  <= '0' ;	y35  <= '0' ;	y36  <= '0' ;
	y37  <= '0' ;	y38  <= '0' ;	y39  <= '0' ;	y40  <= '0' ;
	y41  <= '0' ;	y42  <= '0' ;	y43  <= '0' ;	y44  <= '0' ;
	y45  <= '0' ;
	current_proc888 <= s1;
      elsif (clk'event and clk ='1') then
        proc_proc888;
      end if;
   end process;
end ARC;
