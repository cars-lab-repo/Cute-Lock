module rexm ( clk,rst,
	x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15,
	x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30,
	x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45,
	x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60,
	x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, 
	y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15,
	y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30,
	y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45,
	y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60,
	y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y77, y78, y79, y80, y81, y84, y86, y88, y90,
	y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y102, y110, y112);

input clk, rst, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15,
	x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30,
	x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45,
	x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60,
	x61, x62, x63, x64, x65, x66, x67, x68, x69, x70;
output y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15,
	y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30,
	y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45,
	y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60,
	y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y77, y78, y79, y80, y81, y84, y86, y88, y90,
	y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y102, y110, y112;
reg y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15,
	y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30,
	y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45,
	y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60,
	y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y77, y78, y79, y80, y81, y84, y86, y88, y90,
	y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y102, y110, y112;

parameter s1=1, s2=2, s3=3, s4=4, s5=5, s6=6, s7=7, s8=8, s9=9, s10=10,
	s11=11, s12=12, s13=13, s14=14, s15=15, s16=16, s17=17, s18=18, s19=19, s20=20,
	s21=21, s22=22, s23=23, s24=24, s25=25, s26=26, s27=27, s28=28, s29=29, s30=30,
	s31=31, s32=32, s33=33, s34=34, s35=35, s36=36, s37=37, s38=38, s39=39, s40=40,
	s41=41, s42=42, s43=43, s44=44, s45=45, s46=46, s47=47, s48=48, s49=49, s50=50,
	s51=51, s52=52, s53=53, s54=54, s55=55, s56=56, s57=57, s58=58, s59=59, s60=60,
	s61=61, s62=62, s63=63, s64=64, s65=65, s66=66, s67=67, s68=68, s69=69, s70=70,
	s71=71, s72=72, s73=73, s74=74, s75=75, s76=76, s77=77, s78=78, s79=79, s80=80,
	s81=81, s82=82, s83=83, s84=84, s85=85, s86=86, s87=87, s88=88, s89=89, s90=90,
	s91=91, s92=92, s93=93, s94=94, s95=95, s96=96, s97=97, s98=98, s99=99, s100=100,
	s101=101, s102=102, s103=103, s104=104, s105=105, s106=106, s107=107, s108=108, s109=109, s110=110,
	s111=111, s112=112, s113=113, s114=114, s115=115, s116=116, s117=117, s118=118, s119=119, s120=120,
	s121=121, s122=122, s123=123, s124=124, s125=125, s126=126, s127=127, s128=128, s129=129, s130=130,
	s131=131, s132=132, s133=133, s134=134, s135=135, s136=136, s137=137, s138=138, s139=139, s140=140,
	s141=141, s142=142, s143=143, s144=144, s145=145, s146=146, s147=147, s148=148, s149=149, s150=150,
	s151=151, s152=152, s153=153, s154=154, s155=155, s156=156, s157=157, s158=158, s159=159, s160=160,
	s161=161, s162=162, s163=163, s164=164, s165=165, s166=166, s167=167, s168=168, s169=169, s170=170,
	s171=171, s172=172, s173=173, s174=174, s175=175, s176=176, s177=177, s178=178, s179=179, s180=180,
	s181=181, s182=182, s183=183, s184=184, s185=185, s186=186, s187=187, s188=188, s189=189, s190=190,
	s191=191, s192=192, s193=193, s194=194, s195=195, s196=196, s197=197, s198=198, s199=199, s200=200,
	s201=201, s202=202, s203=203, s204=204, s205=205, s206=206, s207=207, s208=208, s209=209, s210=210,
	s211=211, s212=212, s213=213, s214=214, s215=215, s216=216, s217=217, s218=218, s219=219, s220=220,
	s221=221, s222=222, s223=223, s224=224, s225=225, s226=226, s227=227, s228=228, s229=229, s230=230,
	s231=231, s232=232, s233=233, s234=234, s235=235, s236=236, s237=237, s238=238, s239=239, s240=240,
	s241=241, s242=242, s243=243, s244=244, s245=245, s246=246, s247=247, s248=248, s249=249, s250=250,
	s251=251, s252=252, s253=253, s254=254, s255=255, s256=256, s257=257, s258=258, s259=259, s260=260,
	s261=261, s262=262, s263=263, s264=264, s265=265, s266=266, s267=267, s268=268, s269=269, s270=270,
	s271=271, s272=272, s273=273, s274=274, s275=275, s276=276, s277=277, s278=278, s279=279, s280=280,
	s281=281, s282=282, s283=283, s284=284, s285=285, s286=286, s287=287, s288=288, s289=289, s290=290,
	s291=291, s292=292, s293=293, s294=294, s295=295, s296=296, s297=297, s298=298, s299=299, s300=300,
	s301=301, s302=302, s303=303, s304=304, s305=305, s306=306, s307=307, s308=308, s309=309, s310=310,
	s311=311, s312=312, s313=313, s314=314, s315=315, s316=316, s317=317, s318=318, s319=319, s320=320,
	s321=321, s322=322, s323=323, s324=324, s325=325, s326=326, s327=327, s328=328, s329=329, s330=330,
	s331=331, s332=332, s333=333, s334=334, s335=335, s336=336, s337=337, s338=338, s339=339, s340=340,
	s341=341, s342=342, s343=343, s344=344, s345=345, s346=346, s347=347, s348=348, s349=349, s350=350,
	s351=351, s352=352, s353=353, s354=354, s355=355, s356=356, s357=357, s358=358, s359=359, s360=360,
	s361=361, s362=362, s363=363, s364=364, s365=365, s366=366, s367=367, s368=368, s369=369, s370=370,
	s371=371, s372=372, s373=373, s374=374, s375=375, s376=376, s377=377, s378=378, s379=379, s380=380,
	s381=381, s382=382, s383=383, s384=384, s385=385, s386=386, s387=387, s388=388, s389=389, s390=390,
	s391=391, s392=392, s393=393, s394=394, s395=395, s396=396, s397=397, s398=398, s399=399, s400=400,
	s401=401, s402=402, s403=403, s404=404, s405=405, s406=406, s407=407, s408=408, s409=409, s410=410,
	s411=411, s412=412, s413=413, s414=414, s415=415, s416=416, s417=417, s418=418, s419=419, s420=420,
	s421=421, s422=422, s423=423, s424=424, s425=425, s426=426, s427=427, s428=428, s429=429, s430=430,
	s431=431, s432=432, s433=433, s434=434, s435=435, s436=436, s437=437, s438=438, s439=439, s440=440,
	s441=441, s442=442, s443=443, s444=444, s445=445, s446=446, s447=447, s448=448, s449=449, s450=450,
	s451=451, s452=452, s453=453, s454=454, s455=455, s456=456, s457=457, s458=458, s459=459, s460=460,
	s461=461, s462=462, s463=463, s464=464, s465=465, s466=466, s467=467, s468=468, s469=469, s470=470,
	s471=471, s472=472, s473=473, s474=474, s475=475, s476=476, s477=477, s478=478, s479=479, s480=480,
	s481=481, s482=482, s483=483, s484=484, s485=485, s486=486, s487=487, s488=488, s489=489, s490=490,
	s491=491, s492=492, s493=493, s494=494, s495=495, s496=496, s497=497, s498=498, s499=499, s500=500,
	s501=501, s502=502, s503=503, s504=504, s505=505, s506=506, s507=507, s508=508, s509=509, s510=510,
	s511=511, s512=512, s513=513, s514=514, s515=515, s516=516, s517=517, s518=518, s519=519, s520=520,
	s521=521, s522=522, s523=523, s524=524, s525=525, s526=526, s527=527, s528=528, s529=529, s530=530,
	s531=531, s532=532, s533=533, s534=534, s535=535, s536=536, s537=537, s538=538, s539=539, s540=540,
	s541=541, s542=542, s543=543, s544=544, s545=545, s546=546, s547=547, s548=548, s549=549, s550=550,
	s551=551, s552=552, s553=553, s554=554, s555=555, s556=556, s557=557, s558=558, s559=559, s560=560,
	s561=561, s562=562, s563=563, s564=564, s565=565, s566=566, s567=567, s568=568, s569=569, s570=570,
	s571=571, s572=572, s573=573, s574=574, s575=575, s576=576, s577=577, s578=578, s579=579, s580=580,
	s581=581, s582=582, s583=583, s584=584, s585=585, s586=586, s587=587, s588=588, s589=589, s590=590,
	s591=591, s592=592, s593=593, s594=594, s595=595, s596=596, s597=597, s598=598, s599=599, s600=600,
	s601=601, s602=602, s603=603, s604=604, s605=605, s606=606, s607=607, s608=608, s609=609, s610=610,
	s611=611, s612=612, s613=613, s614=614, s615=615, s616=616, s617=617, s618=618, s619=619, s620=620,
	s621=621, s622=622, s623=623, s624=624, s625=625, s626=626, s627=627, s628=628, s629=629, s630=630,
	s631=631, s632=632, s633=633, s634=634, s635=635, s636=636, s637=637, s638=638, s639=639, s640=640,
	s641=641, s642=642, s643=643, s644=644, s645=645, s646=646, s647=647, s648=648, s649=649, s650=650,
	s651=651, s652=652, s653=653, s654=654, s655=655, s656=656, s657=657, s658=658, s659=659, s660=660,
	s661=661, s662=662, s663=663, s664=664, s665=665, s666=666, s667=667, s668=668, s669=669, s670=670,
	s671=671, s672=672, s673=673, s674=674, s675=675, s676=676, s677=677, s678=678, s679=679, s680=680,
	s681=681, s682=682, s683=683, s684=684, s685=685, s686=686, s687=687, s688=688, s689=689, s690=690,
	s691=691, s692=692, s693=693, s694=694, s695=695, s696=696, s697=697, s698=698, s699=699, s700=700,
	s701=701, s702=702, s703=703, s704=704, s705=705, s706=706, s707=707, s708=708, s709=709, s710=710,
	s711=711, s712=712, s713=713, s714=714, s715=715, s716=716, s717=717, s718=718, s719=719, s720=720,
	s721=721, s722=722, s723=723, s724=724, s725=725, s726=726, s727=727, s728=728, s729=729, s730=730,
	s731=731, s732=732, s733=733, s734=734, s735=735, s736=736, s737=737, s738=738, s739=739, s740=740,
	s741=741, s742=742, s743=743, s744=744, s745=745, s746=746, s747=747, s748=748, s749=749, s750=750,
	s751=751, s752=752, s753=753, s754=754, s755=755, s756=756, s757=757, s758=758, s759=759, s760=760,
	s761=761, s762=762, s763=763, s764=764, s765=765, s766=766, s767=767, s768=768, s769=769, s770=770,
	s771=771, s772=772, s773=773, s774=774, s775=775, s776=776, s777=777, s778=778, s779=779, s780=780,
	s781=781, s782=782, s783=783, s784=784, s785=785, s786=786, s787=787, s788=788, s789=789, s790=790,
	s791=791, s792=792, s793=793, s794=794, s795=795, s796=796, s797=797, s798=798, s799=799, s800=800,
	s801=801, s802=802, s803=803, s804=804, s805=805, s806=806, s807=807, s808=808, s809=809, s810=810,
	s811=811, s812=812, s813=813, s814=814, s815=815, s816=816, s817=817, s818=818, s819=819, s820=820,
	s821=821, s822=822, s823=823, s824=824, s825=825, s826=826, s827=827, s828=828, s829=829, s830=830,
	s831=831, s832=832, s833=833, s834=834, s835=835, s836=836, s837=837, s838=838, s839=839, s840=840,
	s841=841, s842=842, s843=843, s844=844, s845=845, s846=846, s847=847, s848=848, s849=849, s850=850,
	s851=851, s852=852, s853=853, s854=854, s855=855, s856=856, s857=857, s858=858, s859=859, s860=860,
	s861=861, s862=862, s863=863, s864=864, s865=865, s866=866, s867=867, s868=868, s869=869, s870=870,
	s871=871, s872=872, s873=873, s874=874, s875=875, s876=876, s877=877, s878=878, s879=879, s880=880,
	s881=881, s882=882, s883=883, s884=884, s885=885, s886=886, s887=887, s888=888, s889=889, s890=890,
	s891=891, s892=892, s893=893, s894=894, s895=895, s896=896, s897=897, s898=898, s899=899, s900=900,
	s901=901, s902=902, s903=903, s904=904, s905=905, s906=906, s907=907, s908=908, s909=909, s910=910,
	s911=911, s912=912, s913=913, s914=914, s915=915, s916=916, s917=917, s918=918, s919=919, s920=920,
	s921=921, s922=922, s923=923, s924=924, s925=925, s926=926, s927=927, s928=928, s929=929, s930=930,
	s931=931, s932=932, s933=933, s934=934, s935=935, s936=936, s937=937, s938=938, s939=939, s940=940,
	s941=941, s942=942, s943=943, s944=944, s945=945, s946=946, s947=947, s948=948, s949=949, s950=950,
	s951=951, s952=952, s953=953, s954=954, s955=955, s956=956, s957=957, s958=958, s959=959, s960=960,
	s961=961, s962=962, s963=963, s964=964, s965=965, s966=966, s967=967, s968=968, s969=969, s970=970,
	s971=971, s972=972, s973=973, s974=974, s975=975, s976=976, s977=977, s978=978, s979=979, s980=980,
	s981=981, s982=982, s983=983, s984=984, s985=985, s986=986, s987=987, s988=988, s989=989, s990=990,
	s991=991, s992=992, s993=993, s994=994, s995=995, s996=996, s997=997, s998=998, s999=999, s1000=1000,
	s1001=1001, s1002=1002, s1003=1003, s1004=1004, s1005=1005, s1006=1006, s1007=1007, s1008=1008, s1009=1009, s1010=1010,
	s1011=1011, s1012=1012, s1013=1013, s1014=1014, s1015=1015, s1016=1016, s1017=1017, s1018=1018, s1019=1019, s1020=1020,
	s1021=1021, s1022=1022, s1023=1023, s1024=1024, s1025=1025, s1026=1026, s1027=1027, s1028=1028, s1029=1029, s1030=1030,
	s1031=1031, s1032=1032, s1033=1033, s1034=1034, s1035=1035, s1036=1036, s1037=1037, s1038=1038, s1039=1039, s1040=1040,
	s1041=1041, s1042=1042, s1043=1043, s1044=1044, s1045=1045, s1046=1046, s1047=1047, s1048=1048, s1049=1049, s1050=1050,
	s1051=1051, s1052=1052, s1053=1053, s1054=1054, s1055=1055, s1056=1056, s1057=1057, s1058=1058, s1059=1059, s1060=1060,
	s1061=1061, s1062=1062, s1063=1063, s1064=1064, s1065=1065, s1066=1066, s1067=1067, s1068=1068, s1069=1069, s1070=1070,
	s1071=1071, s1072=1072, s1073=1073, s1074=1074, s1075=1075, s1076=1076, s1077=1077, s1078=1078, s1079=1079, s1080=1080,
	s1081=1081, s1082=1082, s1083=1083, s1084=1084, s1085=1085, s1086=1086, s1087=1087, s1088=1088, s1089=1089, s1090=1090,
	s1091=1091, s1092=1092, s1093=1093, s1094=1094, s1095=1095, s1096=1096, s1097=1097, s1098=1098, s1099=1099, s1100=1100,
	s1101=1101, s1102=1102, s1103=1103, s1104=1104, s1105=1105, s1106=1106, s1107=1107, s1108=1108, s1109=1109, s1110=1110,
	s1111=1111, s1112=1112, s1113=1113, s1114=1114, s1115=1115, s1116=1116, s1117=1117, s1118=1118, s1119=1119, s1120=1120,
	s1121=1121, s1122=1122, s1123=1123, s1124=1124, s1125=1125, s1126=1126, s1127=1127, s1128=1128, s1129=1129, s1130=1130,
	s1131=1131, s1132=1132, s1133=1133, s1134=1134, s1135=1135, s1136=1136, s1137=1137, s1138=1138, s1139=1139, s1140=1140,
	s1141=1141, s1142=1142, s1143=1143, s1144=1144, s1145=1145, s1146=1146, s1147=1147, s1148=1148, s1149=1149, s1150=1150,
	s1151=1151, s1152=1152, s1153=1153, s1154=1154, s1155=1155, s1156=1156, s1157=1157, s1158=1158, s1159=1159, s1160=1160,
	s1161=1161, s1162=1162, s1163=1163, s1164=1164, s1165=1165, s1166=1166, s1167=1167, s1168=1168, s1169=1169, s1170=1170,
	s1171=1171, s1172=1172, s1173=1173, s1174=1174, s1175=1175, s1176=1176, s1177=1177, s1178=1178, s1179=1179, s1180=1180,
	s1181=1181, s1182=1182, s1183=1183, s1184=1184, s1185=1185, s1186=1186, s1187=1187, s1188=1188, s1189=1189, s1190=1190,
	s1191=1191, s1192=1192, s1193=1193, s1194=1194, s1195=1195, s1196=1196, s1197=1197, s1198=1198, s1199=1199, s1200=1200,
	s1201=1201, s1202=1202, s1203=1203, s1204=1204, s1205=1205, s1206=1206, s1207=1207, s1208=1208, s1209=1209, s1210=1210,
	s1211=1211, s1212=1212, s1213=1213, s1214=1214, s1215=1215, s1216=1216, s1217=1217, s1218=1218, s1219=1219, s1220=1220,
	s1221=1221, s1222=1222, s1223=1223, s1224=1224, s1225=1225, s1226=1226, s1227=1227, s1228=1228, s1229=1229, s1230=1230,
	s1231=1231, s1232=1232, s1233=1233, s1234=1234, s1235=1235, s1236=1236, s1237=1237, s1238=1238, s1239=1239, s1240=1240,
	s1241=1241, s1242=1242, s1243=1243, s1244=1244, s1245=1245, s1246=1246, s1247=1247, s1248=1248, s1249=1249, s1250=1250,
	s1251=1251, s1252=1252, s1253=1253, s1254=1254, s1255=1255, s1256=1256, s1257=1257, s1258=1258, s1259=1259, s1260=1260,
	s1261=1261, s1262=1262, s1263=1263, s1264=1264, s1265=1265, s1266=1266, s1267=1267, s1268=1268, s1269=1269, s1270=1270,
	s1271=1271, s1272=1272, s1273=1273, s1274=1274, s1275=1275, s1276=1276, s1277=1277, s1278=1278, s1279=1279, s1280=1280,
	s1281=1281, s1282=1282, s1283=1283, s1284=1284, s1285=1285, s1286=1286, s1287=1287, s1288=1288, s1289=1289, s1290=1290,
	s1291=1291, s1292=1292, s1293=1293, s1294=1294, s1295=1295, s1296=1296, s1297=1297, s1298=1298, s1299=1299, s1300=1300,
	s1301=1301, s1302=1302, s1303=1303, s1304=1304, s1305=1305, s1306=1306, s1307=1307, s1308=1308, s1309=1309, s1310=1310,
	s1311=1311, s1312=1312, s1313=1313, s1314=1314, s1315=1315, s1316=1316, s1317=1317, s1318=1318, s1319=1319, s1320=1320,
	s1321=1321, s1322=1322, s1323=1323, s1324=1324, s1325=1325, s1326=1326, s1327=1327, s1328=1328, s1329=1329, s1330=1330,
	s1331=1331, s1332=1332, s1333=1333, s1334=1334, s1335=1335, s1336=1336, s1337=1337, s1338=1338, s1339=1339, s1340=1340,
	s1341=1341, s1342=1342, s1343=1343, s1344=1344, s1345=1345, s1346=1346, s1347=1347, s1348=1348, s1349=1349, s1350=1350,
	s1351=1351, s1352=1352, s1353=1353, s1354=1354, s1355=1355, s1356=1356, s1357=1357, s1358=1358, s1359=1359, s1360=1360,
	s1361=1361, s1362=1362, s1363=1363, s1364=1364, s1365=1365, s1366=1366, s1367=1367, s1368=1368, s1369=1369, s1370=1370,
	s1371=1371, s1372=1372, s1373=1373, s1374=1374, s1375=1375, s1376=1376, s1377=1377, s1378=1378, s1379=1379, s1380=1380,
	s1381=1381, s1382=1382, s1383=1383, s1384=1384, s1385=1385, s1386=1386, s1387=1387, s1388=1388, s1389=1389, s1390=1390,
	s1391=1391, s1392=1392, s1393=1393, s1394=1394, s1395=1395, s1396=1396, s1397=1397, s1398=1398, s1399=1399, s1400=1400,
	s1401=1401, s1402=1402, s1403=1403, s1404=1404, s1405=1405, s1406=1406, s1407=1407, s1408=1408, s1409=1409, s1410=1410,
	s1411=1411, s1412=1412, s1413=1413, s1414=1414, s1415=1415, s1416=1416, s1417=1417, s1418=1418, s1419=1419, s1420=1420,
	s1421=1421, s1422=1422, s1423=1423, s1424=1424, s1425=1425, s1426=1426, s1427=1427, s1428=1428, s1429=1429, s1430=1430,
	s1431=1431, s1432=1432, s1433=1433, s1434=1434, s1435=1435, s1436=1436, s1437=1437, s1438=1438, s1439=1439, s1440=1440,
	s1441=1441, s1442=1442, s1443=1443, s1444=1444, s1445=1445, s1446=1446, s1447=1447, s1448=1448, s1449=1449, s1450=1450,
	s1451=1451, s1452=1452, s1453=1453, s1454=1454, s1455=1455, s1456=1456, s1457=1457, s1458=1458, s1459=1459, s1460=1460,
	s1461=1461, s1462=1462, s1463=1463, s1464=1464, s1465=1465, s1466=1466, s1467=1467, s1468=1468, s1469=1469, s1470=1470,
	s1471=1471, s1472=1472, s1473=1473, s1474=1474, s1475=1475, s1476=1476, s1477=1477, s1478=1478, s1479=1479, s1480=1480,
	s1481=1481, s1482=1482, s1483=1483, s1484=1484, s1485=1485, s1486=1486, s1487=1487, s1488=1488, s1489=1489, s1490=1490,
	s1491=1491, s1492=1492, s1493=1493, s1494=1494, s1495=1495, s1496=1496, s1497=1497, s1498=1498, s1499=1499, s1500=1500,
	s1501=1501, s1502=1502, s1503=1503, s1504=1504, s1505=1505, s1506=1506, s1507=1507, s1508=1508, s1509=1509, s1510=1510,
	s1511=1511, s1512=1512, s1513=1513, s1514=1514, s1515=1515, s1516=1516, s1517=1517, s1518=1518, s1519=1519, s1520=1520,
	s1521=1521, s1522=1522, s1523=1523, s1524=1524, s1525=1525, s1526=1526, s1527=1527, s1528=1528, s1529=1529, s1530=1530,
	s1531=1531, s1532=1532, s1533=1533, s1534=1534, s1535=1535, s1536=1536, s1537=1537, s1538=1538, s1539=1539, s1540=1540,
	s1541=1541, s1542=1542, s1543=1543, s1544=1544, s1545=1545, s1546=1546, s1547=1547, s1548=1548, s1549=1549, s1550=1550,
	s1551=1551, s1552=1552, s1553=1553, s1554=1554, s1555=1555, s1556=1556, s1557=1557, s1558=1558, s1559=1559, s1560=1560,
	s1561=1561, s1562=1562, s1563=1563, s1564=1564, s1565=1565, s1566=1566, s1567=1567, s1568=1568, s1569=1569, s1570=1570,
	s1571=1571, s1572=1572, s1573=1573, s1574=1574, s1575=1575, s1576=1576, s1577=1577, s1578=1578, s1579=1579, s1580=1580,
	s1581=1581, s1582=1582, s1583=1583, s1584=1584, s1585=1585, s1586=1586, s1587=1587, s1588=1588, s1589=1589, s1590=1590,
	s1591=1591, s1592=1592, s1593=1593, s1594=1594, s1595=1595, s1596=1596, s1597=1597, s1598=1598, s1599=1599, s1600=1600,
	s1601=1601, s1602=1602, s1603=1603, s1604=1604, s1605=1605, s1606=1606, s1607=1607, s1608=1608, s1609=1609, s1610=1610,
	s1611=1611, s1612=1612, s1613=1613, s1614=1614, s1615=1615, s1616=1616, s1617=1617, s1618=1618, s1619=1619, s1620=1620,
	s1621=1621, s1622=1622, s1623=1623, s1624=1624, s1625=1625, s1626=1626, s1627=1627, s1628=1628, s1629=1629, s1630=1630,
	s1631=1631, s1632=1632, s1633=1633, s1634=1634, s1635=1635, s1636=1636, s1637=1637, s1638=1638, s1639=1639, s1640=1640,
	s1641=1641, s1642=1642, s1643=1643, s1644=1644, s1645=1645, s1646=1646, s1647=1647, s1648=1648, s1649=1649, s1650=1650,
	s1651=1651, s1652=1652, s1653=1653, s1654=1654, s1655=1655, s1656=1656, s1657=1657, s1658=1658, s1659=1659, s1660=1660,
	s1661=1661, s1662=1662, s1663=1663, s1664=1664, s1665=1665, s1666=1666, s1667=1667, s1668=1668, s1669=1669, s1670=1670,
	s1671=1671, s1672=1672, s1673=1673, s1674=1674, s1675=1675, s1676=1676, s1677=1677, s1678=1678, s1679=1679, s1680=1680,
	s1681=1681, s1682=1682, s1683=1683, s1684=1684, s1685=1685, s1686=1686, s1687=1687, s1688=1688, s1689=1689, s1690=1690,
	s1691=1691, s1692=1692, s1693=1693, s1694=1694, s1695=1695, s1696=1696, s1697=1697, s1698=1698, s1699=1699, s1700=1700,
	s1701=1701, s1702=1702, s1703=1703, s1704=1704, s1705=1705, s1706=1706, s1707=1707, s1708=1708, s1709=1709, s1710=1710,
	s1711=1711, s1712=1712, s1713=1713, s1714=1714, s1715=1715, s1716=1716, s1717=1717, s1718=1718, s1719=1719, s1720=1720,
	s1721=1721, s1722=1722, s1723=1723, s1724=1724, s1725=1725, s1726=1726, s1727=1727, s1728=1728, s1729=1729, s1730=1730,
	s1731=1731, s1732=1732, s1733=1733, s1734=1734, s1735=1735, s1736=1736, s1737=1737, s1738=1738, s1739=1739, s1740=1740,
	s1741=1741, s1742=1742, s1743=1743, s1744=1744, s1745=1745, s1746=1746, s1747=1747, s1748=1748, s1749=1749, s1750=1750,
	s1751=1751, s1752=1752, s1753=1753, s1754=1754, s1755=1755, s1756=1756, s1757=1757, s1758=1758, s1759=1759, s1760=1760,
	s1761=1761, s1762=1762, s1763=1763, s1764=1764, s1765=1765, s1766=1766, s1767=1767, s1768=1768, s1769=1769, s1770=1770,
	s1771=1771, s1772=1772, s1773=1773, s1774=1774, s1775=1775, s1776=1776, s1777=1777, s1778=1778, s1779=1779, s1780=1780,
	s1781=1781, s1782=1782, s1783=1783, s1784=1784, s1785=1785, s1786=1786, s1787=1787, s1788=1788, s1789=1789, s1790=1790,
	s1791=1791, s1792=1792, s1793=1793, s1794=1794, s1795=1795, s1796=1796, s1797=1797, s1798=1798, s1799=1799, s1800=1800,
	s1801=1801, s1802=1802, s1803=1803, s1804=1804, s1805=1805, s1806=1806;
integer pr_state;
integer nx_state;

always@ ( posedge rst or negedge clk )
begin
	if ( rst == 1'b1 )
		pr_state = s1;
	else
		pr_state = nx_state;
end

always@ ( pr_state or x1 or x2 or x3 or x4 or x5 or x6 or x7 or x8 or x9 or x10 or x11 or x12 or x13 or x14 or x15 or 
	x16 or x17 or x18 or x19 or x20 or x21 or x22 or x23 or x24 or x25 or x26 or x27 or x28 or x29 or x30 or 
	x31 or x32 or x33 or x34 or x35 or x36 or x37 or x38 or x39 or x40 or x41 or x42 or x43 or x44 or x45 or 
	x46 or x47 or x48 or x49 or x50 or x51 or x52 or x53 or x54 or x55 or x56 or x57 or x58 or x59 or x60 or 
	x61 or x62 or x63 or x64 or x65 or x66 or x67 or x68 or x69 or x70)
	begin
			y1 = 1'b0;	y2 = 1'b0;	y3 = 1'b0;	y4 = 1'b0;	
			y5 = 1'b0;	y6 = 1'b0;	y7 = 1'b0;	y8 = 1'b0;	
			y9 = 1'b0;	y10 = 1'b0;	y11 = 1'b0;	y12 = 1'b0;	
			y13 = 1'b0;	y14 = 1'b0;	y15 = 1'b0;	y16 = 1'b0;	
			y17 = 1'b0;	y18 = 1'b0;	y19 = 1'b0;	y20 = 1'b0;	
			y21 = 1'b0;	y22 = 1'b0;	y23 = 1'b0;	y24 = 1'b0;	
			y25 = 1'b0;	y26 = 1'b0;	y27 = 1'b0;	y28 = 1'b0;	
			y29 = 1'b0;	y30 = 1'b0;	y31 = 1'b0;	y32 = 1'b0;	
			y33 = 1'b0;	y34 = 1'b0;	y35 = 1'b0;	y36 = 1'b0;	
			y37 = 1'b0;	y38 = 1'b0;	y39 = 1'b0;	y40 = 1'b0;	
			y41 = 1'b0;	y42 = 1'b0;	y43 = 1'b0;	y44 = 1'b0;	
			y45 = 1'b0;	y46 = 1'b0;	y47 = 1'b0;	y48 = 1'b0;	
			y49 = 1'b0;	y50 = 1'b0;	y51 = 1'b0;	y52 = 1'b0;	
			y53 = 1'b0;	y54 = 1'b0;	y55 = 1'b0;	y56 = 1'b0;	
			y57 = 1'b0;	y58 = 1'b0;	y59 = 1'b0;	y60 = 1'b0;	
			y61 = 1'b0;	y62 = 1'b0;	y63 = 1'b0;	y64 = 1'b0;	
			y65 = 1'b0;	y66 = 1'b0;	y67 = 1'b0;	y68 = 1'b0;	
			y69 = 1'b0;	y70 = 1'b0;	y71 = 1'b0;	y72 = 1'b0;	
			y73 = 1'b0;	y74 = 1'b0;	y75 = 1'b0;	y77 = 1'b0;	
			y78 = 1'b0;	y79 = 1'b0;	y80 = 1'b0;	y81 = 1'b0;	
			y84 = 1'b0;	y86 = 1'b0;	y88 = 1'b0;	y90 = 1'b0;	
			y91 = 1'b0;	y92 = 1'b0;	y93 = 1'b0;	y94 = 1'b0;	
			y95 = 1'b0;	y96 = 1'b0;	y97 = 1'b0;	y98 = 1'b0;	
			y99 = 1'b0;	y100 = 1'b0;	y102 = 1'b0;	y110 = 1'b0;	
			y112 = 1'b0;	
		case ( pr_state )
				s1 : if( x69 && x70 && x62 && x65 && x64 && x2 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y8 = 1'b1;	
							nx_state = s2;
						end
					else if( x69 && x70 && x62 && x65 && x64 && x2 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && x62 && x65 && x64 && ~x2 && x1 )
						begin
							y17 = 1'b1;	
							nx_state = s3;
						end
					else if( x69 && x70 && x62 && x65 && x64 && ~x2 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && x66 && x67 && x25 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s4;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && x66 && x67 && ~x25 && x26 && x27 )
						begin
							y14 = 1'b1;	
							nx_state = s5;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && x66 && x67 && ~x25 && x26 && ~x27 && x2 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s6;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && x66 && x67 && ~x25 && x26 && ~x27 && x2 && ~x4 && x5 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	
							nx_state = s7;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && x66 && x67 && ~x25 && x26 && ~x27 && x2 && ~x4 && ~x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && x66 && x67 && ~x25 && x26 && ~x27 && ~x2 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && x66 && x67 && ~x25 && x26 && ~x27 && ~x2 && ~x3 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && x66 && x67 && ~x25 && ~x26 && x27 && x14 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && x66 && x67 && ~x25 && ~x26 && x27 && x14 && ~x12 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && x66 && x67 && ~x25 && ~x26 && x27 && ~x14 && x15 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && x66 && x67 && ~x25 && ~x26 && x27 && ~x14 && x15 && ~x12 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && x66 && x67 && ~x25 && ~x26 && x27 && ~x14 && ~x15 && x16 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && x66 && x67 && ~x25 && ~x26 && x27 && ~x14 && ~x15 && x16 && ~x12 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && x66 && x67 && ~x25 && ~x26 && x27 && ~x14 && ~x15 && ~x16 )
						begin
							y19 = 1'b1;	
							nx_state = s13;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && x66 && x67 && ~x25 && ~x26 && ~x27 && x12 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && x66 && x67 && ~x25 && ~x26 && ~x27 && ~x12 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && x66 && ~x67 && x2 )
						begin
							y1 = 1'b1;	y26 = 1'b1;	y37 = 1'b1;	
							nx_state = s15;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && x66 && ~x67 && ~x2 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && ~x66 && x67 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && ~x66 && ~x67 && x2 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s18;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && ~x66 && ~x67 && ~x2 && x3 && x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s19;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && ~x66 && ~x67 && ~x2 && x3 && ~x6 && x7 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && ~x66 && ~x67 && ~x2 && x3 && ~x6 && ~x7 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s19;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && x1 && ~x66 && ~x67 && ~x2 && ~x3 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	
							nx_state = s20;
						end
					else if( x69 && x70 && x62 && x65 && ~x64 && ~x1 && x67 )
						nx_state = s1;
					else if( x69 && x70 && x62 && x65 && ~x64 && ~x1 && ~x67 && x66 )
						nx_state = s1;
					else if( x69 && x70 && x62 && x65 && ~x64 && ~x1 && ~x67 && ~x66 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && x67 && x2 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && x67 && x2 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && x67 && ~x2 && x32 && x33 && x1 )
						begin
							y15 = 1'b1;	
							nx_state = s22;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && x67 && ~x2 && x32 && x33 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && x67 && ~x2 && x32 && ~x33 && x1 )
						begin
							y3 = 1'b1;	y52 = 1'b1;	
							nx_state = s23;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && x67 && ~x2 && x32 && ~x33 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && x67 && ~x2 && ~x32 && x1 )
						begin
							y3 = 1'b1;	y52 = 1'b1;	
							nx_state = s23;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && x67 && ~x2 && ~x32 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && x12 && x11 && x13 && x1 && x3 && x6 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s24;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && x12 && x11 && x13 && x1 && x3 && ~x6 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && x12 && x11 && x13 && x1 && ~x3 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && x12 && x11 && x13 && ~x1 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s33;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && x12 && x11 && ~x13 && x5 )
						begin
							y5 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s26;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && x12 && x11 && ~x13 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && x12 && ~x11 && x8 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s27;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && x12 && ~x11 && ~x8 && x5 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s28;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && x12 && ~x11 && ~x8 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && ~x12 && x11 && x13 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s29;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && ~x12 && x11 && ~x13 && x14 && x7 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s27;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && ~x12 && x11 && ~x13 && x14 && ~x7 && x1 && x5 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s28;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && ~x12 && x11 && ~x13 && x14 && ~x7 && x1 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && ~x12 && x11 && ~x13 && x14 && ~x7 && ~x1 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s33;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && ~x12 && x11 && ~x13 && ~x14 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s30;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && ~x12 && ~x11 && x14 && x1 && x5 && x13 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s29;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && ~x12 && ~x11 && x14 && x1 && x5 && ~x13 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s28;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && ~x12 && ~x11 && x14 && x1 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && ~x12 && ~x11 && x14 && ~x1 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s33;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && ~x12 && ~x11 && ~x14 && x13 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s31;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && ~x12 && ~x11 && ~x14 && ~x13 && x1 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && x10 && ~x12 && ~x11 && ~x14 && ~x13 && ~x1 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s33;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && x64 && ~x67 && ~x10 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s33;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && ~x64 && x67 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && ~x64 && ~x67 && x6 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s35;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && ~x64 && ~x67 && ~x6 && x7 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && x62 && ~x65 && x66 && ~x64 && ~x67 && ~x6 && ~x7 )
						begin
							y3 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s37;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && x64 && x67 && x2 && x1 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							nx_state = s38;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && x64 && x67 && x2 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x65 && ~x66 && x64 && x67 && ~x2 && x1 )
						begin
							y22 = 1'b1;	
							nx_state = s39;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && x64 && x67 && ~x2 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x65 && ~x66 && x64 && ~x67 && x13 && x10 && x1 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && x64 && ~x67 && x13 && x10 && ~x1 && x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && x64 && ~x67 && x13 && x10 && ~x1 && ~x2 && x15 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && x64 && ~x67 && x13 && x10 && ~x1 && ~x2 && ~x15 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && x64 && ~x67 && x13 && ~x10 && x1 && x2 && x3 && x15 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x65 && ~x66 && x64 && ~x67 && x13 && ~x10 && x1 && x2 && x3 && ~x15 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && x64 && ~x67 && x13 && ~x10 && x1 && x2 && ~x3 && x4 && x5 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && x64 && ~x67 && x13 && ~x10 && x1 && x2 && ~x3 && x4 && ~x5 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && x64 && ~x67 && x13 && ~x10 && x1 && x2 && ~x3 && ~x4 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && x64 && ~x67 && x13 && ~x10 && x1 && ~x2 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s45;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && x64 && ~x67 && x13 && ~x10 && ~x1 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && x64 && ~x67 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s45;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && x64 && ~x67 && ~x13 && ~x12 && x10 && x1 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && x64 && ~x67 && ~x13 && ~x12 && x10 && ~x1 && x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && x64 && ~x67 && ~x13 && ~x12 && x10 && ~x1 && ~x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && x64 && ~x67 && ~x13 && ~x12 && ~x10 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s45;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && x67 && x2 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s46;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && x67 && x2 && ~x1 )
						nx_state = s47;
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && x67 && ~x2 && x1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && x67 && ~x2 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && x18 && x17 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && x18 && x17 && ~x1 && x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && x18 && x17 && ~x1 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && x18 && ~x17 && x19 && x1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && x18 && ~x17 && x19 && ~x1 && x4 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && x18 && ~x17 && x19 && ~x1 && ~x4 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	
							nx_state = s20;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && x18 && ~x17 && ~x19 && x1 && x2 && x4 && x5 && x3 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && x18 && ~x17 && ~x19 && x1 && x2 && x4 && x5 && ~x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && x18 && ~x17 && ~x19 && x1 && x2 && x4 && ~x5 && x3 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && x18 && ~x17 && ~x19 && x1 && x2 && x4 && ~x5 && ~x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && x18 && ~x17 && ~x19 && x1 && x2 && ~x4 && x3 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	
							nx_state = s20;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && x18 && ~x17 && ~x19 && x1 && x2 && ~x4 && ~x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && x18 && ~x17 && ~x19 && x1 && ~x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && x18 && ~x17 && ~x19 && ~x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && ~x18 && x17 && x19 && x1 && x10 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && ~x18 && x17 && x19 && x1 && ~x10 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	
							nx_state = s20;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && ~x18 && x17 && x19 && ~x1 && x6 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && ~x18 && x17 && x19 && ~x1 && ~x6 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && ~x18 && x17 && ~x19 && x1 && x2 && x4 && x5 && x3 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && ~x18 && x17 && ~x19 && x1 && x2 && x4 && x5 && ~x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && ~x18 && x17 && ~x19 && x1 && x2 && x4 && ~x5 && x3 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && ~x18 && x17 && ~x19 && x1 && x2 && x4 && ~x5 && ~x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && ~x18 && x17 && ~x19 && x1 && x2 && ~x4 && x3 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	
							nx_state = s20;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && ~x18 && x17 && ~x19 && x1 && x2 && ~x4 && ~x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && ~x18 && x17 && ~x19 && x1 && ~x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && ~x18 && x17 && ~x19 && ~x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x66 && ~x64 && ~x67 && ~x18 && ~x17 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x69 && x70 && ~x62 && x63 && x66 && x65 && x67 && x64 && x13 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							nx_state = s52;
						end
					else if( x69 && x70 && ~x62 && x63 && x66 && x65 && x67 && x64 && x13 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x66 && x65 && x67 && x64 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s53;
						end
					else if( x69 && x70 && ~x62 && x63 && x66 && x65 && x67 && x64 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x66 && x65 && x67 && ~x64 && x1 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x70 && ~x62 && x63 && x66 && x65 && x67 && ~x64 && ~x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && x70 && ~x62 && x63 && x66 && x65 && ~x67 && x64 && x9 && x8 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x66 && x65 && ~x67 && x64 && x9 && ~x8 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s54;
						end
					else if( x69 && x70 && ~x62 && x63 && x66 && x65 && ~x67 && x64 && ~x9 && x8 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x66 && x65 && ~x67 && x64 && ~x9 && ~x8 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y19 = 1'b1;	
							nx_state = s55;
						end
					else if( x69 && x70 && ~x62 && x63 && x66 && x65 && ~x67 && ~x64 && x6 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && x70 && ~x62 && x63 && x66 && x65 && ~x67 && ~x64 && ~x6 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x66 && ~x65 && x64 && x2 && x67 && x1 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x62 && x63 && x66 && ~x65 && x64 && x2 && x67 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x66 && ~x65 && x64 && x2 && ~x67 && x1 )
						begin
							y2 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							nx_state = s56;
						end
					else if( x69 && x70 && ~x62 && x63 && x66 && ~x65 && x64 && x2 && ~x67 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x66 && ~x65 && x64 && ~x2 && x67 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( x69 && x70 && ~x62 && x63 && x66 && ~x65 && x64 && ~x2 && x67 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x66 && ~x65 && x64 && ~x2 && ~x67 && x1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s6;
						end
					else if( x69 && x70 && ~x62 && x63 && x66 && ~x65 && x64 && ~x2 && ~x67 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x66 && ~x65 && ~x64 && x1 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && x70 && ~x62 && x63 && x66 && ~x65 && ~x64 && x1 && ~x2 && x67 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s57;
						end
					else if( x69 && x70 && ~x62 && x63 && x66 && ~x65 && ~x64 && x1 && ~x2 && ~x67 && x5 && x3 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x66 && ~x65 && ~x64 && x1 && ~x2 && ~x67 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x70 && ~x62 && x63 && x66 && ~x65 && ~x64 && x1 && ~x2 && ~x67 && ~x5 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	
							nx_state = s7;
						end
					else if( x69 && x70 && ~x62 && x63 && x66 && ~x65 && ~x64 && ~x1 && x67 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x66 && ~x65 && ~x64 && ~x1 && ~x67 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && x67 && x15 && x16 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && x67 && x15 && x16 && ~x5 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s60;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && x67 && x15 && x16 && ~x5 && ~x6 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y22 = 1'b1;	
							nx_state = s61;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && x67 && x15 && ~x16 && x1 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && x67 && x15 && ~x16 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && x67 && ~x15 && x1 && x16 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && x67 && ~x15 && x1 && ~x16 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && x67 && ~x15 && ~x1 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && x17 && x1 && x18 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s45;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && x17 && x1 && ~x18 && x15 && x10 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && x17 && x1 && ~x18 && x15 && ~x10 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && x17 && x1 && ~x18 && ~x15 && x2 && x4 && x5 && x3 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && x17 && x1 && ~x18 && ~x15 && x2 && x4 && x5 && ~x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && x17 && x1 && ~x18 && ~x15 && x2 && x4 && ~x5 && x3 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && x17 && x1 && ~x18 && ~x15 && x2 && x4 && ~x5 && ~x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && x17 && x1 && ~x18 && ~x15 && x2 && ~x4 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && x17 && x1 && ~x18 && ~x15 && x2 && ~x4 && ~x3 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && x17 && x1 && ~x18 && ~x15 && ~x2 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s45;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && x17 && ~x1 && x18 && x2 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && x17 && ~x1 && x18 && ~x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && x17 && ~x1 && ~x18 && x15 && x6 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s45;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && x17 && ~x1 && ~x18 && x15 && ~x6 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && x17 && ~x1 && ~x18 && ~x15 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && ~x17 && x18 && x15 && x1 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && ~x17 && x18 && x15 && ~x1 && x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && ~x17 && x18 && x15 && ~x1 && ~x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && ~x17 && x18 && ~x15 && x1 && x2 && x4 && x5 && x3 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && ~x17 && x18 && ~x15 && x1 && x2 && x4 && x5 && ~x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && ~x17 && x18 && ~x15 && x1 && x2 && x4 && ~x5 && x3 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && ~x17 && x18 && ~x15 && x1 && x2 && x4 && ~x5 && ~x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && ~x17 && x18 && ~x15 && x1 && x2 && ~x4 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && ~x17 && x18 && ~x15 && x1 && x2 && ~x4 && ~x3 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && ~x17 && x18 && ~x15 && x1 && ~x2 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s45;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && ~x17 && x18 && ~x15 && ~x1 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && x64 && ~x67 && ~x17 && ~x18 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s45;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && ~x64 && x67 && x15 && x1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && ~x64 && x67 && x15 && ~x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && ~x64 && x67 && ~x15 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && ~x64 && ~x67 && x2 && x1 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && ~x64 && ~x67 && x2 && ~x1 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && x65 && ~x64 && ~x67 && ~x2 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && x67 && x11 && x14 )
						begin
							y5 = 1'b1;	
							nx_state = s64;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && x67 && x11 && ~x14 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s65;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && x67 && ~x11 && x10 && x1 && x14 && x3 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s66;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && x67 && ~x11 && x10 && x1 && x14 && x3 && ~x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && x67 && ~x11 && x10 && x1 && x14 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && x67 && ~x11 && x10 && x1 && ~x14 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s65;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && x67 && ~x11 && x10 && x1 && ~x14 && ~x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && x67 && ~x11 && x10 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y4 = 1'b1;	
							nx_state = s71;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && x67 && ~x11 && ~x10 && x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s68;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && x67 && ~x11 && ~x10 && ~x14 && x1 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && x67 && ~x11 && ~x10 && ~x14 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y4 = 1'b1;	
							nx_state = s71;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && x15 && x10 && x1 && x14 && x3 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s66;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && x15 && x10 && x1 && x14 && x3 && ~x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && x15 && x10 && x1 && x14 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && x15 && x10 && x1 && ~x14 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s65;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && x15 && x10 && x1 && ~x14 && ~x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && x15 && x10 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y4 = 1'b1;	
							nx_state = s71;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && x15 && ~x10 && x14 )
						begin
							y5 = 1'b1;	
							nx_state = s64;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && x15 && ~x10 && ~x14 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s65;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && ~x15 && x11 && x14 && x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && ~x15 && x11 && x14 && ~x8 && x5 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && ~x15 && x11 && x14 && ~x8 && ~x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && ~x15 && x11 && ~x14 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && ~x15 && x11 && ~x14 && ~x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && ~x15 && ~x11 && x14 && x10 && x7 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && ~x15 && ~x11 && x14 && x10 && ~x7 && x1 && x5 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && ~x15 && ~x11 && x14 && x10 && ~x7 && x1 && ~x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && ~x15 && ~x11 && x14 && x10 && ~x7 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y4 = 1'b1;	
							nx_state = s71;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && ~x15 && ~x11 && x14 && ~x10 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s68;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && ~x15 && ~x11 && ~x14 && x1 && x10 && x5 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && ~x15 && ~x11 && ~x14 && x1 && x10 && ~x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && ~x15 && ~x11 && ~x14 && x1 && ~x10 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && x13 && ~x67 && ~x15 && ~x11 && ~x14 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y4 = 1'b1;	
							nx_state = s71;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && x64 && ~x13 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y4 = 1'b1;	
							nx_state = s71;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && ~x64 && x67 && x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s57;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && ~x64 && x67 && x15 && ~x14 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && ~x64 && x67 && ~x15 && x14 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && ~x64 && x67 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && ~x64 && ~x67 && x18 && x14 && x23 && x22 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y5 = 1'b1;	
							y22 = 1'b1;	y23 = 1'b1;	
							nx_state = s72;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && ~x64 && ~x67 && x18 && x14 && x23 && ~x22 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y5 = 1'b1;	
							y22 = 1'b1;	y23 = 1'b1;	
							nx_state = s73;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && ~x64 && ~x67 && x18 && x14 && ~x23 && x22 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y5 = 1'b1;	
							y22 = 1'b1;	y23 = 1'b1;	
							nx_state = s73;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && ~x64 && ~x67 && x18 && x14 && ~x23 && ~x22 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y5 = 1'b1;	
							y22 = 1'b1;	y23 = 1'b1;	
							nx_state = s72;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && ~x64 && ~x67 && x18 && ~x14 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x66 && ~x65 && ~x64 && ~x67 && ~x18 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x2 && x64 && x65 && x66 && x67 && x1 )
						begin
							y35 = 1'b1;	y36 = 1'b1;	
							nx_state = s74;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x2 && x64 && x65 && x66 && x67 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x2 && x64 && x65 && x66 && ~x67 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x2 && x64 && x65 && x66 && ~x67 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x2 && x64 && x65 && ~x66 && x67 && x1 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s76;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x2 && x64 && x65 && ~x66 && x67 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x2 && x64 && x65 && ~x66 && ~x67 && x1 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x2 && x64 && x65 && ~x66 && ~x67 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x2 && x64 && ~x65 && x66 && x67 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s57;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x2 && x64 && ~x65 && x66 && x67 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x2 && x64 && ~x65 && x66 && ~x67 && x1 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x2 && x64 && ~x65 && x66 && ~x67 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x2 && x64 && ~x65 && ~x66 && x67 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y20 = 1'b1;	y38 = 1'b1;	
							nx_state = s79;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x2 && x64 && ~x65 && ~x66 && x67 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x2 && x64 && ~x65 && ~x66 && ~x67 && x1 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y13 = 1'b1;	
							y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s80;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x2 && x64 && ~x65 && ~x66 && ~x67 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x2 && ~x64 && x65 && x66 && x67 && x1 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s81;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x2 && ~x64 && x65 && x66 && x67 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x2 && ~x64 && x65 && x66 && ~x67 && x1 )
						begin
							y7 = 1'b1;	
							nx_state = s82;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x2 && ~x64 && x65 && x66 && ~x67 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x2 && ~x64 && x65 && ~x66 && x67 && x1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y5 = 1'b1;	
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s83;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x2 && ~x64 && x65 && ~x66 && x67 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x2 && ~x64 && x65 && ~x66 && ~x67 && x1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y25 = 1'b1;	
							nx_state = s84;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x2 && ~x64 && x65 && ~x66 && ~x67 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x2 && ~x64 && ~x65 && x67 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s57;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x2 && ~x64 && ~x65 && x67 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x2 && ~x64 && ~x65 && ~x67 && x66 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s57;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x2 && ~x64 && ~x65 && ~x67 && x66 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x2 && ~x64 && ~x65 && ~x67 && ~x66 && x1 )
						begin
							y7 = 1'b1;	
							nx_state = s82;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x2 && ~x64 && ~x65 && ~x67 && ~x66 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x2 && x66 && x67 && x65 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x2 && x66 && x67 && x65 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x2 && x66 && x67 && ~x65 && x64 && x1 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y42 = 1'b1;	
							nx_state = s85;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x2 && x66 && x67 && ~x65 && x64 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x2 && x66 && x67 && ~x65 && ~x64 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x2 && x66 && x67 && ~x65 && ~x64 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x2 && x66 && ~x67 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x2 && x66 && ~x67 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x2 && ~x66 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x2 && ~x66 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && x65 && x22 && x5 && x21 && x1 )
						begin
							y10 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s86;
						end
					else if( x69 && ~x70 && x67 && x66 && x65 && x22 && x5 && x21 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && x65 && x22 && x5 && ~x21 && x1 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( x69 && ~x70 && x67 && x66 && x65 && x22 && x5 && ~x21 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && x65 && x22 && ~x5 && x6 && x1 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x67 && x66 && x65 && x22 && ~x5 && x6 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && x65 && x22 && ~x5 && ~x6 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s57;
						end
					else if( x69 && ~x70 && x67 && x66 && x65 && x22 && ~x5 && ~x6 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && x65 && ~x22 && x4 && x17 && x23 && x1 )
						begin
							y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s1;
						end
					else if( x69 && ~x70 && x67 && x66 && x65 && ~x22 && x4 && x17 && x23 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && x65 && ~x22 && x4 && x17 && ~x23 && x1 )
						begin
							y3 = 1'b1;	y11 = 1'b1;	
							nx_state = s89;
						end
					else if( x69 && ~x70 && x67 && x66 && x65 && ~x22 && x4 && x17 && ~x23 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && x65 && ~x22 && x4 && ~x17 && x23 && x1 )
						begin
							y3 = 1'b1;	y11 = 1'b1;	
							nx_state = s89;
						end
					else if( x69 && ~x70 && x67 && x66 && x65 && ~x22 && x4 && ~x17 && x23 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && x65 && ~x22 && x4 && ~x17 && ~x23 && x1 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x67 && x66 && x65 && ~x22 && x4 && ~x17 && ~x23 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && x65 && ~x22 && ~x4 && x5 && x23 && x1 )
						begin
							y11 = 1'b1;	
							nx_state = s91;
						end
					else if( x69 && ~x70 && x67 && x66 && x65 && ~x22 && ~x4 && x5 && x23 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && x65 && ~x22 && ~x4 && x5 && ~x23 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y10 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s92;
						end
					else if( x69 && ~x70 && x67 && x66 && x65 && ~x22 && ~x4 && x5 && ~x23 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && x65 && ~x22 && ~x4 && ~x5 && x23 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( x69 && ~x70 && x67 && x66 && x65 && ~x22 && ~x4 && ~x5 && x23 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && x65 && ~x22 && ~x4 && ~x5 && ~x23 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s57;
						end
					else if( x69 && ~x70 && x67 && x66 && x65 && ~x22 && ~x4 && ~x5 && ~x23 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && ~x65 && x68 && x1 && x21 && x6 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && x68 && x1 && x21 && ~x6 && x5 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && x68 && x1 && x21 && ~x6 && x5 && ~x18 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && x68 && x1 && x21 && ~x6 && ~x5 && x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && x68 && x1 && x21 && ~x6 && ~x5 && ~x4 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s97;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && x68 && x1 && ~x21 && x4 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && x68 && x1 && ~x21 && ~x4 && x5 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && x68 && x1 && ~x21 && ~x4 && x5 && ~x18 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && x68 && x1 && ~x21 && ~x4 && ~x5 && x6 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && x68 && x1 && ~x21 && ~x4 && ~x5 && ~x6 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s97;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && x68 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && x62 && x5 && x51 && x1 )
						begin
							y17 = 1'b1;	
							nx_state = s98;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && x62 && x5 && x51 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && x62 && x5 && ~x51 && x1 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s99;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && x62 && x5 && ~x51 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && x62 && ~x5 && x2 && x1 )
						begin
							y14 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s100;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && x62 && ~x5 && x2 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && x62 && ~x5 && ~x2 && x1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s101;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && x62 && ~x5 && ~x2 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && x64 && x4 && x5 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s102;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && x64 && x4 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && x64 && ~x4 && x5 && x3 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && x64 && ~x4 && x5 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && x64 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && ~x64 && x2 && x1 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && ~x64 && x2 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && ~x64 && ~x2 && x4 && x1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && ~x64 && ~x2 && x4 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && ~x64 && ~x2 && ~x4 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && ~x64 && ~x2 && ~x4 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && x64 && x5 && x17 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && x64 && x5 && x17 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && x64 && x5 && ~x17 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && x64 && x5 && ~x17 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && x64 && ~x5 && x2 && x1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && x64 && ~x5 && x2 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && x64 && ~x5 && ~x2 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && x64 && ~x5 && ~x2 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && ~x64 && x5 && x18 && x1 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && ~x64 && x5 && x18 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && ~x64 && x5 && ~x18 && x1 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && ~x64 && x5 && ~x18 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && ~x64 && ~x5 && x2 && x1 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && ~x64 && ~x5 && x2 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && ~x64 && ~x5 && ~x2 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x69 && ~x70 && x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && ~x64 && ~x5 && ~x2 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && x21 && x7 && x1 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && x21 && x7 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && x21 && ~x7 && x11 && x2 && x1 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s107;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && x21 && ~x7 && x11 && x2 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && x21 && ~x7 && x11 && ~x2 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && x21 && ~x7 && x11 && ~x2 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && x21 && ~x7 && ~x11 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && x21 && ~x7 && ~x11 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && x22 && x23 && x9 && x1 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && x22 && x23 && x9 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && x22 && x23 && ~x9 && x2 && x3 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s110;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && x22 && x23 && ~x9 && x2 && x3 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && x22 && x23 && ~x9 && x2 && ~x3 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && x22 && x23 && ~x9 && x2 && ~x3 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && x22 && x23 && ~x9 && ~x2 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s111;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && x22 && x23 && ~x9 && ~x2 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && x22 && ~x23 && x4 && x7 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && x22 && ~x23 && x4 && ~x7 && x2 && x1 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s112;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && x22 && ~x23 && x4 && ~x7 && x2 && ~x1 )
						begin
							y3 = 1'b1;	y12 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s113;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && x22 && ~x23 && x4 && ~x7 && ~x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s114;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && x22 && ~x23 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && x23 && x7 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && x23 && x7 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && x23 && ~x7 && x2 && x8 && x1 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s115;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && x23 && ~x7 && x2 && x8 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && x23 && ~x7 && x2 && ~x8 && x1 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s112;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && x23 && ~x7 && x2 && ~x8 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && x23 && ~x7 && ~x2 && x1 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && x23 && ~x7 && ~x2 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && ~x23 && x9 && x1 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && ~x23 && x9 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && ~x23 && ~x9 && x2 && x3 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s110;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && ~x23 && ~x9 && x2 && x3 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && ~x23 && ~x9 && x2 && ~x3 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && ~x23 && ~x9 && x2 && ~x3 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && ~x23 && ~x9 && ~x2 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s111;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && ~x23 && ~x9 && ~x2 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && x65 && ~x68 && x9 && x1 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	y12 = 1'b1;	
							nx_state = s116;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && ~x68 && x9 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && x65 && ~x68 && ~x9 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s117;
						end
					else if( x69 && ~x70 && x67 && ~x66 && x65 && ~x68 && ~x9 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && x20 && x4 && x19 && x2 )
						nx_state = s118;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && x20 && x4 && x19 && ~x2 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && x20 && x4 && ~x19 && x2 )
						nx_state = s47;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && x20 && x4 && ~x19 && ~x2 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && x20 && ~x4 && x3 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && x20 && ~x4 && x3 && ~x2 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && x20 && ~x4 && ~x3 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && x20 && ~x4 && ~x3 && ~x2 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && ~x20 && x21 && x4 && x19 && x1 )
						begin
							y3 = 1'b1;	y20 = 1'b1;	
							nx_state = s120;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && ~x20 && x21 && x4 && x19 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && ~x20 && x21 && x4 && ~x19 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && ~x20 && x21 && x4 && ~x19 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && ~x20 && x21 && ~x4 && x5 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && ~x20 && x21 && ~x4 && x5 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && ~x20 && x21 && ~x4 && ~x5 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && ~x20 && x21 && ~x4 && ~x5 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x5 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x5 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x5 && x4 && x1 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y21 = 1'b1;	
							nx_state = s121;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x5 && x4 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x5 && ~x4 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x5 && ~x4 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && x24 && x26 && x6 && x1 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s122;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && x24 && x26 && x6 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && x24 && x26 && ~x6 && x5 && x1 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && x24 && x26 && ~x6 && x5 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && x24 && x26 && ~x6 && ~x5 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && x24 && x26 && ~x6 && ~x5 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && x24 && ~x26 && x5 && x18 && x1 )
						begin
							y14 = 1'b1;	
							nx_state = s124;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && x24 && ~x26 && x5 && x18 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && x24 && ~x26 && x5 && ~x18 && x1 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && x24 && ~x26 && x5 && ~x18 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && x24 && ~x26 && ~x5 && x2 && x1 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s126;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && x24 && ~x26 && ~x5 && x2 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && x24 && ~x26 && ~x5 && ~x2 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && x24 && ~x26 && ~x5 && ~x2 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && x26 && x6 && x2 && x17 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s126;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && x26 && x6 && x2 && ~x17 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s122;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && x26 && x6 && ~x2 && x5 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s35;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && x26 && x6 && ~x2 && ~x5 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s101;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && x26 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x3 && x17 && x1 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x3 && x17 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x3 && ~x17 && x1 )
						begin
							y14 = 1'b1;	
							nx_state = s124;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x3 && ~x17 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && ~x3 && x4 && x1 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && ~x3 && x4 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && ~x3 && ~x4 && x1 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && ~x3 && ~x4 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && x6 && x1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && x6 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && ~x6 && x5 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && ~x6 && x5 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && ~x6 && ~x5 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && ~x6 && ~x5 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && ~x26 && x6 && x19 && x1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && ~x26 && x6 && x19 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && ~x26 && x6 && ~x19 && x1 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && ~x26 && x6 && ~x19 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && ~x26 && ~x6 && x2 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && ~x26 && ~x6 && x2 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && ~x26 && ~x6 && ~x2 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( x69 && ~x70 && x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && ~x26 && ~x6 && ~x2 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && x68 && x1 && x21 && x20 && x3 && x19 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && x68 && x1 && x21 && x20 && x3 && ~x19 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s129;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && x68 && x1 && x21 && x20 && ~x3 && x4 )
						begin
							y22 = 1'b1;	
							nx_state = s130;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && x68 && x1 && x21 && x20 && ~x3 && ~x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && x68 && x1 && x21 && ~x20 && x6 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s130;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && x68 && x1 && x21 && ~x20 && x6 && ~x17 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s131;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && x68 && x1 && x21 && ~x20 && ~x6 && x4 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s132;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && x68 && x1 && x21 && ~x20 && ~x6 && ~x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && x68 && x1 && ~x21 && x6 && x20 && x17 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && x68 && x1 && ~x21 && x6 && x20 && ~x17 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	
							nx_state = s133;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && x68 && x1 && ~x21 && x6 && ~x20 && x17 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	
							nx_state = s133;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && x68 && x1 && ~x21 && x6 && ~x20 && ~x17 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && x68 && x1 && ~x21 && ~x6 && x5 )
						begin
							y22 = 1'b1;	
							nx_state = s130;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && x68 && x1 && ~x21 && ~x6 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && x68 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && x60 && x5 && x4 && x17 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && x60 && x5 && x4 && ~x17 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s135;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && x60 && x5 && ~x4 && x6 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y24 = 1'b1;	
							nx_state = s136;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && x60 && x5 && ~x4 && ~x6 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && x60 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && x62 && x59 && x19 && x1 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && x62 && x59 && x19 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && x62 && x59 && ~x19 && x1 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && x62 && x59 && ~x19 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && x62 && ~x59 && x6 && x1 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s139;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && x62 && ~x59 && x6 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && x62 && ~x59 && ~x6 && x1 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && x62 && ~x59 && ~x6 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && ~x62 && x3 && x17 && x1 )
						nx_state = s141;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && ~x62 && x3 && x17 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && ~x62 && x3 && ~x17 && x1 )
						nx_state = s142;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && ~x62 && x3 && ~x17 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && ~x62 && ~x3 && x6 && x1 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && ~x62 && ~x3 && x6 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && ~x62 && ~x3 && ~x6 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && ~x62 && ~x3 && ~x6 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && x60 && x3 && x17 && x1 )
						nx_state = s141;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && x60 && x3 && x17 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && x60 && x3 && ~x17 && x1 )
						nx_state = s142;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && x60 && x3 && ~x17 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && x60 && ~x3 && x6 && x1 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && x60 && ~x3 && x6 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && x60 && ~x3 && ~x6 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && x60 && ~x3 && ~x6 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && x62 && x3 && x1 )
						nx_state = s142;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && x62 && x3 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && x62 && ~x3 && x5 && x1 )
						nx_state = s143;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && x62 && ~x3 && x5 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && x62 && ~x3 && ~x5 && x15 && x16 && x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && x62 && ~x3 && ~x5 && x15 && x16 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && x62 && ~x3 && ~x5 && x15 && ~x16 && x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && x62 && ~x3 && ~x5 && x15 && ~x16 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && x62 && ~x3 && ~x5 && ~x15 && x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && x62 && ~x3 && ~x5 && ~x15 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && ~x62 && x6 && x1 )
						nx_state = s142;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && ~x62 && x6 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && ~x62 && ~x6 && x2 && x1 )
						nx_state = s143;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && ~x62 && ~x6 && x2 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && ~x62 && ~x6 && ~x2 && x1 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x69 && ~x70 && ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && ~x62 && ~x6 && ~x2 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && x21 && x68 && x3 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && x21 && x68 && ~x3 && x18 && x19 )
						begin
							y25 = 1'b1;	y26 = 1'b1;	
							nx_state = s1;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && x21 && x68 && ~x3 && x18 && ~x19 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && x21 && x68 && ~x3 && ~x18 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s149;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && x21 && ~x68 && x6 && x17 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && x21 && ~x68 && x6 && ~x17 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s150;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && x21 && ~x68 && ~x6 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s151;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && x21 && ~x68 && ~x6 && ~x2 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && ~x21 && x22 && x68 && x3 )
						begin
							y8 = 1'b1;	y18 = 1'b1;	
							nx_state = s152;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x3 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && x23 && x5 && x19 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && x23 && x5 && ~x19 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y13 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s1;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && x23 && ~x5 && x6 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && x23 && ~x5 && ~x6 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s57;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && ~x23 && x4 && x17 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && ~x23 && x4 && ~x17 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && ~x23 && ~x4 && x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s57;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && ~x23 && ~x4 && ~x5 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && ~x21 && ~x22 && x68 && x9 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s107;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && ~x21 && ~x22 && x68 && ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x5 && x17 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x5 && ~x17 && x23 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x5 && ~x17 && ~x23 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && ~x5 && x6 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && ~x5 && ~x6 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s57;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && x22 && x19 && x20 && x21 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && x22 && x19 && x20 && ~x21 && x68 && x3 )
						begin
							y25 = 1'b1;	y26 = 1'b1;	
							nx_state = s1;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && x22 && x19 && x20 && ~x21 && x68 && ~x3 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && x22 && x19 && x20 && ~x21 && ~x68 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && x22 && x19 && ~x20 && x21 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && x22 && x19 && ~x20 && ~x21 && x68 && x3 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && x22 && x19 && ~x20 && ~x21 && x68 && ~x3 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && x22 && x19 && ~x20 && ~x21 && ~x68 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && x22 && ~x19 && x21 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && x22 && ~x19 && ~x21 && x68 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && x22 && ~x19 && ~x21 && x68 && ~x3 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && x22 && ~x19 && ~x21 && ~x68 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && x21 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && x17 && x10 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && x17 && ~x10 && x68 && x16 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && x17 && ~x10 && x68 && ~x16 && x15 && x14 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && x17 && ~x10 && x68 && ~x16 && x15 && ~x14 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && x17 && ~x10 && x68 && ~x16 && x15 && ~x14 && ~x3 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && x17 && ~x10 && x68 && ~x16 && ~x15 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && x17 && ~x10 && x68 && ~x16 && ~x15 && ~x3 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && x17 && ~x10 && ~x68 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && x14 && x68 && x16 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && x14 && x68 && x16 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && x14 && x68 && x16 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && x14 && x68 && ~x16 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && x14 && ~x68 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && x15 && x16 && x10 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && x15 && x16 && ~x10 && x68 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && x15 && x16 && ~x10 && x68 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && x15 && x16 && ~x10 && x68 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && x15 && x16 && ~x10 && x68 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && x15 && x16 && ~x10 && ~x68 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && x15 && ~x16 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && ~x15 && x68 && x16 && x10 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && ~x15 && x68 && x16 && ~x10 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && ~x15 && x68 && x16 && ~x10 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && ~x15 && x68 && x16 && ~x10 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && ~x15 && x68 && ~x16 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && ~x15 && ~x68 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && x68 && x10 && x1 )
						begin
							y28 = 1'b1;	y29 = 1'b1;	
							nx_state = s159;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && x68 && x10 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && x68 && ~x10 && x1 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && x68 && ~x10 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && x21 && x4 && x20 && x1 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && x21 && x4 && x20 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && x21 && x4 && ~x20 && x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && x21 && x4 && ~x20 && ~x18 && x1 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && x21 && x4 && ~x20 && ~x18 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && x21 && ~x4 && x3 && x1 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && x21 && ~x4 && x3 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && x21 && ~x4 && ~x3 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && x21 && ~x4 && ~x3 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && x2 && x20 && x23 && x1 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s161;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && x2 && x20 && x23 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && x2 && x20 && ~x23 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && x2 && ~x20 && x23 && x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && x2 && ~x20 && x23 && ~x19 && x1 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && x2 && ~x20 && x23 && ~x19 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && x2 && ~x20 && ~x23 && x4 && x19 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s161;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && x2 && ~x20 && ~x23 && x4 && ~x19 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && x2 && ~x20 && ~x23 && ~x4 && x3 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && x2 && ~x20 && ~x23 && ~x4 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x2 && x3 && x23 && x1 )
						begin
							y31 = 1'b1;	
							nx_state = s164;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x2 && x3 && x23 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x2 && x3 && ~x23 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x2 && ~x3 && x23 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x2 && ~x3 && x23 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x2 && ~x3 && ~x23 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && x19 && x23 && x1 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && x19 && x23 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && x19 && ~x23 && x1 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							nx_state = s165;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && x19 && ~x23 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && x4 && x23 && x18 && x1 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && x4 && x23 && x18 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && x4 && x23 && ~x18 && x1 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							nx_state = s165;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && x4 && x23 && ~x18 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && x4 && ~x23 && x20 && x1 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s166;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && x4 && ~x23 && x20 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && x4 && ~x23 && ~x20 && x1 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && x4 && ~x23 && ~x20 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && ~x4 && x3 && x23 && x1 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && ~x4 && x3 && x23 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && ~x4 && x3 && ~x23 && x1 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s161;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && ~x4 && x3 && ~x23 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && ~x4 && ~x3 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && ~x4 && ~x3 && ~x1 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && x21 && x68 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && x21 && x68 && ~x6 && x10 && x11 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s168;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && x21 && x68 && ~x6 && x10 && ~x11 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && x21 && x68 && ~x6 && ~x10 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && x21 && ~x68 && x10 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s169;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && x21 && ~x68 && ~x10 && x12 && x11 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && x21 && ~x68 && ~x10 && x12 && ~x11 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s170;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && x21 && ~x68 && ~x10 && ~x12 && x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && x21 && ~x68 && ~x10 && ~x12 && ~x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && x9 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s171;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && x10 && x18 && x19 && x11 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && x10 && x18 && x19 && ~x11 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s168;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && x10 && x18 && ~x19 && x12 && x16 && x11 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && x10 && x18 && ~x19 && x12 && x16 && ~x11 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s168;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && x10 && x18 && ~x19 && x12 && ~x16 && x11 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s168;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && x10 && x18 && ~x19 && x12 && ~x16 && ~x11 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && x10 && x18 && ~x19 && ~x12 && x11 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && x10 && x18 && ~x19 && ~x12 && ~x11 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s168;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && x10 && ~x18 && x11 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s168;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && x10 && ~x18 && ~x11 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && ~x10 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && x3 )
						begin
							y8 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s172;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && ~x3 && x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y9 = 1'b1;	
							nx_state = s173;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && ~x3 && x11 && ~x2 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && ~x3 && ~x11 && x9 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && ~x3 && ~x11 && ~x9 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && x68 && x11 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && x68 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && x20 && x13 && x9 && x11 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && x20 && x13 && x9 && ~x11 && x2 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && x20 && x13 && x9 && ~x11 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && x20 && x13 && ~x9 && x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s174;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && x20 && x13 && ~x9 && ~x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && x20 && ~x13 && x2 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && x20 && ~x13 && ~x2 && x9 && x11 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && x20 && ~x13 && ~x2 && x9 && ~x11 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && x20 && ~x13 && ~x2 && ~x9 && x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s174;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && x20 && ~x13 && ~x2 && ~x9 && ~x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && ~x20 && x2 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && ~x20 && ~x2 && x9 && x11 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && ~x20 && ~x2 && x9 && ~x11 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && ~x20 && ~x2 && ~x9 && x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s174;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && ~x20 && ~x2 && ~x9 && ~x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && ~x19 && x2 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && ~x19 && ~x2 && x9 && x11 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && ~x19 && ~x2 && x9 && ~x11 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && ~x19 && ~x2 && ~x9 && x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s174;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && ~x19 && ~x2 && ~x9 && ~x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && ~x1 && x68 && x22 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && ~x1 && x68 && ~x22 && x21 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && ~x1 && x68 && ~x22 && ~x21 && x11 && x3 && x6 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s175;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && ~x1 && x68 && ~x22 && ~x21 && x11 && x3 && ~x6 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && ~x1 && x68 && ~x22 && ~x21 && x11 && ~x3 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && ~x1 && x68 && ~x22 && ~x21 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x66 && ~x65 && ~x1 && ~x68 )
						nx_state = s1;
					else if( ~x69 && x70 && x63 && x62 && x11 && x10 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s176;
						end
					else if( ~x69 && x70 && x63 && x62 && x11 && ~x10 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s177;
						end
					else if( ~x69 && x70 && x63 && x62 && ~x11 && x10 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x69 && x70 && x63 && x62 && ~x11 && ~x10 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x69 && x70 && x63 && x62 && ~x11 && ~x10 && ~x1 && x2 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x69 && x70 && x63 && x62 && ~x11 && ~x10 && ~x1 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && x11 && x43 && x13 && x32 && x3 && x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s99;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && x11 && x43 && x13 && x32 && x3 && ~x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && x11 && x43 && x13 && x32 && ~x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && x11 && x43 && x13 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && x11 && x43 && ~x13 && x5 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s181;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && x11 && x43 && ~x13 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && x11 && ~x43 && x44 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && x11 && ~x43 && ~x44 && x14 && x7 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && x11 && ~x43 && ~x44 && x14 && ~x7 && x1 && x5 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s183;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && x11 && ~x43 && ~x44 && x14 && ~x7 && x1 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && x11 && ~x43 && ~x44 && x14 && ~x7 && ~x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && x11 && ~x43 && ~x44 && ~x14 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && ~x11 && x12 && x8 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && ~x11 && x12 && ~x8 && x5 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s183;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && ~x11 && x12 && ~x8 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && ~x11 && ~x12 && x13 && x45 && x32 && x36 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && ~x11 && ~x12 && x13 && x45 && x32 && ~x36 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && ~x11 && ~x12 && x13 && x45 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && ~x11 && ~x12 && x13 && ~x45 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && ~x11 && ~x12 && ~x13 && x1 && x14 && x5 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s183;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && ~x11 && ~x12 && ~x13 && x1 && x14 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && ~x11 && ~x12 && ~x13 && x1 && ~x14 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && x64 && ~x11 && ~x12 && ~x13 && ~x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && ~x64 && x15 && x12 && x23 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && ~x64 && x15 && x12 && ~x23 && x4 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && ~x64 && x15 && x12 && ~x23 && ~x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && ~x64 && x15 && ~x12 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && ~x64 && ~x15 && x39 && x46 && x48 && x36 )
						nx_state = s1;
					else if( ~x69 && x70 && x63 && ~x62 && x10 && ~x64 && ~x15 && x39 && x46 && x48 && ~x36 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && ~x64 && ~x15 && x39 && x46 && ~x48 && x36 )
						nx_state = s1;
					else if( ~x69 && x70 && x63 && ~x62 && x10 && ~x64 && ~x15 && x39 && x46 && ~x48 && ~x36 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && ~x64 && ~x15 && x39 && ~x46 && x36 )
						nx_state = s1;
					else if( ~x69 && x70 && x63 && ~x62 && x10 && ~x64 && ~x15 && x39 && ~x46 && ~x36 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && x63 && ~x62 && x10 && ~x64 && ~x15 && ~x39 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && x64 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && x15 && x1 && x22 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s190;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && x15 && x1 && ~x22 && x2 && x11 && x5 && x3 )
						nx_state = s1;
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && x15 && x1 && ~x22 && x2 && x11 && x5 && ~x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && x15 && x1 && ~x22 && x2 && x11 && ~x5 && x3 )
						nx_state = s1;
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && x15 && x1 && ~x22 && x2 && x11 && ~x5 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && x15 && x1 && ~x22 && x2 && ~x11 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && x15 && x1 && ~x22 && x2 && ~x11 && ~x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && x15 && x1 && ~x22 && ~x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && x15 && ~x1 && x11 && x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && x15 && ~x1 && x11 && ~x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && x15 && ~x1 && ~x11 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && ~x15 && x11 && x34 && x8 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && ~x15 && x11 && x34 && ~x8 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && ~x15 && x11 && x34 && ~x8 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && ~x15 && x11 && ~x34 && x32 && x7 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && ~x15 && x11 && ~x34 && x32 && ~x7 && x43 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && ~x15 && x11 && ~x34 && x32 && ~x7 && x43 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && ~x15 && x11 && ~x34 && x32 && ~x7 && ~x43 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && ~x15 && x11 && ~x34 && ~x32 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && ~x15 && ~x11 && x12 && x20 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && ~x15 && ~x11 && x12 && ~x20 && x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && ~x15 && ~x11 && x12 && ~x20 && ~x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && ~x15 && ~x11 && ~x12 && x13 && x1 && x3 && x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && ~x15 && ~x11 && ~x12 && x13 && x1 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && ~x15 && ~x11 && ~x12 && x13 && x1 && ~x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && ~x15 && ~x11 && ~x12 && x13 && ~x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && x63 && ~x62 && ~x10 && ~x64 && ~x15 && ~x11 && ~x12 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && x70 && ~x63 && x64 && x15 && x16 && x62 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s193;
						end
					else if( ~x69 && x70 && ~x63 && x64 && x15 && x16 && x62 && ~x5 && x6 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s194;
						end
					else if( ~x69 && x70 && ~x63 && x64 && x15 && x16 && x62 && ~x5 && ~x6 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s195;
						end
					else if( ~x69 && x70 && ~x63 && x64 && x15 && x16 && ~x62 && x5 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x70 && ~x63 && x64 && x15 && x16 && ~x62 && ~x5 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x69 && x70 && ~x63 && x64 && x15 && x16 && ~x62 && ~x5 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x69 && x70 && ~x63 && x64 && x15 && ~x16 && x62 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( ~x69 && x70 && ~x63 && x64 && x15 && ~x16 && x62 && ~x1 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x63 && x64 && x15 && ~x16 && ~x62 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x63 && x64 && x15 && ~x16 && ~x62 && ~x1 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x63 && x64 && ~x15 && x16 && x62 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( ~x69 && x70 && ~x63 && x64 && ~x15 && x16 && ~x62 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x63 && x64 && ~x15 && ~x16 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x69 && x70 && ~x63 && x64 && ~x15 && ~x16 && ~x1 && x62 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( ~x69 && x70 && ~x63 && x64 && ~x15 && ~x16 && ~x1 && ~x62 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && x10 && x39 && x44 && x41 && x36 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && x10 && x39 && x44 && x41 && ~x36 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && x10 && x39 && x44 && ~x41 && x36 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && x10 && x39 && x44 && ~x41 && ~x36 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && x10 && x39 && ~x44 && x36 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && x10 && x39 && ~x44 && ~x36 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && x10 && ~x39 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s201;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && ~x10 && x11 && x34 && x8 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && ~x10 && x11 && x34 && ~x8 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && ~x10 && x11 && x34 && ~x8 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && ~x10 && x11 && ~x34 && x32 && x7 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && ~x10 && x11 && ~x34 && x32 && ~x7 && x26 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && ~x10 && x11 && ~x34 && x32 && ~x7 && x26 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && ~x10 && x11 && ~x34 && x32 && ~x7 && ~x26 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && ~x10 && x11 && ~x34 && ~x32 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && ~x10 && ~x11 && x12 && x20 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && ~x10 && ~x11 && x12 && ~x20 && x2 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && ~x10 && ~x11 && x12 && ~x20 && ~x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && ~x10 && ~x11 && ~x12 && x13 && x1 && x3 && x6 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && ~x10 && ~x11 && ~x12 && x13 && x1 && x3 && ~x6 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && ~x10 && ~x11 && ~x12 && x13 && x1 && ~x3 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && ~x10 && ~x11 && ~x12 && x13 && ~x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && x14 && ~x10 && ~x11 && ~x12 && ~x13 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && ~x14 && x10 && x11 && x1 && x2 && x4 && x5 && x3 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && ~x14 && x10 && x11 && x1 && x2 && x4 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && ~x14 && x10 && x11 && x1 && x2 && x4 && ~x5 && x3 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && ~x14 && x10 && x11 && x1 && x2 && x4 && ~x5 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && ~x14 && x10 && x11 && x1 && x2 && ~x4 && x3 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && ~x14 && x10 && x11 && x1 && x2 && ~x4 && ~x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && ~x14 && x10 && x11 && x1 && ~x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && ~x14 && x10 && x11 && ~x1 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && ~x14 && x10 && ~x11 && x12 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && ~x14 && x10 && ~x11 && ~x12 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && ~x14 && ~x10 && x11 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && ~x14 && ~x10 && x11 && ~x1 && x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && ~x14 && ~x10 && x11 && ~x1 && ~x2 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && ~x14 && ~x10 && ~x11 && x12 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && ~x14 && ~x10 && ~x11 && x12 && ~x1 && x4 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && ~x14 && ~x10 && ~x11 && x12 && ~x1 && ~x4 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && ~x14 && ~x10 && ~x11 && ~x12 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s206;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && ~x14 && ~x10 && ~x11 && ~x12 && ~x1 && x2 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && ~x14 && ~x10 && ~x11 && ~x12 && ~x1 && ~x2 && x9 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && x62 && ~x14 && ~x10 && ~x11 && ~x12 && ~x1 && ~x2 && ~x9 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && x17 && x18 && x40 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s45;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && x17 && x18 && ~x40 && x2 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && x17 && x18 && ~x40 && ~x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && x17 && ~x18 && x19 && x1 && x10 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && x17 && ~x18 && x19 && x1 && ~x10 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && x17 && ~x18 && x19 && ~x1 && x6 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s45;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && x17 && ~x18 && x19 && ~x1 && ~x6 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && x17 && ~x18 && ~x19 && x1 && x39 && x4 && x5 && x3 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && x17 && ~x18 && ~x19 && x1 && x39 && x4 && x5 && ~x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && x17 && ~x18 && ~x19 && x1 && x39 && x4 && ~x5 && x3 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && x17 && ~x18 && ~x19 && x1 && x39 && x4 && ~x5 && ~x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && x17 && ~x18 && ~x19 && x1 && x39 && ~x4 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && x17 && ~x18 && ~x19 && x1 && x39 && ~x4 && ~x3 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && x17 && ~x18 && ~x19 && x1 && ~x39 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s45;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && x17 && ~x18 && ~x19 && ~x1 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && ~x17 && x18 && x40 && x19 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && ~x17 && x18 && x40 && ~x19 && x39 && x4 && x5 && x3 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && ~x17 && x18 && x40 && ~x19 && x39 && x4 && x5 && ~x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && ~x17 && x18 && x40 && ~x19 && x39 && x4 && ~x5 && x3 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && ~x17 && x18 && x40 && ~x19 && x39 && x4 && ~x5 && ~x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && ~x17 && x18 && x40 && ~x19 && x39 && ~x4 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && ~x17 && x18 && x40 && ~x19 && x39 && ~x4 && ~x3 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && ~x17 && x18 && x40 && ~x19 && ~x39 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s45;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && ~x17 && x18 && ~x40 && x19 && x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && ~x17 && x18 && ~x40 && x19 && ~x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && ~x17 && x18 && ~x40 && ~x19 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x70 && ~x63 && ~x64 && ~x62 && ~x17 && ~x18 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s45;
						end
					else if( ~x69 && ~x70 && x46 && x44 && x10 && x45 && x39 && x36 && x35 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && x46 && x44 && x10 && x45 && x39 && x36 && ~x35 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x46 && x44 && x10 && x45 && x39 && ~x36 && x43 && x42 && x40 )
						begin
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x69 && ~x70 && x46 && x44 && x10 && x45 && x39 && ~x36 && x43 && x42 && ~x40 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x69 && ~x70 && x46 && x44 && x10 && x45 && x39 && ~x36 && x43 && ~x42 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x46 && x44 && x10 && x45 && x39 && ~x36 && ~x43 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x69 && ~x70 && x46 && x44 && x10 && x45 && ~x39 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x69 && ~x70 && x46 && x44 && x10 && ~x45 && x3 && x7 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x69 && ~x70 && x46 && x44 && x10 && ~x45 && x3 && ~x7 && x1 && x5 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x70 && x46 && x44 && x10 && ~x45 && x3 && ~x7 && x1 && ~x5 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s209;
						end
					else if( ~x69 && ~x70 && x46 && x44 && x10 && ~x45 && x3 && ~x7 && ~x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && x46 && x44 && x10 && ~x45 && ~x3 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && x46 && x44 && ~x10 && x45 && x11 && x34 && x8 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && ~x70 && x46 && x44 && ~x10 && x45 && x11 && x34 && ~x8 && x5 )
						begin
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x69 && ~x70 && x46 && x44 && ~x10 && x45 && x11 && x34 && ~x8 && ~x5 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x46 && x44 && ~x10 && x45 && x11 && ~x34 && x32 && x7 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && ~x70 && x46 && x44 && ~x10 && x45 && x11 && ~x34 && x32 && ~x7 && x22 && x5 )
						begin
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x69 && ~x70 && x46 && x44 && ~x10 && x45 && x11 && ~x34 && x32 && ~x7 && x22 && ~x5 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x46 && x44 && ~x10 && x45 && x11 && ~x34 && x32 && ~x7 && ~x22 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x69 && ~x70 && x46 && x44 && ~x10 && x45 && x11 && ~x34 && ~x32 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x69 && ~x70 && x46 && x44 && ~x10 && x45 && ~x11 && x12 && x20 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x69 && ~x70 && x46 && x44 && ~x10 && x45 && ~x11 && x12 && ~x20 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && x46 && x44 && ~x10 && x45 && ~x11 && x12 && ~x20 && ~x2 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x70 && x46 && x44 && ~x10 && x45 && ~x11 && ~x12 && x13 && x1 && x3 && x6 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && ~x70 && x46 && x44 && ~x10 && x45 && ~x11 && ~x12 && x13 && x1 && x3 && ~x6 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x46 && x44 && ~x10 && x45 && ~x11 && ~x12 && x13 && x1 && ~x3 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x46 && x44 && ~x10 && x45 && ~x11 && ~x12 && x13 && ~x1 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x69 && ~x70 && x46 && x44 && ~x10 && x45 && ~x11 && ~x12 && ~x13 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x69 && ~x70 && x46 && x44 && ~x10 && ~x45 && x3 && x1 && x5 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x70 && x46 && x44 && ~x10 && ~x45 && x3 && x1 && ~x5 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s209;
						end
					else if( ~x69 && ~x70 && x46 && x44 && ~x10 && ~x45 && x3 && ~x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && x46 && x44 && ~x10 && ~x45 && ~x3 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && x47 && x7 && x45 && x9 && x5 && x3 && x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && x47 && x7 && x45 && x9 && x5 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && x47 && x7 && x45 && x9 && x5 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && x47 && x7 && x45 && x9 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && x47 && x7 && x45 && ~x9 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && x47 && x7 && ~x45 && x8 && x1 && x3 && x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && x47 && x7 && ~x45 && x8 && x1 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && x47 && x7 && ~x45 && x8 && x1 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && x47 && x7 && ~x45 && x8 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && x47 && x7 && ~x45 && ~x8 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && x47 && ~x7 && x1 && x45 && x15 && x5 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	
							nx_state = s213;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && x47 && ~x7 && x1 && x45 && x15 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && x47 && ~x7 && x1 && x45 && ~x15 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && x47 && ~x7 && x1 && ~x45 && x8 && x5 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	
							nx_state = s213;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && x47 && ~x7 && x1 && ~x45 && x8 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && x47 && ~x7 && x1 && ~x45 && ~x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && x47 && ~x7 && ~x1 && x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && x47 && ~x7 && ~x1 && ~x8 && x2 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && x47 && ~x7 && ~x1 && ~x8 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && x11 && x12 && x10 && x5 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && x11 && x12 && x10 && ~x5 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && x11 && x12 && ~x10 && x8 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && x11 && x12 && ~x10 && ~x8 && x5 )
						begin
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && x11 && x12 && ~x10 && ~x8 && ~x5 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && x11 && ~x12 && x10 && x1 && x5 && x13 )
						begin
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && x11 && ~x12 && x10 && x1 && x5 && ~x13 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && x11 && ~x12 && x10 && x1 && ~x5 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && x11 && ~x12 && x10 && ~x1 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && x11 && ~x12 && ~x10 && x13 && x7 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && x11 && ~x12 && ~x10 && x13 && ~x7 && x1 && x5 )
						begin
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && x11 && ~x12 && ~x10 && x13 && ~x7 && x1 && ~x5 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && x11 && ~x12 && ~x10 && x13 && ~x7 && ~x1 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && x11 && ~x12 && ~x10 && ~x13 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && ~x11 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && ~x11 && ~x10 && x12 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && ~x11 && ~x10 && x12 && ~x1 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && ~x11 && ~x10 && x12 && ~x1 && ~x2 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && ~x11 && ~x10 && ~x12 && x13 && x1 && x3 && x6 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && ~x11 && ~x10 && ~x12 && x13 && x1 && x3 && ~x6 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && ~x11 && ~x10 && ~x12 && x13 && x1 && ~x3 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && ~x11 && ~x10 && ~x12 && x13 && ~x1 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && x45 && ~x11 && ~x10 && ~x12 && ~x13 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && ~x45 && x9 && x11 && x1 && x5 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && ~x45 && x9 && x11 && x1 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && ~x45 && x9 && x11 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && ~x45 && x9 && ~x11 && x7 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && ~x45 && x9 && ~x11 && ~x7 && x1 && x5 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && ~x45 && x9 && ~x11 && ~x7 && x1 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && ~x45 && x9 && ~x11 && ~x7 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && ~x45 && ~x9 && x10 && x11 && x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && ~x45 && ~x9 && x10 && x11 && ~x8 && x5 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && ~x45 && ~x9 && x10 && x11 && ~x8 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && ~x45 && ~x9 && x10 && ~x11 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							nx_state = s214;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && ~x45 && ~x9 && x10 && ~x11 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && ~x45 && ~x9 && ~x10 && x1 && x11 && x3 && x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && ~x45 && ~x9 && ~x10 && x1 && x11 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && ~x45 && ~x9 && ~x10 && x1 && x11 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && ~x45 && ~x9 && ~x10 && x1 && ~x11 && x5 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s176;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && ~x45 && ~x9 && ~x10 && x1 && ~x11 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x46 && ~x44 && ~x47 && ~x45 && ~x9 && ~x10 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && x44 && x10 && x11 && x1 && x2 && x4 && x5 && x3 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x46 && x45 && x44 && x10 && x11 && x1 && x2 && x4 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && x44 && x10 && x11 && x1 && x2 && x4 && ~x5 && x3 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x46 && x45 && x44 && x10 && x11 && x1 && x2 && x4 && ~x5 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && x44 && x10 && x11 && x1 && x2 && ~x4 && x3 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && x44 && x10 && x11 && x1 && x2 && ~x4 && ~x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && x44 && x10 && x11 && x1 && ~x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && x44 && x10 && x11 && ~x1 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && x44 && x10 && ~x11 && x12 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && x44 && x10 && ~x11 && ~x12 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s215;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && x44 && ~x10 && x11 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && x44 && ~x10 && x11 && ~x1 && x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && x44 && ~x10 && x11 && ~x1 && ~x2 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && x44 && ~x10 && ~x11 && x12 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && x44 && ~x10 && ~x11 && x12 && ~x1 && x4 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && x44 && ~x10 && ~x11 && x12 && ~x1 && ~x4 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && x44 && ~x10 && ~x11 && ~x12 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s216;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && x44 && ~x10 && ~x11 && ~x12 && ~x1 && x2 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && x44 && ~x10 && ~x11 && ~x12 && ~x1 && ~x2 && x9 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && x44 && ~x10 && ~x11 && ~x12 && ~x1 && ~x2 && ~x9 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && x47 && x10 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && x47 && x10 && ~x1 && x4 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && x47 && x10 && ~x1 && ~x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && x47 && ~x10 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && x47 && ~x10 && ~x1 && x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && x47 && ~x10 && ~x1 && ~x2 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && x12 && x11 && x10 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && x12 && x11 && ~x10 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s177;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && x12 && ~x11 && x10 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s176;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && x12 && ~x11 && ~x10 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && x12 && ~x11 && ~x10 && ~x1 && x2 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && x12 && ~x11 && ~x10 && ~x1 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && ~x12 && x9 && x11 && x1 && x5 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && ~x12 && x9 && x11 && x1 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && ~x12 && x9 && x11 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && ~x12 && x9 && ~x11 && x7 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && ~x12 && x9 && ~x11 && ~x7 && x1 && x5 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && ~x12 && x9 && ~x11 && ~x7 && x1 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && ~x12 && x9 && ~x11 && ~x7 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && ~x12 && ~x9 && x10 && x11 && x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && ~x12 && ~x9 && x10 && x11 && ~x8 && x5 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && ~x12 && ~x9 && x10 && x11 && ~x8 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && ~x12 && ~x9 && x10 && ~x11 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							nx_state = s214;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && ~x12 && ~x9 && x10 && ~x11 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && ~x12 && ~x9 && ~x10 && x1 && x11 && x3 && x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && ~x12 && ~x9 && ~x10 && x1 && x11 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && ~x12 && ~x9 && ~x10 && x1 && x11 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && ~x12 && ~x9 && ~x10 && x1 && ~x11 && x5 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s176;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && ~x12 && ~x9 && ~x10 && x1 && ~x11 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x46 && x45 && ~x44 && ~x47 && ~x12 && ~x9 && ~x10 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && x47 && x10 && x12 && x23 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && x47 && x10 && x12 && ~x23 && x4 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && x47 && x10 && x12 && ~x23 && ~x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && x47 && x10 && ~x12 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && x47 && ~x10 && x1 && x22 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s190;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && x47 && ~x10 && x1 && ~x22 && x2 && x11 && x5 && x3 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && x47 && ~x10 && x1 && ~x22 && x2 && x11 && x5 && ~x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && x47 && ~x10 && x1 && ~x22 && x2 && x11 && ~x5 && x3 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && x47 && ~x10 && x1 && ~x22 && x2 && x11 && ~x5 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && x47 && ~x10 && x1 && ~x22 && x2 && ~x11 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && x47 && ~x10 && x1 && ~x22 && x2 && ~x11 && ~x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && x47 && ~x10 && x1 && ~x22 && ~x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && x47 && ~x10 && ~x1 && x11 && x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && x47 && ~x10 && ~x1 && x11 && ~x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && x47 && ~x10 && ~x1 && ~x11 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && ~x47 && x9 && x16 && x8 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && ~x47 && x9 && x16 && ~x8 && x5 )
						begin
							y7 = 1'b1;	
							nx_state = s82;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && ~x47 && x9 && x16 && ~x8 && ~x5 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && ~x47 && x9 && ~x16 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && ~x47 && ~x9 && x10 && x5 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && ~x47 && ~x9 && x10 && ~x5 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && ~x47 && ~x9 && ~x10 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && ~x47 && ~x9 && ~x10 && ~x1 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && x44 && ~x47 && ~x9 && ~x10 && ~x1 && ~x2 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && x11 && x12 && x10 && x13 && x7 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && x11 && x12 && x10 && x13 && ~x7 && x1 && x5 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && x11 && x12 && x10 && x13 && ~x7 && x1 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && x11 && x12 && x10 && x13 && ~x7 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && x11 && x12 && x10 && ~x13 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							nx_state = s214;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && x11 && x12 && x10 && ~x13 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && x11 && x12 && ~x10 && x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && x11 && x12 && ~x10 && ~x8 && x5 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && x11 && x12 && ~x10 && ~x8 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && x11 && ~x12 && x10 && x1 && x5 && x13 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && x11 && ~x12 && x10 && x1 && x5 && ~x13 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s176;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && x11 && ~x12 && x10 && x1 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && x11 && ~x12 && x10 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && x11 && ~x12 && ~x10 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s177;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && ~x11 && x10 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && ~x11 && ~x10 && x12 && x1 && x3 && x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && ~x11 && ~x10 && x12 && x1 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && ~x11 && ~x10 && x12 && x1 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && ~x11 && ~x10 && x12 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && ~x11 && ~x10 && ~x12 && x13 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && ~x11 && ~x10 && ~x12 && x13 && ~x1 && x2 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && ~x11 && ~x10 && ~x12 && x13 && ~x1 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && ~x46 && ~x45 && ~x44 && ~x11 && ~x10 && ~x12 && ~x13 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s176;
						end
					else nx_state = s1;
				s2 : if( x64 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s218;
						end
					else if( ~x64 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x64 && ~x3 && x1 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s46;
						end
					else if( ~x64 && ~x3 && x1 && ~x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x64 && ~x3 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else nx_state = s2;
				s3 : if( x70 && x62 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							y8 = 1'b1;	
							nx_state = s219;
						end
					else if( x70 && ~x62 && x64 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	
							nx_state = s220;
						end
					else if( x70 && ~x62 && ~x64 && x65 && x66 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( x70 && ~x62 && ~x64 && x65 && ~x66 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x70 && ~x62 && ~x64 && ~x65 )
						begin
							y3 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s223;
						end
					else if( ~x70 && x66 && x21 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && x66 && ~x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s224;
						end
					else if( ~x70 && ~x66 && x68 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && ~x66 && ~x68 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s225;
						end
					else nx_state = s3;
				s4 : if( 1'b1 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else nx_state = s4;
				s5 : if( x70 && x62 && x64 )
						begin
							y22 = 1'b1;	
							nx_state = s130;
						end
					else if( x70 && x62 && ~x64 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x70 && x62 && ~x64 && ~x7 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x70 && ~x62 && x63 )
						begin
							y6 = 1'b1;	y17 = 1'b1;	y34 = 1'b1;	
							nx_state = s226;
						end
					else if( x70 && ~x62 && ~x63 && x21 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x70 && ~x62 && ~x63 && ~x21 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else if( ~x70 && x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x22 && x23 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x22 && ~x23 && x18 && x14 )
						nx_state = s47;
					else if( ~x70 && ~x21 && x22 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s47;
					else if( ~x70 && ~x21 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x70 && ~x21 && ~x22 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x70 && ~x21 && ~x22 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 && x23 && ~x19 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else nx_state = s5;
				s6 : if( x70 && x62 && x66 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x70 && x62 && ~x66 && x3 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s230;
						end
					else if( x70 && x62 && ~x66 && x3 && ~x2 )
						nx_state = s6;
					else if( x70 && x62 && ~x66 && ~x3 && x4 && x2 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	
							nx_state = s231;
						end
					else if( x70 && x62 && ~x66 && ~x3 && x4 && ~x2 )
						nx_state = s6;
					else if( x70 && x62 && ~x66 && ~x3 && ~x4 && x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x70 && x62 && ~x66 && ~x3 && ~x4 && ~x2 )
						nx_state = s6;
					else if( x70 && ~x62 && x64 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s232;
						end
					else if( x70 && ~x62 && ~x64 && x15 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && ~x64 && ~x15 && x3 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s230;
						end
					else if( x70 && ~x62 && ~x64 && ~x15 && x3 && ~x2 )
						nx_state = s6;
					else if( x70 && ~x62 && ~x64 && ~x15 && ~x3 && x4 && x2 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	
							nx_state = s231;
						end
					else if( x70 && ~x62 && ~x64 && ~x15 && ~x3 && x4 && ~x2 )
						nx_state = s6;
					else if( x70 && ~x62 && ~x64 && ~x15 && ~x3 && ~x4 && x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x70 && ~x62 && ~x64 && ~x15 && ~x3 && ~x4 && ~x2 )
						nx_state = s6;
					else if( ~x70 && x66 && x16 && x21 && x7 && x10 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x70 && x66 && x16 && x21 && x7 && ~x10 )
						begin
							y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s233;
						end
					else if( ~x70 && x66 && x16 && x21 && ~x7 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x70 && x66 && x16 && ~x21 && x7 && x10 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x70 && x66 && x16 && ~x21 && x7 && ~x10 )
						begin
							y4 = 1'b1;	y18 = 1'b1;	
							nx_state = s234;
						end
					else if( ~x70 && x66 && x16 && ~x21 && ~x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x70 && x66 && ~x16 && x17 && x9 && x21 && x10 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x70 && x66 && ~x16 && x17 && x9 && x21 && ~x10 && x13 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x70 && x66 && ~x16 && x17 && x9 && x21 && ~x10 && ~x13 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x66 && ~x16 && x17 && x9 && x21 && ~x10 && ~x13 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x66 && ~x16 && x17 && x9 && x21 && ~x10 && ~x13 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && x17 && x9 && x21 && ~x10 && ~x13 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && x17 && x9 && ~x21 && x10 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x70 && x66 && ~x16 && x17 && x9 && ~x21 && ~x10 && x13 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x70 && x66 && ~x16 && x17 && x9 && ~x21 && ~x10 && ~x13 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x70 && x66 && ~x16 && x17 && x9 && ~x21 && ~x10 && ~x13 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x70 && x66 && ~x16 && x17 && x9 && ~x21 && ~x10 && ~x13 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && x17 && x9 && ~x21 && ~x10 && ~x13 && ~x20 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && x17 && ~x9 && x21 && x10 && x11 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x70 && x66 && ~x16 && x17 && ~x9 && x21 && x10 && ~x11 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x66 && ~x16 && x17 && ~x9 && x21 && x10 && ~x11 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x66 && ~x16 && x17 && ~x9 && x21 && x10 && ~x11 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && x17 && ~x9 && x21 && x10 && ~x11 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && x17 && ~x9 && x21 && ~x10 && x12 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x70 && x66 && ~x16 && x17 && ~x9 && x21 && ~x10 && ~x12 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x66 && ~x16 && x17 && ~x9 && x21 && ~x10 && ~x12 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x66 && ~x16 && x17 && ~x9 && x21 && ~x10 && ~x12 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && x17 && ~x9 && x21 && ~x10 && ~x12 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && x17 && ~x9 && ~x21 && x10 && x11 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x70 && x66 && ~x16 && x17 && ~x9 && ~x21 && x10 && ~x11 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x70 && x66 && ~x16 && x17 && ~x9 && ~x21 && x10 && ~x11 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x70 && x66 && ~x16 && x17 && ~x9 && ~x21 && x10 && ~x11 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && x17 && ~x9 && ~x21 && x10 && ~x11 && ~x20 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && x17 && ~x9 && ~x21 && ~x10 && x12 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x70 && x66 && ~x16 && x17 && ~x9 && ~x21 && ~x10 && ~x12 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x70 && x66 && ~x16 && x17 && ~x9 && ~x21 && ~x10 && ~x12 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x70 && x66 && ~x16 && x17 && ~x9 && ~x21 && ~x10 && ~x12 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && x17 && ~x9 && ~x21 && ~x10 && ~x12 && ~x20 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && ~x17 && x7 )
						begin
							y4 = 1'b1;	y17 = 1'b1;	
							nx_state = s235;
						end
					else if( ~x70 && x66 && ~x16 && ~x17 && ~x7 && x21 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x70 && x66 && ~x16 && ~x17 && ~x7 && ~x21 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x70 && ~x66 && x21 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && ~x66 && x21 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && ~x66 && x21 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x70 && ~x66 && x21 && ~x3 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x21 && x22 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x70 && ~x66 && ~x21 && x22 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x70 && ~x66 && ~x21 && x22 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x21 && x22 && ~x6 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x21 && ~x22 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x70 && ~x66 && ~x21 && ~x22 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x70 && ~x66 && ~x21 && ~x22 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x21 && ~x22 && ~x8 )
						nx_state = s1;
					else nx_state = s6;
				s7 : if( x62 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x62 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s238;
						end
					else if( ~x62 && ~x13 )
						begin
							y6 = 1'b1;	
							nx_state = s239;
						end
					else nx_state = s7;
				s8 : if( x70 && x25 && x9 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x70 && x25 && ~x9 )
						begin
							y13 = 1'b1;	
							nx_state = s240;
						end
					else if( x70 && ~x25 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x70 && x65 && x66 && x67 && x23 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && x67 && ~x23 && x6 && x15 && x8 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && x66 && x67 && ~x23 && x6 && x15 && ~x8 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && x65 && x66 && x67 && ~x23 && x6 && ~x15 && x16 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && x66 && x67 && ~x23 && x6 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( ~x70 && x65 && x66 && x67 && ~x23 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && x66 && ~x67 && x60 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && x61 && x62 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && x61 && ~x62 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && x16 && x12 && x7 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && x16 && x12 && ~x7 && x14 && x11 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && x16 && x12 && ~x7 && x14 && ~x11 )
						begin
							y15 = 1'b1;	
							nx_state = s243;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && x16 && x12 && ~x7 && ~x14 )
						nx_state = s47;
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && x16 && ~x12 && x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && x16 && ~x12 && ~x7 && x13 && x11 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && x16 && ~x12 && ~x7 && x13 && ~x11 )
						begin
							y15 = 1'b1;	
							nx_state = s243;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && x16 && ~x12 && ~x7 && ~x13 )
						nx_state = s47;
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && ~x16 && x11 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s244;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && ~x16 && x11 && ~x7 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s245;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && ~x16 && x11 && ~x7 && ~x12 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && ~x16 && ~x11 && x6 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && ~x16 && ~x11 && ~x6 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && ~x16 && ~x11 && ~x6 && ~x2 && x12 && x7 )
						begin
							y11 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && ~x16 && ~x11 && ~x6 && ~x2 && x12 && ~x7 )
						begin
							y11 = 1'b1;	
							nx_state = s248;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && ~x16 && ~x11 && ~x6 && ~x2 && ~x12 && x7 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && ~x16 && ~x11 && ~x6 && ~x2 && ~x12 && ~x7 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && x6 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && x7 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && x7 && ~x2 && x12 )
						begin
							y11 = 1'b1;	
							nx_state = s250;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && x7 && ~x2 && ~x12 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && x12 && x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && x12 && x11 && ~x2 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s251;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && x12 && ~x11 && x9 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && x12 && ~x11 && x9 && ~x2 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s251;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && x12 && ~x11 && ~x9 )
						nx_state = s47;
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && ~x12 && x11 && x10 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && ~x12 && x11 && x10 && ~x2 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s251;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && ~x12 && x11 && ~x10 )
						nx_state = s47;
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && ~x12 && ~x11 && x8 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && ~x12 && ~x11 && x8 && ~x2 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s251;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && ~x12 && ~x11 && ~x8 )
						nx_state = s47;
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && ~x16 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && ~x16 && ~x2 && x7 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && ~x16 && ~x2 && ~x7 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s139;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 && ~x62 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && x16 && x13 && x18 && x15 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && x16 && x13 && x18 && ~x15 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && x16 && x13 && ~x18 && x14 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && x16 && x13 && ~x18 && ~x14 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && x16 && ~x13 && x14 && x18 && x15 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && x16 && ~x13 && x14 && x18 && ~x15 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s253;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && x16 && ~x13 && x14 && ~x18 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s253;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && x16 && ~x13 && ~x14 && x18 && x15 && x6 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && x16 && ~x13 && ~x14 && x18 && x15 && ~x6 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && x16 && ~x13 && ~x14 && x18 && x15 && ~x6 && x4 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x21 && x17 && x16 && ~x13 && ~x14 && x18 && x15 && ~x6 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x21 && x17 && x16 && ~x13 && ~x14 && x18 && ~x15 && x5 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && x16 && ~x13 && ~x14 && x18 && ~x15 && ~x5 && x4 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && x16 && ~x13 && ~x14 && x18 && ~x15 && ~x5 && x4 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x21 && x17 && x16 && ~x13 && ~x14 && x18 && ~x15 && ~x5 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x21 && x17 && x16 && ~x13 && ~x14 && ~x18 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && x13 && x18 && x15 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && x13 && x18 && ~x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && x13 && x18 && ~x15 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && x13 && ~x18 && x14 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && x13 && ~x18 && x14 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && x13 && ~x18 && x14 && ~x2 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && x13 && ~x18 && ~x14 && x12 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && x13 && ~x18 && ~x14 && x12 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && x13 && ~x18 && ~x14 && x12 && ~x2 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && x13 && ~x18 && ~x14 && ~x12 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && x13 && ~x18 && ~x14 && ~x12 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && x13 && ~x18 && ~x14 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && x13 && ~x18 && ~x14 && ~x12 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && x18 && x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && x18 && x15 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && x18 && ~x15 && x12 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && x18 && ~x15 && x12 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && x18 && ~x15 && ~x12 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && x18 && ~x15 && ~x12 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && x18 && ~x15 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && x18 && ~x15 && ~x12 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && ~x18 && x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && ~x18 && x11 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && ~x18 && x11 && ~x2 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && ~x18 && ~x11 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && ~x18 && ~x11 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && ~x18 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && ~x18 && ~x11 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && x15 && x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && x15 && x11 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && x15 && ~x11 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && x15 && ~x11 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && x15 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && x15 && ~x11 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && ~x15 && x10 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && ~x15 && x10 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && ~x15 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && ~x15 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && ~x15 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && ~x15 && ~x10 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && ~x18 && x10 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && ~x18 && x10 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && ~x18 && x10 && ~x2 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && ~x18 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && ~x18 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && ~x18 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && ~x18 && ~x10 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x21 && ~x17 && x16 && x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x65 && ~x66 && x21 && ~x17 && x16 && x14 && ~x13 && x15 && x18 && x12 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && x65 && ~x66 && x21 && ~x17 && x16 && x14 && ~x13 && x15 && x18 && ~x12 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s256;
						end
					else if( ~x70 && x65 && ~x66 && x21 && ~x17 && x16 && x14 && ~x13 && x15 && ~x18 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && x65 && ~x66 && x21 && ~x17 && x16 && x14 && ~x13 && ~x15 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s258;
						end
					else if( ~x70 && x65 && ~x66 && x21 && ~x17 && x16 && ~x14 && x15 && x18 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && x65 && ~x66 && x21 && ~x17 && x16 && ~x14 && x15 && x18 && ~x13 )
						begin
							y24 = 1'b1;	
							nx_state = s259;
						end
					else if( ~x70 && x65 && ~x66 && x21 && ~x17 && x16 && ~x14 && x15 && ~x18 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s259;
						end
					else if( ~x70 && x65 && ~x66 && x21 && ~x17 && x16 && ~x14 && x15 && ~x18 && ~x13 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s256;
						end
					else if( ~x70 && x65 && ~x66 && x21 && ~x17 && x16 && ~x14 && ~x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && x21 && ~x17 && x16 && ~x14 && ~x15 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && x21 && ~x17 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && x13 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && x21 && ~x17 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( ~x70 && x65 && ~x66 && x21 && ~x17 && ~x16 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && x21 && ~x17 && ~x16 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && x21 && ~x17 && ~x16 && ~x2 && ~x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s35;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && x10 && x15 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s253;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && x10 && ~x15 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && ~x10 && x15 && x6 && x14 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s261;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && ~x10 && x15 && x6 && ~x14 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && ~x10 && x15 && ~x6 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && ~x10 && x15 && ~x6 && x4 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && ~x10 && x15 && ~x6 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && ~x10 && ~x15 && x5 && x14 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && ~x10 && ~x15 && x5 && ~x14 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && ~x10 && ~x15 && ~x5 && x4 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && ~x10 && ~x15 && ~x5 && x4 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && ~x10 && ~x15 && ~x5 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && x13 && x15 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && x13 && ~x15 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s261;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && ~x13 && x15 && x6 && x14 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && ~x13 && x15 && x6 && ~x14 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && ~x13 && x15 && ~x6 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && ~x13 && x15 && ~x6 && x4 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && ~x13 && x15 && ~x6 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && ~x13 && ~x15 && x5 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && ~x13 && ~x15 && x5 && ~x14 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && ~x13 && ~x15 && ~x5 && x4 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && ~x13 && ~x15 && ~x5 && x4 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && ~x13 && ~x15 && ~x5 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && x13 && x15 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && x13 && ~x15 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s253;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && x14 && x19 && x15 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && x14 && x19 && ~x15 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s261;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && x14 && ~x19 && x15 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s261;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && x14 && ~x19 && ~x15 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && ~x14 && x15 && x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && ~x14 && x15 && ~x6 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && ~x14 && x15 && ~x6 && x4 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && ~x14 && x15 && ~x6 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && ~x14 && ~x15 && x5 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && ~x14 && ~x15 && ~x5 && x4 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && ~x14 && ~x15 && ~x5 && x4 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && ~x14 && ~x15 && ~x5 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && x19 && x10 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && x19 && ~x10 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && x19 && ~x10 && ~x2 && x14 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && x19 && ~x10 && ~x2 && x14 && ~x3 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && x19 && ~x10 && ~x2 && ~x14 && x12 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && x19 && ~x10 && ~x2 && ~x14 && x12 && ~x3 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && x19 && ~x10 && ~x2 && ~x14 && ~x12 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && x19 && ~x10 && ~x2 && ~x14 && ~x12 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && x19 && ~x10 && ~x2 && ~x14 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && x19 && ~x10 && ~x2 && ~x14 && ~x12 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && ~x19 && x13 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s253;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && ~x19 && ~x13 && x14 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && ~x19 && ~x13 && x14 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && ~x19 && ~x13 && x14 && ~x2 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && ~x19 && ~x13 && ~x14 && x11 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && ~x19 && ~x13 && ~x14 && ~x11 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && ~x19 && ~x13 && ~x14 && ~x11 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && ~x19 && ~x13 && ~x14 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && ~x19 && ~x13 && ~x14 && ~x11 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && x10 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && x14 && x13 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && x14 && x13 && ~x3 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && x14 && ~x13 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && x14 && ~x13 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && x14 && ~x13 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && x14 && ~x13 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && ~x14 && x11 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && ~x14 && x11 && ~x3 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && ~x14 && ~x11 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && ~x14 && ~x11 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && ~x14 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && ~x14 && ~x11 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && x13 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && x13 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && ~x13 && x14 && x12 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && ~x13 && x14 && ~x12 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && ~x13 && x14 && ~x12 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && ~x13 && x14 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && ~x13 && x14 && ~x12 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && ~x13 && ~x14 && x10 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && ~x13 && ~x14 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && ~x13 && ~x14 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && ~x13 && ~x14 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && ~x13 && ~x14 && ~x10 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && x13 && x15 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && x13 && ~x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && x13 && ~x15 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && x14 && x15 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && x14 && x15 && ~x3 && x19 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && x14 && x15 && ~x3 && ~x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && x14 && ~x15 && x12 && x19 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && x14 && ~x15 && x12 && x19 && ~x3 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && x14 && ~x15 && x12 && ~x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && x14 && ~x15 && ~x12 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && x14 && ~x15 && ~x12 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && x14 && ~x15 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && x14 && ~x15 && ~x12 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && x15 && x11 && x19 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && x15 && x11 && x19 && ~x3 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && x15 && x11 && ~x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && x15 && ~x11 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && x15 && ~x11 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && x15 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && x15 && ~x11 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && ~x15 && x10 && x19 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && ~x15 && x10 && x19 && ~x3 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && ~x15 && x10 && ~x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && ~x15 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && ~x15 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && ~x15 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && ~x15 && ~x10 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && x13 && x15 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && x13 && ~x15 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s253;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && ~x13 && x15 && x6 && x14 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && ~x13 && x15 && x6 && ~x14 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && ~x13 && x15 && ~x6 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && ~x13 && x15 && ~x6 && x4 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && ~x13 && x15 && ~x6 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && ~x13 && ~x15 && x5 && x14 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s261;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && ~x13 && ~x15 && x5 && ~x14 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && ~x13 && ~x15 && ~x5 && x4 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && ~x13 && ~x15 && ~x5 && x4 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && ~x13 && ~x15 && ~x5 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && ~x18 && x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && ~x18 && x14 && ~x13 && x15 && x16 )
						begin
							y26 = 1'b1;	
							nx_state = s262;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && ~x18 && x14 && ~x13 && x15 && ~x16 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && ~x18 && x14 && ~x13 && ~x15 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && ~x18 && ~x14 && x15 && x13 )
						begin
							y26 = 1'b1;	
							nx_state = s262;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && ~x18 && ~x14 && x15 && ~x13 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && ~x18 && ~x14 && ~x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && ~x18 && ~x14 && ~x15 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && ~x18 && ~x14 && ~x15 && ~x2 && ~x3 && x13 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	
							nx_state = s263;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && ~x18 && ~x14 && ~x15 && ~x2 && ~x3 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && x13 && x20 && x14 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && x13 && x20 && ~x14 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && x13 && ~x20 && x15 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && x13 && ~x20 && ~x15 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && x14 && x20 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s253;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && x14 && ~x20 && x15 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && x14 && ~x20 && ~x15 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s253;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && ~x14 && x20 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && ~x14 && ~x20 && x15 && x6 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && ~x14 && ~x20 && x15 && ~x6 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && ~x14 && ~x20 && x15 && ~x6 && x4 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && ~x14 && ~x20 && x15 && ~x6 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && ~x14 && ~x20 && ~x15 && x5 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && ~x14 && ~x20 && ~x15 && ~x5 && x4 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && ~x14 && ~x20 && ~x15 && ~x5 && x4 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && ~x14 && ~x20 && ~x15 && ~x5 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && x20 && x14 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && x20 && x14 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && x20 && x14 && ~x2 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && x20 && ~x14 && x12 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && x20 && ~x14 && x12 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && x20 && ~x14 && x12 && ~x2 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && x20 && ~x14 && ~x12 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && x20 && ~x14 && ~x12 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && x20 && ~x14 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && x20 && ~x14 && ~x12 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && ~x20 && x15 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && ~x20 && ~x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && ~x20 && ~x15 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && x20 && x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && x20 && x11 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && x20 && x11 && ~x2 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && x20 && ~x11 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && x20 && ~x11 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && x20 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && x20 && ~x11 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && ~x20 && x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && ~x20 && x15 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && ~x20 && ~x15 && x12 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && ~x20 && ~x15 && x12 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && ~x20 && ~x15 && ~x12 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && ~x20 && ~x15 && ~x12 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && ~x20 && ~x15 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && ~x20 && ~x15 && ~x12 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && x20 && x10 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && x20 && x10 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && x20 && x10 && ~x2 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && x20 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && x20 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && x20 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && x20 && ~x10 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && x15 && x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && x15 && x11 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && x15 && ~x11 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && x15 && ~x11 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && x15 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && x15 && ~x11 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && ~x15 && x10 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && ~x15 && x10 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && ~x15 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && ~x15 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && ~x15 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && ~x15 && ~x10 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && x18 && x19 && x10 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && x18 && x19 && ~x10 && x15 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && x18 && x19 && ~x10 && ~x15 )
						begin
							y26 = 1'b1;	
							nx_state = s262;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && x18 && ~x19 && x13 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && x18 && ~x19 && ~x13 && x15 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	
							nx_state = s263;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && x18 && ~x19 && ~x13 && ~x15 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && ~x18 && x19 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && ~x18 && x19 && ~x13 && x15 )
						begin
							y26 = 1'b1;	
							nx_state = s262;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && ~x18 && x19 && ~x13 && ~x15 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && ~x18 && ~x19 && x13 )
						begin
							y26 = 1'b1;	
							nx_state = s262;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && ~x18 && ~x19 && ~x13 && x15 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && ~x18 && ~x19 && ~x13 && ~x15 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && x15 && x19 && x18 && x10 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	
							nx_state = s263;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && x15 && x19 && x18 && ~x10 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && x15 && x19 && ~x18 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && x15 && x19 && ~x18 && ~x13 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && x15 && ~x19 && x13 )
						nx_state = s47;
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && x15 && ~x19 && ~x13 && x18 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && x15 && ~x19 && ~x13 && x18 && ~x3 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && x15 && ~x19 && ~x13 && ~x18 && x3 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	
							nx_state = s263;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && x15 && ~x19 && ~x13 && ~x18 && ~x3 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && x2 && x18 && x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && x2 && x18 && ~x19 && x13 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && x2 && x18 && ~x19 && ~x13 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s264;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && x2 && ~x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && x19 && x18 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && x19 && x18 && ~x10 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && x19 && ~x18 && x13 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	
							nx_state = s263;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && x19 && ~x18 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && ~x19 && x13 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && ~x19 && ~x13 && x18 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && ~x19 && ~x13 && ~x18 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s264;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && ~x16 && x18 && x19 && x10 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && ~x16 && x18 && x19 && ~x10 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && ~x16 && x18 && x19 && ~x10 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && ~x16 && x18 && x19 && ~x10 && ~x2 && ~x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s35;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && ~x16 && x18 && ~x19 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && ~x16 && x18 && ~x19 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && ~x16 && x18 && ~x19 && ~x2 && ~x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s35;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && ~x16 && ~x18 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && ~x16 && ~x18 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && x22 && ~x16 && ~x18 && ~x2 && ~x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s35;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && x15 && x13 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && x15 && ~x13 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && x15 && ~x13 && ~x2 && x14 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && x15 && ~x13 && ~x2 && x14 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && x15 && ~x13 && ~x2 && ~x14 && x11 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && x15 && ~x13 && ~x2 && ~x14 && x11 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && x15 && ~x13 && ~x2 && ~x14 && ~x11 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && x15 && ~x13 && ~x2 && ~x14 && ~x11 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && x15 && ~x13 && ~x2 && ~x14 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && x15 && ~x13 && ~x2 && ~x14 && ~x11 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && x13 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && x14 && x12 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && x14 && x12 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && x14 && ~x12 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && x14 && ~x12 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && x14 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && x14 && ~x12 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && ~x14 && x10 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && ~x14 && x10 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && ~x14 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && ~x14 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && ~x14 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && ~x14 && ~x10 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && ~x18 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && ~x18 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && ~x18 && ~x2 && ~x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s35;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && x14 && ~x13 && x15 && x20 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && x14 && ~x13 && x15 && ~x20 && x12 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && x14 && ~x13 && x15 && ~x20 && ~x12 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && x14 && ~x13 && ~x15 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s264;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && ~x14 && x15 && x20 && x13 )
						begin
							y26 = 1'b1;	
							nx_state = s262;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && ~x14 && x15 && x20 && ~x13 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && ~x14 && x15 && ~x20 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && ~x14 && x15 && ~x20 && ~x13 )
						begin
							y26 = 1'b1;	
							nx_state = s262;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && ~x14 && ~x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && ~x14 && ~x15 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && x13 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && ~x16 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && ~x16 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && ~x16 && ~x2 && ~x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s35;
						end
					else if( ~x70 && ~x65 && x21 && x68 && x16 && x17 && x10 && x15 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && ~x65 && x21 && x68 && x16 && x17 && x10 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x70 && ~x65 && x21 && x68 && x16 && x17 && ~x10 && x15 && x7 && x14 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s253;
						end
					else if( ~x70 && ~x65 && x21 && x68 && x16 && x17 && ~x10 && x15 && x7 && ~x14 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x70 && ~x65 && x21 && x68 && x16 && x17 && ~x10 && x15 && ~x7 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x65 && x21 && x68 && x16 && x17 && ~x10 && x15 && ~x7 && x9 && ~x8 && x14 )
						nx_state = s8;
					else if( ~x70 && ~x65 && x21 && x68 && x16 && x17 && ~x10 && x15 && ~x7 && x9 && ~x8 && ~x14 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x21 && x68 && x16 && x17 && ~x10 && x15 && ~x7 && ~x9 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x21 && x68 && x16 && x17 && ~x10 && ~x15 && x8 && x14 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s267;
						end
					else if( ~x70 && ~x65 && x21 && x68 && x16 && x17 && ~x10 && ~x15 && x8 && ~x14 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x70 && ~x65 && x21 && x68 && x16 && x17 && ~x10 && ~x15 && ~x8 && x9 && x14 )
						nx_state = s8;
					else if( ~x70 && ~x65 && x21 && x68 && x16 && x17 && ~x10 && ~x15 && ~x8 && x9 && ~x14 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x65 && x21 && x68 && x16 && x17 && ~x10 && ~x15 && ~x8 && x9 && ~x14 && ~x7 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x21 && x68 && x16 && x17 && ~x10 && ~x15 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x21 && x68 && x16 && ~x17 && x14 && x10 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x65 && x21 && x68 && x16 && ~x17 && x14 && ~x10 && x15 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x70 && ~x65 && x21 && x68 && x16 && ~x17 && x14 && ~x10 && x15 && ~x13 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( ~x70 && ~x65 && x21 && x68 && x16 && ~x17 && x14 && ~x10 && ~x15 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	
							nx_state = s268;
						end
					else if( ~x70 && ~x65 && x21 && x68 && x16 && ~x17 && ~x14 && x2 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s269;
						end
					else if( ~x70 && ~x65 && x21 && x68 && x16 && ~x17 && ~x14 && ~x2 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && x21 && x68 && x16 && ~x17 && ~x14 && ~x2 && ~x4 && x15 && x10 )
						begin
							y11 = 1'b1;	
							nx_state = s248;
						end
					else if( ~x70 && ~x65 && x21 && x68 && x16 && ~x17 && ~x14 && ~x2 && ~x4 && x15 && ~x10 )
						begin
							y11 = 1'b1;	
							nx_state = s250;
						end
					else if( ~x70 && ~x65 && x21 && x68 && x16 && ~x17 && ~x14 && ~x2 && ~x4 && ~x15 && x10 )
						begin
							y2 = 1'b1;	y16 = 1'b1;	y24 = 1'b1;	
							nx_state = s270;
						end
					else if( ~x70 && ~x65 && x21 && x68 && x16 && ~x17 && ~x14 && ~x2 && ~x4 && ~x15 && ~x10 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && x2 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s269;
						end
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && x10 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && x10 && ~x4 )
						begin
							y11 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && x15 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && x15 && ~x4 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && x13 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && x13 && ~x4 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && ~x13 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && ~x13 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && ~x13 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && ~x13 && ~x9 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && x12 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && x12 && ~x4 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && ~x12 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && ~x12 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && ~x12 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && ~x12 && ~x9 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && x11 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && x11 && ~x4 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && ~x11 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && ~x11 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && ~x11 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && ~x11 && ~x9 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && ~x17 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && ~x17 && ~x4 && x10 )
						begin
							y11 = 1'b1;	
							nx_state = s272;
						end
					else if( ~x70 && ~x65 && x21 && x68 && ~x16 && ~x2 && ~x17 && ~x4 && ~x10 )
						begin
							y11 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x70 && ~x65 && x21 && ~x68 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( ~x70 && ~x65 && ~x21 && x22 && x68 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x70 && ~x65 && ~x21 && x22 && x68 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x70 && ~x65 && ~x21 && x22 && x68 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && x22 && x68 && ~x7 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && x22 && ~x68 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x70 && ~x65 && ~x21 && x22 && ~x68 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x70 && ~x65 && ~x21 && x22 && ~x68 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && x22 && ~x68 && x23 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && x22 && ~x68 && ~x23 && x18 && x14 )
						nx_state = s47;
					else if( ~x70 && ~x65 && ~x21 && x22 && ~x68 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s47;
					else if( ~x70 && ~x65 && ~x21 && x22 && ~x68 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && x22 && ~x68 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && ~x22 && x68 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x65 && ~x21 && ~x22 && ~x68 && x23 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s274;
						end
					else if( ~x70 && ~x65 && ~x21 && ~x22 && ~x68 && ~x23 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s275;
						end
					else nx_state = s8;
				s9 : if( x65 && x70 && x62 && x66 && x2 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s6;
						end
					else if( x65 && x70 && x62 && x66 && x2 && ~x4 && x5 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x70 && x62 && x66 && x2 && ~x4 && ~x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x65 && x70 && x62 && x66 && ~x2 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x65 && x70 && x62 && x66 && ~x2 && ~x3 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x65 && x70 && x62 && ~x66 && x5 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	
							nx_state = s276;
						end
					else if( x65 && x70 && x62 && ~x66 && ~x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s6;
						end
					else if( x65 && x70 && ~x62 && x63 && x15 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s6;
						end
					else if( x65 && x70 && ~x62 && x63 && ~x15 && x5 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	
							nx_state = s276;
						end
					else if( x65 && x70 && ~x62 && x63 && ~x15 && ~x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s6;
						end
					else if( x65 && x70 && ~x62 && ~x63 )
						begin
							y39 = 1'b1;	
							nx_state = s277;
						end
					else if( x65 && ~x70 && x16 && x11 && x12 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s278;
						end
					else if( x65 && ~x70 && x16 && x11 && ~x12 && x13 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s278;
						end
					else if( x65 && ~x70 && x16 && x11 && ~x12 && ~x13 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( x65 && ~x70 && x16 && ~x11 && x13 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s135;
						end
					else if( x65 && ~x70 && x16 && ~x11 && ~x13 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x65 && ~x70 && ~x16 && x17 && x11 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x65 && ~x70 && ~x16 && x17 && x11 && ~x13 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x65 && ~x70 && ~x16 && x17 && ~x11 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x65 && ~x70 && ~x16 && ~x17 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x65 && x70 && x62 && x18 && x17 && x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	
							nx_state = s20;
						end
					else if( ~x65 && x70 && x62 && x18 && x17 && ~x1 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && x70 && x62 && x18 && x17 && ~x1 && ~x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x65 && x70 && x62 && x18 && ~x17 && x19 && x5 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x65 && x70 && x62 && x18 && ~x17 && x19 && ~x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && x70 && x62 && x18 && ~x17 && ~x19 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x65 && x70 && x62 && ~x18 && x17 && x7 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s215;
						end
					else if( ~x65 && x70 && x62 && ~x18 && x17 && ~x7 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s280;
						end
					else if( ~x65 && x70 && x62 && ~x18 && ~x17 && x19 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	
							nx_state = s20;
						end
					else if( ~x65 && x70 && x62 && ~x18 && ~x17 && ~x19 && x5 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x65 && x70 && x62 && ~x18 && ~x17 && ~x19 && x5 && ~x3 && x4 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( ~x65 && x70 && x62 && ~x18 && ~x17 && ~x19 && x5 && ~x3 && ~x4 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && x70 && x62 && ~x18 && ~x17 && ~x19 && ~x5 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x65 && x70 && ~x62 && x63 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s238;
						end
					else if( ~x65 && x70 && ~x62 && x63 && ~x13 )
						begin
							y6 = 1'b1;	
							nx_state = s239;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && x19 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && x19 && ~x3 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && x19 && ~x3 && ~x4 && x5 && x12 )
						begin
							y54 = 1'b1;	
							nx_state = s281;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && x19 && ~x3 && ~x4 && x5 && ~x12 )
						begin
							y55 = 1'b1;	
							nx_state = s282;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && x19 && ~x3 && ~x4 && ~x5 && x6 && x12 && x11 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && x19 && ~x3 && ~x4 && ~x5 && x6 && x12 && ~x11 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && x19 && ~x3 && ~x4 && ~x5 && x6 && x12 && ~x11 && x9 && ~x10 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && x19 && ~x3 && ~x4 && ~x5 && x6 && x12 && ~x11 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && x19 && ~x3 && ~x4 && ~x5 && x6 && ~x12 && x10 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && x19 && ~x3 && ~x4 && ~x5 && x6 && ~x12 && ~x10 && x9 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && x19 && ~x3 && ~x4 && ~x5 && x6 && ~x12 && ~x10 && x9 && ~x11 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && x19 && ~x3 && ~x4 && ~x5 && x6 && ~x12 && ~x10 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && x19 && ~x3 && ~x4 && ~x5 && ~x6 && x12 )
						begin
							y58 = 1'b1;	y59 = 1'b1;	
							nx_state = s284;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && x19 && ~x3 && ~x4 && ~x5 && ~x6 && ~x12 )
						begin
							y56 = 1'b1;	y57 = 1'b1;	
							nx_state = s284;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && x17 )
						begin
							y53 = 1'b1;	
							nx_state = s285;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && x6 && x12 && x5 )
						begin
							y45 = 1'b1;	
							nx_state = s286;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && x6 && x12 && ~x5 && x14 )
						begin
							y47 = 1'b1;	
							nx_state = s287;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && x6 && x12 && ~x5 && ~x14 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && x6 && x12 && ~x5 && ~x14 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && x6 && x12 && ~x5 && ~x14 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && x6 && x12 && ~x5 && ~x14 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && x6 && ~x12 && x5 )
						begin
							y5 = 1'b1;	
							nx_state = s64;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && x6 && ~x12 && ~x5 && x13 )
						begin
							y47 = 1'b1;	
							nx_state = s287;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && x6 && ~x12 && ~x5 && ~x13 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && x6 && ~x12 && ~x5 && ~x13 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && x6 && ~x12 && ~x5 && ~x13 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && x6 && ~x12 && ~x5 && ~x13 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && ~x6 && x5 && x12 && x16 )
						begin
							y47 = 1'b1;	
							nx_state = s287;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && ~x6 && x5 && x12 && ~x16 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && ~x6 && x5 && x12 && ~x16 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && ~x6 && x5 && x12 && ~x16 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && ~x6 && x5 && x12 && ~x16 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && ~x6 && x5 && ~x12 && x15 )
						begin
							y47 = 1'b1;	
							nx_state = s287;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && ~x6 && x5 && ~x12 && ~x15 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && ~x6 && x5 && ~x12 && ~x15 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && ~x6 && x5 && ~x12 && ~x15 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && ~x6 && x5 && ~x12 && ~x15 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x18 && ~x19 && ~x17 && ~x3 && ~x4 && ~x6 && ~x5 )
						begin
							y47 = 1'b1;	
							nx_state = s287;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && ~x18 && x5 && x19 && x12 && x6 )
						begin
							y26 = 1'b1;	
							nx_state = s262;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && ~x18 && x5 && x19 && x12 && ~x6 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && ~x18 && x5 && x19 && ~x12 && x6 )
						begin
							y25 = 1'b1;	
							nx_state = s238;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && ~x18 && x5 && x19 && ~x12 && ~x6 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && ~x18 && x5 && x19 && ~x12 && ~x6 && ~x3 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && ~x18 && x5 && x19 && ~x12 && ~x6 && ~x3 && ~x4 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y29 = 1'b1;	
							nx_state = s288;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && ~x18 && x5 && ~x19 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && ~x18 && x5 && ~x19 && ~x3 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && ~x18 && x5 && ~x19 && ~x3 && ~x4 && x6 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && ~x18 && x5 && ~x19 && ~x3 && ~x4 && ~x6 )
						begin
							y17 = 1'b1;	
							nx_state = s98;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && ~x18 && ~x5 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && ~x18 && ~x5 && ~x3 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && ~x18 && ~x5 && ~x3 && ~x4 && x19 && x12 && x6 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && ~x18 && ~x5 && ~x3 && ~x4 && x19 && x12 && ~x6 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && ~x18 && ~x5 && ~x3 && ~x4 && x19 && ~x12 && x6 )
						begin
							y30 = 1'b1;	
							nx_state = s291;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && ~x18 && ~x5 && ~x3 && ~x4 && x19 && ~x12 && ~x6 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && ~x18 && ~x5 && ~x3 && ~x4 && ~x19 )
						begin
							y16 = 1'b1;	
							nx_state = s293;
						end
					else if( ~x65 && ~x70 && x66 && x62 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && x63 && x64 && x17 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && x63 && x64 && x17 && ~x13 && x12 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && x63 && x64 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x66 && ~x62 && x63 && x64 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x66 && ~x62 && x63 && ~x64 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s294;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && x64 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s295;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && x14 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && x14 && ~x8 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && ~x14 && x7 && x8 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s296;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && ~x14 && x7 && ~x8 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s297;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && ~x14 && ~x7 && x8 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && x19 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && x19 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && ~x14 && ~x7 && ~x8 && x13 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && x19 && x12 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && x19 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && x7 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && x7 && ~x3 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && x7 && ~x3 && ~x4 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && ~x7 && x9 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && ~x7 && x9 && ~x3 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && ~x7 && x9 && ~x3 && ~x4 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && ~x7 && ~x9 && x3 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && ~x7 && ~x9 && ~x3 && x19 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && ~x7 && ~x9 && ~x3 && x19 && ~x13 && x12 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && ~x7 && ~x9 && ~x3 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && ~x7 && ~x9 && ~x3 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && x7 && x11 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && x7 && x11 && ~x3 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && x7 && x11 && ~x3 && ~x4 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && x7 && ~x11 && x3 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && x7 && ~x11 && ~x3 && x19 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && x7 && ~x11 && ~x3 && x19 && ~x13 && x12 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && x7 && ~x11 && ~x3 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && x7 && ~x11 && ~x3 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && ~x7 && x10 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && ~x7 && x10 && ~x3 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && ~x7 && x10 && ~x3 && ~x4 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && x3 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x3 && x19 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x3 && x19 && ~x13 && x12 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x3 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x3 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && ~x16 && x15 && x7 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s298;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && ~x16 && x15 && ~x7 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && ~x16 && x15 && ~x7 && ~x3 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && ~x16 && x15 && ~x7 && ~x3 && ~x4 && x8 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && ~x16 && x15 && ~x7 && ~x3 && ~x4 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && ~x16 && ~x15 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && ~x16 && ~x15 && ~x3 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && ~x16 && ~x15 && ~x3 && ~x4 && x14 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y28 = 1'b1;	
							nx_state = s299;
						end
					else if( ~x65 && ~x70 && x66 && ~x62 && ~x63 && ~x64 && ~x16 && ~x15 && ~x3 && ~x4 && ~x14 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s294;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && x26 && x17 && x11 && x13 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s300;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && x26 && x17 && x11 && ~x13 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && x26 && x17 && ~x11 && x12 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && x26 && x17 && ~x11 && x12 && ~x13 )
						begin
							y14 = 1'b1;	
							nx_state = s124;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && x26 && x17 && ~x11 && ~x12 && x13 && x14 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s301;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && x26 && x17 && ~x11 && ~x12 && x13 && ~x14 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && x26 && x17 && ~x11 && ~x12 && x13 && ~x14 && x18 && ~x15 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && x26 && x17 && ~x11 && ~x12 && x13 && ~x14 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && x26 && x17 && ~x11 && ~x12 && ~x13 && x15 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s301;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && x26 && x17 && ~x11 && ~x12 && ~x13 && ~x15 && x18 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && x26 && x17 && ~x11 && ~x12 && ~x13 && ~x15 && x18 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && x26 && x17 && ~x11 && ~x12 && ~x13 && ~x15 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && x26 && ~x17 && x13 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && x26 && ~x17 && ~x13 && x12 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && x26 && ~x17 && ~x13 && ~x12 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && x26 && ~x17 && ~x13 && ~x12 && ~x2 && x11 && x4 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s126;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && x26 && ~x17 && ~x13 && ~x12 && ~x2 && x11 && ~x4 )
						begin
							y8 = 1'b1;	y17 = 1'b1;	y23 = 1'b1;	
							nx_state = s303;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && x26 && ~x17 && ~x13 && ~x12 && ~x2 && ~x11 && x4 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && x26 && ~x17 && ~x13 && ~x12 && ~x2 && ~x11 && ~x4 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s304;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && x11 && x13 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && x11 && ~x13 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && ~x11 && x12 && x13 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && ~x11 && x12 && ~x13 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && ~x11 && ~x12 && x13 && x14 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s306;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && ~x11 && ~x12 && x13 && ~x14 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && ~x11 && ~x12 && x13 && ~x14 && x20 && ~x15 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && ~x11 && ~x12 && x13 && ~x14 && ~x20 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && ~x11 && ~x12 && ~x13 && x15 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s306;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && ~x11 && ~x12 && ~x13 && ~x15 && x20 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && ~x11 && ~x12 && ~x13 && ~x15 && x20 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && ~x11 && ~x12 && ~x13 && ~x15 && ~x20 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && x11 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && x11 && ~x3 && x12 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && x11 && ~x3 && x12 && ~x4 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s256;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && x11 && ~x3 && ~x12 && x13 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && x11 && ~x3 && ~x12 && x13 && ~x4 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s308;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && x11 && ~x3 && ~x12 && ~x13 && x4 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s304;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && x11 && ~x3 && ~x12 && ~x13 && ~x4 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && ~x11 && x13 && x12 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s35;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && ~x11 && x13 && ~x12 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s308;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && ~x11 && ~x13 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && ~x11 && ~x13 && ~x12 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && ~x11 && ~x13 && ~x12 && ~x3 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && ~x11 && ~x13 && ~x12 && ~x3 && ~x4 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s309;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && x11 && x9 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && x11 && x9 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && x11 && x9 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && x11 && x9 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && x11 && ~x9 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && x11 && ~x9 && ~x2 && x4 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && x11 && ~x9 && ~x2 && ~x4 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s304;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && ~x11 && x12 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && ~x11 && x12 && ~x2 && x4 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && ~x11 && x12 && ~x2 && ~x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && ~x11 && ~x12 && x8 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && ~x11 && ~x12 && x8 && ~x2 && x4 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && ~x11 && ~x12 && x8 && ~x2 && ~x4 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s304;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && ~x11 && ~x12 && ~x8 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && ~x11 && ~x12 && ~x8 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && ~x11 && ~x12 && ~x8 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && ~x11 && ~x12 && ~x8 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && x11 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && x11 && ~x2 && x4 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && x11 && ~x2 && ~x4 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && x12 && x10 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && x12 && x10 && ~x2 && x4 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && x12 && x10 && ~x2 && ~x4 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s304;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && x12 && ~x10 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && x12 && ~x10 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && x12 && ~x10 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && x12 && ~x10 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && ~x12 && x9 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && ~x12 && x9 && ~x2 && x4 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && ~x12 && x9 && ~x2 && ~x4 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s304;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && ~x12 && ~x9 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && ~x12 && ~x9 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && ~x12 && ~x9 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && ~x12 && ~x9 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && ~x17 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && ~x17 && ~x2 && x4 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && x26 && ~x17 && ~x2 && ~x4 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && x11 && x9 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && x11 && x9 && ~x4 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && x11 && ~x9 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && x11 && ~x9 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && x11 && ~x9 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && x11 && ~x9 && ~x20 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && ~x11 && x12 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && ~x11 && x12 && ~x4 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && ~x11 && ~x12 && x7 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && ~x11 && ~x12 && x7 && ~x4 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && ~x11 && ~x12 && ~x7 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && ~x11 && ~x12 && ~x7 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && ~x11 && ~x12 && ~x7 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && ~x11 && ~x12 && ~x7 && ~x20 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && x11 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s311;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && x11 && ~x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && x12 && x10 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && x12 && x10 && ~x4 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && x12 && ~x10 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && x12 && ~x10 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && x12 && ~x10 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && x12 && ~x10 && ~x20 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && x8 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && x8 && ~x4 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && ~x8 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && ~x8 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && ~x8 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && ~x8 && ~x20 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && ~x17 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && ~x17 && ~x4 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s258;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && ~x24 && x25 && x26 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && ~x24 && x25 && ~x26 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && ~x24 && x25 && ~x26 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && ~x24 && x25 && ~x26 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && ~x24 && x25 && ~x26 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x26 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x26 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x26 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x26 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && ~x67 && x68 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && x21 && x10 && x11 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && x21 && x10 && ~x11 )
						nx_state = s9;
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && x21 && ~x10 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s170;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s313;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && x19 && x15 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y17 = 1'b1;	
							nx_state = s314;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && x19 && ~x15 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							nx_state = s315;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && x15 && x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s316;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && x15 && ~x14 && x16 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s316;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && x15 && ~x14 && ~x16 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && x15 && ~x14 && ~x16 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && x15 && ~x14 && ~x16 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && x15 && ~x14 && ~x16 && ~x5 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && ~x15 && x14 && x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s316;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && ~x15 && x14 && ~x18 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && ~x15 && x14 && ~x18 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && ~x15 && x14 && ~x18 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && ~x15 && x14 && ~x18 && ~x5 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && ~x15 && ~x14 && x17 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s316;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && ~x5 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && ~x20 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && ~x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && ~x22 && x10 && x19 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && ~x22 && x10 && x19 && ~x15 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	
							nx_state = s315;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && ~x22 && x10 && ~x19 && x20 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && ~x22 && x10 && ~x19 && ~x20 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( ~x65 && ~x70 && ~x66 && ~x67 && ~x68 && ~x21 && ~x22 && ~x10 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s170;
						end
					else nx_state = s9;
				s10 : if( x69 && x65 && x66 && x2 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s6;
						end
					else if( x69 && x65 && x66 && x2 && ~x4 && x5 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	
							nx_state = s7;
						end
					else if( x69 && x65 && x66 && x2 && ~x4 && ~x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && x65 && x66 && ~x2 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x65 && x66 && ~x2 && ~x3 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x69 && x65 && ~x66 && x6 && x4 && x5 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s18;
						end
					else if( x69 && x65 && ~x66 && x6 && x4 && x5 && ~x1 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( x69 && x65 && ~x66 && x6 && x4 && ~x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x65 && ~x66 && x6 && ~x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( x69 && x65 && ~x66 && ~x6 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x65 && x66 && x4 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( x69 && ~x65 && x66 && x4 && ~x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x65 && x66 && ~x4 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x65 && ~x66 && x18 && x17 && x4 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s320;
						end
					else if( x69 && ~x65 && ~x66 && x18 && x17 && ~x4 && x1 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x65 && ~x66 && x18 && x17 && ~x4 && x1 && ~x3 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x65 && ~x66 && x18 && x17 && ~x4 && ~x1 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x65 && ~x66 && x18 && ~x17 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x65 && ~x66 && ~x18 && x17 && x11 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x69 && ~x65 && ~x66 && ~x18 && x17 && ~x11 && x16 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x65 && ~x66 && ~x18 && x17 && ~x11 && ~x16 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x66 && ~x18 && ~x17 && x19 && x1 && x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x65 && ~x66 && ~x18 && ~x17 && x19 && x1 && ~x2 && x3 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x65 && ~x66 && ~x18 && ~x17 && x19 && x1 && ~x2 && ~x3 )
						nx_state = s10;
					else if( x69 && ~x65 && ~x66 && ~x18 && ~x17 && x19 && ~x1 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && ~x65 && ~x66 && ~x18 && ~x17 && ~x19 && x2 && x1 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && ~x65 && ~x66 && ~x18 && ~x17 && ~x19 && x2 && x1 && ~x3 && x4 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x65 && ~x66 && ~x18 && ~x17 && ~x19 && x2 && x1 && ~x3 && ~x4 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x65 && ~x66 && ~x18 && ~x17 && ~x19 && x2 && ~x1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x65 && ~x66 && ~x18 && ~x17 && ~x19 && ~x2 && x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	
							nx_state = s20;
						end
					else if( x69 && ~x65 && ~x66 && ~x18 && ~x17 && ~x19 && ~x2 && ~x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && x70 && x62 && x64 && x10 && x61 && x39 && x46 && x51 && x36 )
						nx_state = s10;
					else if( ~x69 && x70 && x62 && x64 && x10 && x61 && x39 && x46 && x51 && ~x36 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x69 && x70 && x62 && x64 && x10 && x61 && x39 && x46 && ~x51 && x36 )
						nx_state = s10;
					else if( ~x69 && x70 && x62 && x64 && x10 && x61 && x39 && x46 && ~x51 && ~x36 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && x70 && x62 && x64 && x10 && x61 && x39 && ~x46 && x36 )
						nx_state = s10;
					else if( ~x69 && x70 && x62 && x64 && x10 && x61 && x39 && ~x46 && ~x36 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && x70 && x62 && x64 && x10 && x61 && ~x39 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s201;
						end
					else if( ~x69 && x70 && x62 && x64 && x10 && ~x61 && x11 && x1 && x2 && x4 && x5 && x3 )
						nx_state = s10;
					else if( ~x69 && x70 && x62 && x64 && x10 && ~x61 && x11 && x1 && x2 && x4 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && x70 && x62 && x64 && x10 && ~x61 && x11 && x1 && x2 && x4 && ~x5 && x3 )
						nx_state = s10;
					else if( ~x69 && x70 && x62 && x64 && x10 && ~x61 && x11 && x1 && x2 && x4 && ~x5 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && x70 && x62 && x64 && x10 && ~x61 && x11 && x1 && x2 && ~x4 && x3 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && x62 && x64 && x10 && ~x61 && x11 && x1 && x2 && ~x4 && ~x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && x62 && x64 && x10 && ~x61 && x11 && x1 && ~x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && x70 && x62 && x64 && x10 && ~x61 && x11 && ~x1 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x70 && x62 && x64 && x10 && ~x61 && ~x11 && x12 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && x70 && x62 && x64 && x10 && ~x61 && ~x11 && ~x12 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && x11 && x61 && x34 && x8 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && x11 && x61 && x34 && ~x8 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && x11 && x61 && x34 && ~x8 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && x11 && x61 && ~x34 && x32 && x7 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && x11 && x61 && ~x34 && x32 && ~x7 && x54 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && x11 && x61 && ~x34 && x32 && ~x7 && x54 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && x11 && x61 && ~x34 && x32 && ~x7 && ~x54 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && x11 && x61 && ~x34 && ~x32 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && x11 && ~x61 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && x11 && ~x61 && ~x1 && x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && x11 && ~x61 && ~x1 && ~x2 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && ~x11 && x12 && x61 && x20 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && ~x11 && x12 && x61 && ~x20 && x2 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && ~x11 && x12 && x61 && ~x20 && ~x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && ~x11 && x12 && ~x61 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && ~x11 && x12 && ~x61 && ~x1 && x4 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && ~x11 && x12 && ~x61 && ~x1 && ~x4 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && ~x11 && ~x12 && x61 && x13 && x1 && x3 && x6 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && ~x11 && ~x12 && x61 && x13 && x1 && x3 && ~x6 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && ~x11 && ~x12 && x61 && x13 && x1 && ~x3 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && ~x11 && ~x12 && x61 && x13 && ~x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && ~x11 && ~x12 && x61 && ~x13 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && ~x11 && ~x12 && ~x61 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s206;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && ~x11 && ~x12 && ~x61 && ~x1 && x2 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && ~x11 && ~x12 && ~x61 && ~x1 && ~x2 && x9 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x10 && ~x11 && ~x12 && ~x61 && ~x1 && ~x2 && ~x9 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && x62 && ~x64 && x14 && x30 && x43 )
						nx_state = s10;
					else if( ~x69 && x70 && x62 && ~x64 && x14 && x30 && ~x43 && x18 && x41 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && x62 && ~x64 && x14 && x30 && ~x43 && x18 && ~x41 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x70 && x62 && ~x64 && x14 && x30 && ~x43 && ~x18 && x34 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x70 && x62 && ~x64 && x14 && x30 && ~x43 && ~x18 && ~x34 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && x62 && ~x64 && x14 && ~x30 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && x62 && ~x64 && ~x14 && x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && x62 && ~x64 && ~x14 && ~x11 && x1 && x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && x62 && ~x64 && ~x14 && ~x11 && x1 && ~x2 && x3 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x70 && x62 && ~x64 && ~x14 && ~x11 && x1 && ~x2 && ~x3 )
						nx_state = s10;
					else if( ~x69 && x70 && x62 && ~x64 && ~x14 && ~x11 && ~x1 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x46 && x47 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x46 && x47 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x46 && ~x47 && x34 && x2 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s322;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x46 && ~x47 && x34 && ~x2 )
						nx_state = s10;
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x46 && ~x47 && ~x34 && x4 && x2 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x46 && ~x47 && ~x34 && x4 && ~x2 )
						nx_state = s10;
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x46 && ~x47 && ~x34 && ~x4 && x32 && x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x46 && ~x47 && ~x34 && ~x4 && x32 && ~x2 )
						nx_state = s10;
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x46 && ~x47 && ~x34 && ~x4 && ~x32 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x46 && ~x47 && ~x34 && ~x4 && ~x32 && ~x2 )
						nx_state = s10;
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x46 && x16 && x35 && x5 && x1 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x46 && x16 && x35 && x5 && ~x1 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x46 && x16 && x35 && ~x5 && x32 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x46 && x16 && x35 && ~x5 && ~x32 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x46 && x16 && ~x35 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x46 && x16 && ~x35 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x46 && ~x16 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && x15 && x11 && x25 && x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && x15 && x11 && x25 && ~x3 && x5 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && x15 && x11 && x25 && ~x3 && ~x5 )
						nx_state = s10;
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && x15 && x11 && ~x25 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && x15 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && ~x15 && x44 && x40 && x48 && x47 )
						nx_state = s10;
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && ~x15 && x44 && x40 && x48 && ~x47 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && ~x15 && x44 && x40 && ~x48 && x47 )
						nx_state = s10;
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && ~x15 && x44 && x40 && ~x48 && ~x47 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && ~x15 && x44 && ~x40 && x47 )
						nx_state = s10;
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && ~x15 && x44 && ~x40 && ~x47 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && ~x15 && x44 && ~x40 && ~x47 && ~x34 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && ~x15 && ~x44 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && x16 && x15 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && x16 && x15 && ~x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && x16 && ~x15 && x4 && x5 && x1 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && x16 && ~x15 && x4 && x5 && ~x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && x16 && ~x15 && x4 && ~x5 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && x16 && ~x15 && x4 && ~x5 && ~x1 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && x16 && ~x15 && ~x4 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && x16 && ~x15 && ~x4 && ~x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && ~x16 && x15 && x2 && x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s326;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && ~x16 && x15 && x2 && ~x3 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && ~x16 && x15 && x2 && ~x3 && ~x4 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && ~x16 && x15 && x2 && ~x3 && ~x4 && ~x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && ~x16 && x15 && ~x2 )
						nx_state = s10;
					else if( ~x69 && x70 && ~x62 && ~x63 && ~x16 && ~x15 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( ~x69 && ~x70 && x45 && x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && ~x70 && x45 && ~x11 && x1 && x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && ~x70 && x45 && ~x11 && x1 && ~x2 && x3 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && ~x70 && x45 && ~x11 && x1 && ~x2 && ~x3 )
						nx_state = s10;
					else if( ~x69 && ~x70 && x45 && ~x11 && ~x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && ~x45 && x11 && x25 && x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && ~x70 && ~x45 && x11 && x25 && ~x3 && x5 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && ~x70 && ~x45 && x11 && x25 && ~x3 && ~x5 )
						nx_state = s10;
					else if( ~x69 && ~x70 && ~x45 && x11 && ~x25 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else nx_state = s10;
				s11 : if( x69 && x70 && x62 && x25 && x7 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x70 && x62 && x25 && ~x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && x70 && x62 && ~x25 && x26 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && x70 && x62 && ~x25 && x26 && ~x7 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && x70 && x62 && ~x25 && ~x26 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && x70 && x62 && ~x25 && ~x26 && ~x12 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && x70 && ~x62 && x63 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 )
						begin
							y3 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s327;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x65 && x66 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x65 && x66 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x65 && x66 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x65 && x66 && ~x23 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x65 && ~x66 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x65 && ~x66 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x65 && ~x66 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x65 && ~x66 && ~x15 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && ~x65 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s328;
						end
					else if( x69 && ~x70 && x65 && x66 && x67 && x23 && x18 && x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && ~x70 && x65 && x66 && x67 && x23 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && ~x70 && x65 && x66 && x67 && x23 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x66 && x67 && x23 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x66 && x67 && ~x23 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && x61 && x60 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && x61 && x60 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && x61 && x60 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && x61 && x60 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && x61 && ~x60 && x62 && x2 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && x61 && ~x60 && x62 && ~x2 && x20 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	
							nx_state = s330;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && x61 && ~x60 && x62 && ~x2 && ~x20 && x16 && x11 && x12 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s278;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && x61 && ~x60 && x62 && ~x2 && ~x20 && x16 && x11 && ~x12 && x13 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s278;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && x61 && ~x60 && x62 && ~x2 && ~x20 && x16 && x11 && ~x12 && ~x13 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && x61 && ~x60 && x62 && ~x2 && ~x20 && x16 && ~x11 && x13 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s135;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && x61 && ~x60 && x62 && ~x2 && ~x20 && x16 && ~x11 && ~x13 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && x61 && ~x60 && x62 && ~x2 && ~x20 && ~x16 && x17 && x11 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && x61 && ~x60 && x62 && ~x2 && ~x20 && ~x16 && x17 && x11 && ~x13 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && x61 && ~x60 && x62 && ~x2 && ~x20 && ~x16 && x17 && ~x11 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && x61 && ~x60 && x62 && ~x2 && ~x20 && ~x16 && ~x17 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && x61 && ~x60 && ~x62 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && x61 && ~x60 && ~x62 && ~x7 )
						nx_state = s118;
					else if( x69 && ~x70 && x65 && x66 && ~x67 && ~x61 && x60 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && ~x61 && x60 && ~x7 )
						nx_state = s118;
					else if( x69 && ~x70 && x65 && x66 && ~x67 && ~x61 && ~x60 && x62 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && ~x61 && ~x60 && ~x62 )
						nx_state = s331;
					else if( x69 && ~x70 && x65 && ~x66 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && x65 && ~x66 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && ~x66 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && ~x66 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && x15 && x9 )
						begin
							y31 = 1'b1;	
							nx_state = s164;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && x15 && ~x9 && x6 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && x15 && ~x9 && ~x6 )
						begin
							y31 = 1'b1;	
							nx_state = s164;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && x9 && x8 )
						begin
							y31 = 1'b1;	
							nx_state = s164;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && x9 && ~x8 && x10 )
						begin
							y31 = 1'b1;	
							nx_state = s164;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && x9 && ~x8 && ~x10 && x18 && x14 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && x9 && ~x8 && ~x10 && x18 && ~x14 && x13 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && x9 && ~x8 && ~x10 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && x9 && ~x8 && ~x10 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && ~x9 && x8 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s164;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && ~x9 && x8 && ~x12 && x18 && x14 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && ~x9 && x8 && ~x12 && x18 && ~x14 && x13 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && ~x9 && x8 && ~x12 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && ~x9 && x8 && ~x12 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && ~x9 && ~x8 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s164;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && ~x9 && ~x8 && ~x11 && x18 && x14 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && ~x9 && ~x8 && ~x11 && x18 && ~x14 && x13 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && ~x9 && ~x8 && ~x11 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && ~x9 && ~x8 && ~x11 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && ~x15 && ~x16 && x6 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s333;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x22 && ~x15 && ~x16 && ~x6 )
						begin
							y31 = 1'b1;	
							nx_state = s164;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && ~x22 )
						begin
							y31 = 1'b1;	
							nx_state = s164;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x21 && x68 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x21 && ~x68 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x21 && ~x68 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x21 && ~x68 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x21 && ~x68 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && x22 && x68 && x17 && x10 && x15 && x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s334;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && x22 && x68 && x17 && x10 && x15 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && x22 && x68 && x17 && x10 && ~x15 && x16 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && x22 && x68 && x17 && x10 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && x22 && x68 && x17 && ~x10 && x6 )
						begin
							y13 = 1'b1;	y16 = 1'b1;	
							nx_state = s335;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && x22 && x68 && x17 && ~x10 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && x22 && x68 && ~x17 && x18 && x6 && x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && x22 && x68 && ~x17 && x18 && x6 && ~x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && x22 && x68 && ~x17 && x18 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && x22 && x68 && ~x17 && ~x18 && x6 && x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && x22 && x68 && ~x17 && ~x18 && x6 && ~x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s107;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && x22 && x68 && ~x17 && ~x18 && ~x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && x22 && ~x68 && x23 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && x22 && ~x68 && ~x23 && x18 && x14 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && x22 && ~x68 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && x22 && ~x68 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && x22 && ~x68 && ~x23 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && ~x22 && x68 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && ~x22 && x68 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && ~x22 && x68 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && ~x22 && x68 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x21 && ~x22 && ~x68 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && x20 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && ~x20 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && x21 && x9 && x3 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && x21 && x9 && ~x3 && x4 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && x21 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && x21 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && ~x22 )
						nx_state = s1;
					else if( ~x69 )
						nx_state = s1;
					else nx_state = s11;
				s12 : if( x69 && x70 && x64 && x7 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s337;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && x32 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s337;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && x15 && x14 && x13 && x5 )
						begin
							y6 = 1'b1;	y35 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s338;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && x15 && x14 && x13 && ~x5 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y27 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s339;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && x15 && x14 && ~x13 && x8 && x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s340;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && x15 && x14 && ~x13 && x8 && ~x5 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && x15 && x14 && ~x13 && ~x8 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && x15 && x14 && ~x13 && ~x8 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && x15 && x14 && ~x13 && ~x8 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && x15 && x14 && ~x13 && ~x8 && ~x10 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && x15 && ~x14 && x13 && x31 && x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s340;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && x15 && ~x14 && x13 && x31 && ~x5 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && x15 && ~x14 && x13 && ~x31 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && x15 && ~x14 && x13 && ~x31 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && x15 && ~x14 && x13 && ~x31 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && x15 && ~x14 && x13 && ~x31 && ~x10 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && x15 && ~x14 && ~x13 && x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s340;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && x15 && ~x14 && ~x13 && ~x5 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && ~x15 && x13 && x14 && x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s343;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && ~x15 && x13 && x14 && ~x5 )
						begin
							y53 = 1'b1;	
							nx_state = s344;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && ~x15 && x13 && ~x14 && x16 && x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s340;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && ~x15 && x13 && ~x14 && x16 && ~x5 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && ~x15 && x13 && ~x14 && ~x16 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && ~x15 && x13 && ~x14 && ~x16 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && ~x15 && x13 && ~x14 && ~x16 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && ~x15 && x13 && ~x14 && ~x16 && ~x10 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && ~x15 && ~x13 && x14 && x30 && x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s340;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && ~x15 && ~x13 && x14 && x30 && ~x5 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && ~x15 && ~x13 && x14 && ~x30 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && ~x15 && ~x13 && x14 && ~x30 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && ~x15 && ~x13 && x14 && ~x30 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && ~x15 && ~x13 && x14 && ~x30 && ~x10 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && x9 && ~x15 && ~x13 && ~x14 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s345;
						end
					else if( x69 && x70 && x64 && ~x7 && x33 && ~x32 && ~x9 )
						begin
							y6 = 1'b1;	y40 = 1'b1;	y41 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s346;
						end
					else if( x69 && x70 && x64 && ~x7 && ~x33 && x9 && x13 && x32 && x15 && x14 )
						begin
							y6 = 1'b1;	y35 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s338;
						end
					else if( x69 && x70 && x64 && ~x7 && ~x33 && x9 && x13 && x32 && x15 && ~x14 && x16 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s347;
						end
					else if( x69 && x70 && x64 && ~x7 && ~x33 && x9 && x13 && x32 && x15 && ~x14 && ~x16 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s348;
						end
					else if( x69 && x70 && x64 && ~x7 && ~x33 && x9 && x13 && x32 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s349;
						end
					else if( x69 && x70 && x64 && ~x7 && ~x33 && x9 && x13 && x32 && ~x15 && ~x14 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s350;
						end
					else if( x69 && x70 && x64 && ~x7 && ~x33 && x9 && x13 && ~x32 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y35 = 1'b1;	y40 = 1'b1;	
							nx_state = s351;
						end
					else if( x69 && x70 && x64 && ~x7 && ~x33 && x9 && ~x13 && x32 && x15 && x14 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s352;
						end
					else if( x69 && x70 && x64 && ~x7 && ~x33 && x9 && ~x13 && x32 && x15 && ~x14 && x17 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x7 && ~x33 && x9 && ~x13 && x32 && x15 && ~x14 && ~x17 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s353;
						end
					else if( x69 && x70 && x64 && ~x7 && ~x33 && x9 && ~x13 && x32 && ~x15 && x14 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s354;
						end
					else if( x69 && x70 && x64 && ~x7 && ~x33 && x9 && ~x13 && x32 && ~x15 && ~x14 && x18 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x7 && ~x33 && x9 && ~x13 && x32 && ~x15 && ~x14 && ~x18 )
						nx_state = s12;
					else if( x69 && x70 && x64 && ~x7 && ~x33 && x9 && ~x13 && ~x32 && x4 && x6 )
						begin
							y6 = 1'b1;	y35 = 1'b1;	y40 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s355;
						end
					else if( x69 && x70 && x64 && ~x7 && ~x33 && x9 && ~x13 && ~x32 && x4 && ~x6 )
						begin
							y15 = 1'b1;	
							nx_state = s22;
						end
					else if( x69 && x70 && x64 && ~x7 && ~x33 && x9 && ~x13 && ~x32 && ~x4 )
						begin
							y15 = 1'b1;	
							nx_state = s356;
						end
					else if( x69 && x70 && x64 && ~x7 && ~x33 && ~x9 )
						begin
							y6 = 1'b1;	y40 = 1'b1;	y41 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s346;
						end
					else if( x69 && x70 && ~x64 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x21 && x5 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( x69 && ~x70 && x66 && x21 && ~x5 && x19 && x15 && x10 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s274;
						end
					else if( x69 && ~x70 && x66 && x21 && ~x5 && x19 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x70 && x66 && x21 && ~x5 && x19 && x15 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s124;
						end
					else if( x69 && ~x70 && x66 && x21 && ~x5 && x19 && ~x15 && x16 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && x66 && x21 && ~x5 && x19 && ~x15 && ~x16 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s357;
						end
					else if( x69 && ~x70 && x66 && x21 && ~x5 && ~x19 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( x69 && ~x70 && x66 && ~x21 && x22 && x23 && x3 && x15 && x10 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s363;
						end
					else if( x69 && ~x70 && x66 && ~x21 && x22 && x23 && x3 && x15 && ~x10 && x12 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s358;
						end
					else if( x69 && ~x70 && x66 && ~x21 && x22 && x23 && x3 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( x69 && ~x70 && x66 && ~x21 && x22 && x23 && x3 && ~x15 && x16 && x10 && x12 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s361;
						end
					else if( x69 && ~x70 && x66 && ~x21 && x22 && x23 && x3 && ~x15 && x16 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s360;
						end
					else if( x69 && ~x70 && x66 && ~x21 && x22 && x23 && x3 && ~x15 && x16 && ~x10 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s361;
						end
					else if( x69 && ~x70 && x66 && ~x21 && x22 && x23 && x3 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s362;
						end
					else if( x69 && ~x70 && x66 && ~x21 && x22 && x23 && ~x3 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s363;
						end
					else if( x69 && ~x70 && x66 && ~x21 && x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && x66 && ~x21 && ~x22 && x15 && x4 && x7 )
						nx_state = s47;
					else if( x69 && ~x70 && x66 && ~x21 && ~x22 && x15 && x4 && ~x7 && x23 && x9 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s361;
						end
					else if( x69 && ~x70 && x66 && ~x21 && ~x22 && x15 && x4 && ~x7 && x23 && ~x9 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && ~x70 && x66 && ~x21 && ~x22 && x15 && x4 && ~x7 && ~x23 && x9 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s365;
						end
					else if( x69 && ~x70 && x66 && ~x21 && ~x22 && x15 && x4 && ~x7 && ~x23 && ~x9 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s363;
						end
					else if( x69 && ~x70 && x66 && ~x21 && ~x22 && x15 && ~x4 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x69 && ~x70 && x66 && ~x21 && ~x22 && ~x15 && x16 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x69 && ~x70 && x66 && ~x21 && ~x22 && ~x15 && ~x16 && x23 && x4 )
						begin
							y14 = 1'b1;	
							nx_state = s366;
						end
					else if( x69 && ~x70 && x66 && ~x21 && ~x22 && ~x15 && ~x16 && x23 && ~x4 )
						begin
							y14 = 1'b1;	
							nx_state = s124;
						end
					else if( x69 && ~x70 && x66 && ~x21 && ~x22 && ~x15 && ~x16 && ~x23 && x4 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s367;
						end
					else if( x69 && ~x70 && x66 && ~x21 && ~x22 && ~x15 && ~x16 && ~x23 && ~x4 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( x69 && ~x70 && ~x66 && x67 && x24 && x26 && x20 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x66 && x67 && x24 && x26 && ~x20 && x21 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x66 && x67 && x24 && x26 && ~x20 && ~x21 && x22 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x66 && x67 && x24 && x26 && ~x20 && ~x21 && ~x22 && x23 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x66 && x67 && x24 && x26 && ~x20 && ~x21 && ~x22 && ~x23 && x16 && x11 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( x69 && ~x70 && ~x66 && x67 && x24 && x26 && ~x20 && ~x21 && ~x22 && ~x23 && x16 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && ~x66 && x67 && x24 && x26 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && x13 && x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && ~x66 && x67 && x24 && x26 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && x13 && ~x11 && x12 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( x69 && ~x70 && ~x66 && x67 && x24 && x26 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && x13 && ~x11 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && ~x66 && x67 && x24 && x26 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && ~x13 && x11 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && ~x70 && ~x66 && x67 && x24 && x26 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && ~x13 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && ~x66 && x67 && x24 && x26 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s35;
						end
					else if( x69 && ~x70 && ~x66 && x67 && x24 && ~x26 && x16 && x11 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s368;
						end
					else if( x69 && ~x70 && ~x66 && x67 && x24 && ~x26 && x16 && x11 && ~x12 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( x69 && ~x70 && ~x66 && x67 && x24 && ~x26 && x16 && ~x11 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s300;
						end
					else if( x69 && ~x70 && ~x66 && x67 && x24 && ~x26 && ~x16 && x17 && x11 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x66 && x67 && x24 && ~x26 && ~x16 && x17 && x11 && ~x13 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s122;
						end
					else if( x69 && ~x70 && ~x66 && x67 && x24 && ~x26 && ~x16 && x17 && ~x11 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x66 && x67 && x24 && ~x26 && ~x16 && ~x17 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && x25 && x26 && x4 && x15 && x10 && x11 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && x25 && x26 && x4 && x15 && x10 && ~x11 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && x25 && x26 && x4 && x15 && x10 && ~x11 && ~x12 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s301;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && x25 && x26 && x4 && x15 && ~x10 && x12 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s369;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && x25 && x26 && x4 && x15 && ~x10 && ~x12 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && x25 && x26 && x4 && ~x15 && x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && x25 && x26 && x4 && ~x15 && ~x16 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && x25 && x26 && ~x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && x25 && ~x26 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && x25 && ~x26 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && x25 && ~x26 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && x25 && ~x26 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && x10 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && x10 && ~x12 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s300;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && ~x10 && x11 && x12 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s309;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && ~x10 && x11 && ~x12 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s300;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && ~x10 && ~x11 && x12 && x13 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s370;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && ~x10 && ~x11 && x12 && ~x13 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && ~x10 && ~x11 && x12 && ~x13 && x18 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && ~x10 && ~x11 && x12 && ~x13 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && ~x10 && ~x11 && ~x12 && x14 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s370;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && ~x10 && ~x11 && ~x12 && ~x14 && x18 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && ~x10 && ~x11 && ~x12 && ~x14 && x18 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && ~x10 && ~x11 && ~x12 && ~x14 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && x12 && x10 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && x12 && x10 && ~x2 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && x12 && x10 && ~x2 && ~x4 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s372;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && x12 && ~x10 && x11 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && x12 && ~x10 && ~x11 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && x12 && ~x10 && ~x11 && ~x2 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && x12 && ~x10 && ~x11 && ~x2 && ~x4 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s372;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && ~x12 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && ~x12 && ~x2 && x11 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && ~x12 && ~x2 && x11 && ~x4 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s372;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && ~x12 && ~x2 && ~x11 && x10 && x4 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && ~x12 && ~x2 && ~x11 && x10 && ~x4 )
						begin
							y14 = 1'b1;	
							nx_state = s124;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && ~x12 && ~x2 && ~x11 && ~x10 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && ~x12 && ~x2 && ~x11 && ~x10 && ~x4 )
						begin
							y8 = 1'b1;	y17 = 1'b1;	y23 = 1'b1;	
							nx_state = s303;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && x10 && x12 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && x10 && ~x12 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && ~x10 && x11 && x12 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s300;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && ~x10 && x11 && ~x12 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s309;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && ~x10 && ~x11 && x12 && x13 )
						begin
							y8 = 1'b1;	
							nx_state = s373;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && ~x10 && ~x11 && x12 && ~x13 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && ~x10 && ~x11 && x12 && ~x13 && x17 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && ~x10 && ~x11 && x12 && ~x13 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && ~x10 && ~x11 && ~x12 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s373;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && ~x10 && ~x11 && ~x12 && ~x14 && x17 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && ~x10 && ~x11 && ~x12 && ~x14 && x17 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && ~x10 && ~x11 && ~x12 && ~x14 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && x10 && x8 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && x10 && x8 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && x10 && x8 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && x10 && x8 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && x10 && ~x8 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && x10 && ~x8 && ~x3 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && x10 && ~x8 && ~x3 && ~x5 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && ~x10 && x7 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && ~x10 && x7 && ~x3 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && ~x10 && x7 && ~x3 && ~x5 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && ~x10 && ~x7 && x11 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && ~x10 && ~x7 && x11 && ~x3 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && ~x10 && ~x7 && x11 && ~x3 && ~x5 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && ~x10 && ~x7 && ~x11 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && ~x10 && ~x7 && ~x11 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && ~x10 && ~x7 && ~x11 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && ~x10 && ~x7 && ~x11 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && x10 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && x10 && ~x3 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && x10 && ~x3 && ~x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && x11 && x9 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && x11 && x9 && ~x3 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && x11 && x9 && ~x3 && ~x5 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && ~x11 && x8 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && ~x11 && x8 && ~x3 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && ~x11 && x8 && ~x3 && ~x5 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && x10 && x8 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && x10 && x8 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && x10 && x8 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && x10 && x8 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && x10 && ~x8 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && x10 && ~x8 && ~x2 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && x10 && ~x8 && ~x2 && ~x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && ~x10 && x7 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && ~x10 && x7 && ~x2 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && ~x10 && x7 && ~x2 && ~x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && ~x10 && ~x7 && x11 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && ~x10 && ~x7 && x11 && ~x2 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && ~x10 && ~x7 && x11 && ~x2 && ~x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && ~x10 && ~x7 && ~x11 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && ~x10 && ~x7 && ~x11 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && ~x10 && ~x7 && ~x11 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && ~x10 && ~x7 && ~x11 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && x10 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && x10 && ~x2 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s271;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && x10 && ~x2 && ~x4 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && x11 && x9 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && x11 && x9 && ~x2 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && x11 && x9 && ~x2 && ~x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && x11 && ~x9 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && x11 && ~x9 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && x11 && ~x9 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && x11 && ~x9 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && ~x11 && x8 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && ~x11 && x8 && ~x2 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && ~x11 && x8 && ~x2 && ~x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && ~x11 && ~x8 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && ~x11 && ~x8 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && ~x11 && ~x8 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && ~x11 && ~x8 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && ~x17 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && ~x17 && ~x2 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && ~x17 && ~x2 && ~x4 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s372;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && x12 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && x12 && ~x3 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && x12 && ~x3 && ~x5 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && x15 && x11 && x10 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && x15 && x11 && x10 && ~x3 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && x15 && x11 && x10 && ~x3 && ~x5 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && x15 && x11 && ~x10 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && x15 && ~x11 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && x15 && ~x11 && ~x3 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && x15 && ~x11 && ~x3 && ~x5 && x10 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s300;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && x15 && ~x11 && ~x3 && ~x5 && ~x10 )
						begin
							y14 = 1'b1;	
							nx_state = s124;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && ~x15 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && ~x15 && ~x3 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && ~x15 && ~x3 && ~x5 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && x68 && x12 && x7 && x19 && x17 )
						begin
							y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s374;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && x68 && x12 && x7 && x19 && ~x17 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s376;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && x68 && x12 && x7 && ~x19 && x20 )
						begin
							y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s374;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && x68 && x12 && x7 && ~x19 && ~x20 )
						begin
							y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s375;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && x68 && x12 && ~x7 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s376;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && x68 && ~x12 && x19 && x7 && x17 )
						begin
							y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s374;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && x68 && ~x12 && x19 && x7 && ~x17 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s377;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && x68 && ~x12 && x19 && ~x7 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s376;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && x68 && ~x12 && ~x19 && x20 && x17 && x14 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s376;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && x68 && ~x12 && ~x19 && x20 && x17 && ~x14 && x16 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s376;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && x68 && ~x12 && ~x19 && x20 && x17 && ~x14 && ~x16 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && x68 && ~x12 && ~x19 && x20 && ~x17 && x16 && x15 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s376;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && x68 && ~x12 && ~x19 && x20 && ~x17 && x16 && ~x15 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && x68 && ~x12 && ~x19 && x20 && ~x17 && ~x16 && x13 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s376;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && x68 && ~x12 && ~x19 && x20 && ~x17 && ~x16 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && x68 && ~x12 && ~x19 && ~x20 && x7 )
						begin
							y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s378;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && x68 && ~x12 && ~x19 && ~x20 && ~x7 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s376;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && ~x68 && x19 && x7 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y17 = 1'b1;	
							nx_state = s314;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && ~x68 && x19 && ~x7 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && x15 && x14 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && x15 && ~x14 && x16 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && x15 && ~x14 && ~x16 && x9 && x3 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && x15 && ~x14 && ~x16 && x9 && ~x3 && x4 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && x15 && ~x14 && ~x16 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && x15 && ~x14 && ~x16 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && ~x15 && x14 && x18 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && ~x15 && x14 && ~x18 && x9 && x3 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && ~x15 && x14 && ~x18 && x9 && ~x3 && x4 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && ~x15 && x14 && ~x18 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && ~x15 && x14 && ~x18 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && ~x15 && ~x14 && x17 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x9 && x3 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x9 && ~x3 && x4 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && ~x68 && ~x19 && ~x20 && x7 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && x21 && ~x68 && ~x19 && ~x20 && ~x7 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && x22 && x68 && x12 && x18 && x17 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s379;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && x22 && x68 && x12 && x18 && ~x17 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s380;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && x22 && x68 && x12 && ~x18 && x19 && x17 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s379;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && x22 && x68 && x12 && ~x18 && x19 && ~x17 && x3 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s381;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && x22 && x68 && x12 && ~x18 && x19 && ~x17 && ~x3 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s382;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && x22 && x68 && x12 && ~x18 && ~x19 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s379;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && x22 && x68 && ~x12 && x18 && x17 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s379;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && x22 && x68 && ~x12 && x18 && ~x17 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s6;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && x22 && x68 && ~x12 && ~x18 && x19 )
						begin
							y4 = 1'b1;	y21 = 1'b1;	
							nx_state = s377;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && x22 && x68 && ~x12 && ~x18 && ~x19 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && x22 && ~x68 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && x68 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && x13 && x20 && x15 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && x13 && x20 && ~x15 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && x13 && ~x20 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && x14 && x20 && x15 )
						begin
							y22 = 1'b1;	y25 = 1'b1;	
							nx_state = s315;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && x14 && x20 && ~x15 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	y23 = 1'b1;	
							nx_state = s383;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && x14 && ~x20 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && x20 && x15 && x6 )
						begin
							y8 = 1'b1;	
							nx_state = s373;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && x20 && x15 && ~x6 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && x20 && x15 && ~x6 && x4 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && x20 && x15 && ~x6 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && x20 && ~x15 && x5 )
						begin
							y8 = 1'b1;	
							nx_state = s373;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && x20 && ~x15 && ~x5 && x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && x20 && ~x15 && ~x5 && x4 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && x20 && ~x15 && ~x5 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && ~x20 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s384;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && ~x20 && ~x3 && x7 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y17 = 1'b1;	
							nx_state = s314;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && ~x20 && ~x3 && ~x7 && x15 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s358;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && ~x20 && ~x3 && ~x7 && ~x15 )
						begin
							y2 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s385;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s384;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && x14 && x18 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s315;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && x14 && ~x18 && x15 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s315;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && x14 && ~x18 && ~x15 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && x14 && ~x18 && ~x15 && x4 && ~x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && x14 && ~x18 && ~x15 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && x14 && ~x18 && ~x15 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && ~x14 && x15 && x16 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s315;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && ~x14 && x15 && ~x16 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && ~x14 && x15 && ~x16 && x4 && ~x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && ~x14 && x15 && ~x16 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && ~x14 && x15 && ~x16 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && ~x14 && ~x15 && x17 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s315;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && ~x14 && ~x15 && ~x17 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && ~x14 && ~x15 && ~x17 && x4 && ~x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && ~x14 && ~x15 && ~x17 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && ~x14 && ~x15 && ~x17 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && ~x20 && x7 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y17 = 1'b1;	
							nx_state = s314;
						end
					else if( x69 && ~x70 && ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && ~x20 && ~x7 )
						begin
							y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s386;
						end
					else if( ~x69 && x44 && x45 && x38 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && x44 && x45 && ~x38 && x41 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && x44 && x45 && ~x38 && ~x41 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s387;
						end
					else if( ~x69 && x44 && ~x45 && x4 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && x44 && ~x45 && ~x4 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x69 && ~x44 && x10 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && ~x44 && ~x10 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x44 && ~x10 && ~x4 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s387;
						end
					else nx_state = s12;
				s13 : if( x62 && x64 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x62 && x64 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x62 && x64 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x62 && x64 && ~x19 )
						nx_state = s1;
					else if( x62 && ~x64 && x18 && x17 && x19 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y17 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s389;
						end
					else if( x62 && ~x64 && x18 && x17 && ~x19 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x62 && ~x64 && x18 && ~x17 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x62 && ~x64 && ~x18 && x17 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x62 && ~x64 && ~x18 && ~x17 && x19 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x62 && ~x64 && ~x18 && ~x17 && ~x19 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x62 && x63 && x65 && x66 && x31 && x5 )
						begin
							y23 = 1'b1;	y51 = 1'b1;	y58 = 1'b1;	
							nx_state = s390;
						end
					else if( ~x62 && x63 && x65 && x66 && x31 && ~x5 && x22 )
						begin
							y51 = 1'b1;	
							nx_state = s391;
						end
					else if( ~x62 && x63 && x65 && x66 && x31 && ~x5 && ~x22 )
						begin
							y44 = 1'b1;	y45 = 1'b1;	
							nx_state = s392;
						end
					else if( ~x62 && x63 && x65 && x66 && ~x31 && x5 )
						begin
							y65 = 1'b1;	
							nx_state = s393;
						end
					else if( ~x62 && x63 && x65 && x66 && ~x31 && ~x5 )
						begin
							y71 = 1'b1;	
							nx_state = s394;
						end
					else if( ~x62 && x63 && x65 && ~x66 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y55 = 1'b1;	
							y58 = 1'b1;	y69 = 1'b1;	
							nx_state = s395;
						end
					else if( ~x62 && x63 && ~x65 )
						begin
							y32 = 1'b1;	y33 = 1'b1;	
							nx_state = s396;
						end
					else if( ~x62 && ~x63 )
						begin
							y2 = 1'b1;	y15 = 1'b1;	y31 = 1'b1;	
							nx_state = s397;
						end
					else nx_state = s13;
				s14 : if( x69 && x70 && x62 && x66 && x25 && x8 )
						begin
							y2 = 1'b1;	y19 = 1'b1;	
							nx_state = s398;
						end
					else if( x69 && x70 && x62 && x66 && x25 && ~x8 )
						begin
							y1 = 1'b1;	y17 = 1'b1;	
							nx_state = s398;
						end
					else if( x69 && x70 && x62 && x66 && ~x25 && x13 )
						begin
							y13 = 1'b1;	
							nx_state = s240;
						end
					else if( x69 && x70 && x62 && x66 && ~x25 && ~x13 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && x70 && x62 && ~x66 && x13 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && x62 && ~x66 && x13 && ~x11 && x6 && x4 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	
							nx_state = s231;
						end
					else if( x69 && x70 && x62 && ~x66 && x13 && ~x11 && x6 && ~x4 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x70 && x62 && ~x66 && x13 && ~x11 && ~x6 && x5 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	
							nx_state = s276;
						end
					else if( x69 && x70 && x62 && ~x66 && x13 && ~x11 && ~x6 && ~x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s6;
						end
					else if( x69 && x70 && x62 && ~x66 && ~x13 && x14 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x69 && x70 && x62 && ~x66 && ~x13 && ~x14 && x9 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x69 && x70 && x62 && ~x66 && ~x13 && ~x14 && ~x9 && x6 && x2 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x69 && x70 && x62 && ~x66 && ~x13 && ~x14 && ~x9 && x6 && ~x2 )
						nx_state = s14;
					else if( x69 && x70 && x62 && ~x66 && ~x13 && ~x14 && ~x9 && ~x6 && x8 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x69 && x70 && x62 && ~x66 && ~x13 && ~x14 && ~x9 && ~x6 && ~x8 )
						nx_state = s14;
					else if( x69 && x70 && ~x62 && x63 && x64 && x67 && x11 && x7 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x64 && x67 && x11 && ~x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && x67 && ~x11 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && x10 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && ~x10 && x15 && x7 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && ~x10 && x15 && ~x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && ~x10 && ~x15 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x64 && x65 && x66 && x7 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x64 && x65 && x66 && ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x64 && x65 && ~x66 && x15 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x64 && x65 && ~x66 && ~x15 && x13 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x64 && x65 && ~x66 && ~x15 && x13 && ~x11 && x6 && x4 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	
							nx_state = s231;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x64 && x65 && ~x66 && ~x15 && x13 && ~x11 && x6 && ~x4 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x64 && x65 && ~x66 && ~x15 && x13 && ~x11 && ~x6 && x5 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	
							nx_state = s276;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x64 && x65 && ~x66 && ~x15 && x13 && ~x11 && ~x6 && ~x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s6;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x64 && x65 && ~x66 && ~x15 && ~x13 && x14 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x64 && x65 && ~x66 && ~x15 && ~x13 && ~x14 && x9 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x64 && x65 && ~x66 && ~x15 && ~x13 && ~x14 && ~x9 && x6 && x2 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x64 && x65 && ~x66 && ~x15 && ~x13 && ~x14 && ~x9 && x6 && ~x2 )
						nx_state = s14;
					else if( x69 && x70 && ~x62 && x63 && ~x64 && x65 && ~x66 && ~x15 && ~x13 && ~x14 && ~x9 && ~x6 && x8 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x64 && x65 && ~x66 && ~x15 && ~x13 && ~x14 && ~x9 && ~x6 && ~x8 )
						nx_state = s14;
					else if( x69 && x70 && ~x62 && x63 && ~x64 && ~x65 && x66 && x11 )
						begin
							y14 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s401;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x64 && ~x65 && x66 && ~x11 )
						begin
							y10 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s402;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x64 && ~x65 && ~x66 && x12 )
						begin
							y17 = 1'b1;	
							nx_state = s98;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x64 && ~x65 && ~x66 && ~x12 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x64 && ~x65 && ~x66 && ~x12 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x64 && ~x65 && ~x66 && ~x12 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x64 && ~x65 && ~x66 && ~x12 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x6 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x6 && ~x7 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x6 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && x23 && x24 && x10 && x11 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && x23 && x24 && x10 && ~x11 && x12 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && x23 && x24 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && x23 && x24 && ~x10 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && x23 && ~x24 )
						begin
							y31 = 1'b1;	
							nx_state = s164;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && x9 && x10 && x24 && x11 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && x9 && x10 && x24 && ~x11 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && x9 && x10 && ~x24 && x8 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && x9 && x10 && ~x24 && ~x8 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && x9 && ~x10 && x24 && x13 && x14 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && x9 && ~x10 && x24 && x13 && ~x14 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && x9 && ~x10 && x24 && x13 && ~x14 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && x9 && ~x10 && x24 && x13 && ~x14 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && x9 && ~x10 && x24 && x13 && ~x14 && ~x20 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && x9 && ~x10 && x24 && ~x13 && x15 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && x9 && ~x10 && x24 && ~x13 && ~x15 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && x9 && ~x10 && x24 && ~x13 && ~x15 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && x9 && ~x10 && x24 && ~x13 && ~x15 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && x9 && ~x10 && x24 && ~x13 && ~x15 && ~x20 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && x9 && ~x10 && ~x24 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && x9 && ~x10 && ~x24 && ~x8 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && ~x9 && x24 && x16 && x17 && x18 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && ~x9 && x24 && x16 && x17 && ~x18 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && ~x9 && x24 && x16 && x17 && ~x18 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && ~x9 && x24 && x16 && x17 && ~x18 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && ~x9 && x24 && x16 && x17 && ~x18 && ~x20 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && ~x9 && x24 && x16 && ~x17 && x19 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && ~x9 && x24 && x16 && ~x17 && ~x19 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && ~x9 && x24 && x16 && ~x17 && ~x19 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && ~x9 && x24 && x16 && ~x17 && ~x19 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && ~x9 && x24 && x16 && ~x17 && ~x19 && ~x20 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && ~x9 && x24 && ~x16 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && ~x9 && ~x24 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && ~x9 && ~x24 && x8 && ~x10 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && x67 && ~x23 && ~x9 && ~x24 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s98;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && ~x67 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && ~x67 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && ~x67 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x66 && ~x67 && ~x23 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && ~x66 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x67 && x65 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x66 && x67 && x65 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x66 && x67 && x65 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x67 && x65 && x22 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x67 && x65 && ~x22 && x18 && x13 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && ~x70 && x66 && x67 && x65 && ~x22 && x18 && x13 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x66 && x67 && x65 && ~x22 && x18 && ~x13 && x12 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && ~x70 && x66 && x67 && x65 && ~x22 && x18 && ~x13 && x12 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x66 && x67 && x65 && ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x67 && x65 && ~x22 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x68 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x68 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x68 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x68 && x21 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x68 && ~x21 )
						begin
							y10 = 1'b1;	
							nx_state = s405;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x68 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x68 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x68 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x68 && x62 && ~x61 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x68 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x68 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x68 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x68 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x68 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x68 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x68 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && x65 && ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x66 && ~x67 && x65 && ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x66 && ~x67 && x65 && ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && x65 && ~x21 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && x21 && x68 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && x21 && x68 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && x21 && x68 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && x21 && x68 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && x21 && ~x68 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x68 && x22 && x9 && x7 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x68 && x22 && x9 && ~x7 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x68 && x22 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x68 && ~x22 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x68 && ~x22 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x68 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x68 && ~x22 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x68 && x23 && x22 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x68 && x23 && ~x22 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x68 && x23 && ~x22 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x68 && x23 && ~x22 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x68 && x23 && ~x22 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x68 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x21 && x67 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x21 && x67 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x21 && x67 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && x21 && x67 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && x21 && ~x67 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x21 && ~x67 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x21 && ~x67 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x21 && ~x67 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && x21 && ~x67 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x67 && x22 && x18 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x67 && x22 && x18 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x67 && x22 && x18 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x67 && x22 && x18 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x67 && x22 && ~x18 && x10 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s252;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x67 && x22 && ~x18 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x67 && x22 && ~x18 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x67 && x22 && ~x18 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x67 && x22 && ~x18 && ~x10 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x67 && ~x22 && x19 && x10 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s252;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x67 && ~x22 && x19 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x67 && ~x22 && x19 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x67 && ~x22 && x19 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x67 && ~x22 && x19 && ~x10 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x67 && ~x22 && ~x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x67 && ~x22 && ~x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x67 && ~x22 && ~x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x67 && ~x22 && ~x19 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x67 && x23 && x22 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x67 && x23 && x22 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x67 && x23 && x22 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x67 && x23 && x22 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x67 && x23 && x22 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x67 && x23 && ~x22 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s406;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x67 && ~x23 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s406;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x20 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else if( ~x69 && x70 && x7 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( ~x69 && ~x70 && x44 && x17 )
						begin
							y8 = 1'b1;	y17 = 1'b1;	
							nx_state = s408;
						end
					else if( ~x69 && ~x70 && x44 && ~x17 && x18 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && ~x70 && x44 && ~x17 && ~x18 )
						nx_state = s14;
					else if( ~x69 && ~x70 && ~x44 && x45 && x46 && x47 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( ~x69 && ~x70 && ~x44 && x45 && x46 && ~x47 && x10 )
						begin
							y8 = 1'b1;	y17 = 1'b1;	
							nx_state = s408;
						end
					else if( ~x69 && ~x70 && ~x44 && x45 && x46 && ~x47 && ~x10 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && ~x70 && ~x44 && x45 && x46 && ~x47 && ~x10 && ~x4 )
						nx_state = s14;
					else if( ~x69 && ~x70 && ~x44 && x45 && ~x46 && x12 && x7 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x44 && x45 && ~x46 && x12 && ~x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( ~x69 && ~x70 && ~x44 && x45 && ~x46 && ~x12 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x45 && x46 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x45 && ~x46 && x10 && x11 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x45 && ~x46 && x10 && ~x11 && x7 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x44 && ~x45 && ~x46 && x10 && ~x11 && ~x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x45 && ~x46 && ~x10 && x12 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x45 && ~x46 && ~x10 && ~x12 && x7 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x44 && ~x45 && ~x46 && ~x10 && ~x12 && ~x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else nx_state = s14;
				s15 : if( 1'b1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y37 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s409;
						end
					else nx_state = s15;
				s16 : if( x69 && x70 && x62 && x64 && x65 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x69 && x70 && x62 && x64 && x65 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x69 && x70 && x62 && x64 && x65 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( x69 && x70 && x62 && x64 && x65 && ~x21 )
						nx_state = s1;
					else if( x69 && x70 && x62 && x64 && ~x65 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x69 && x70 && x62 && x64 && ~x65 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x69 && x70 && x62 && x64 && ~x65 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && x62 && x64 && ~x65 && ~x19 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x64 && x66 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x66 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x66 && ~x8 && x9 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x66 && ~x8 && ~x9 && x10 && x6 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x66 && ~x8 && ~x9 && x10 && ~x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x66 && ~x8 && ~x9 && ~x10 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x66 && ~x8 && ~x9 && ~x10 && ~x11 )
						nx_state = s16;
					else if( x69 && x70 && ~x62 && x64 && x63 )
						begin
							y3 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s411;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && x66 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && x66 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && x66 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && x66 && ~x14 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && x20 && x9 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && x20 && ~x9 && x5 && x3 && x12 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && x20 && ~x9 && x5 && x3 && x12 && ~x8 && x7 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && x20 && ~x9 && x5 && x3 && x12 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && x20 && ~x9 && x5 && x3 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && x20 && ~x9 && x5 && ~x3 && x6 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && x20 && ~x9 && x5 && ~x3 && x6 && ~x7 && x12 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && x20 && ~x9 && x5 && ~x3 && x6 && ~x7 && x12 && ~x8 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && x20 && ~x9 && x5 && ~x3 && x6 && ~x7 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && x20 && ~x9 && x5 && ~x3 && ~x6 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && x20 && ~x9 && x5 && ~x3 && ~x6 && ~x8 && x12 && x7 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && x20 && ~x9 && x5 && ~x3 && ~x6 && ~x8 && x12 && ~x7 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && x20 && ~x9 && x5 && ~x3 && ~x6 && ~x8 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && x20 && ~x9 && ~x5 && x6 && x3 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && x20 && ~x9 && ~x5 && x6 && ~x3 )
						begin
							y21 = 1'b1;	y38 = 1'b1;	
							nx_state = s412;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && x20 && ~x9 && ~x5 && ~x6 && x3 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && x20 && ~x9 && ~x5 && ~x6 && ~x3 )
						begin
							y22 = 1'b1;	y29 = 1'b1;	
							nx_state = s412;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && ~x20 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && ~x20 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && ~x20 && ~x4 && ~x5 && x15 )
						begin
							y26 = 1'b1;	
							nx_state = s413;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x21 && ~x20 && ~x4 && ~x5 && ~x15 )
						begin
							y35 = 1'b1;	
							nx_state = s414;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && ~x4 && x20 && x9 && x8 && x7 && x6 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && ~x4 && x20 && x9 && x8 && x7 && ~x6 && x5 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && ~x4 && x20 && x9 && x8 && x7 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && ~x4 && x20 && x9 && x8 && ~x7 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && ~x4 && x20 && x9 && ~x8 && x10 )
						begin
							y21 = 1'b1;	y38 = 1'b1;	
							nx_state = s412;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && ~x4 && x20 && x9 && ~x8 && ~x10 )
						begin
							y22 = 1'b1;	y29 = 1'b1;	
							nx_state = s412;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && ~x4 && x20 && ~x9 && x8 && x10 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s415;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && ~x4 && x20 && ~x9 && x8 && ~x10 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s301;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && ~x4 && x20 && ~x9 && ~x8 && x10 && x11 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && ~x4 && x20 && ~x9 && ~x8 && x10 && ~x11 && x7 && x6 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && ~x4 && x20 && ~x9 && ~x8 && x10 && ~x11 && x7 && ~x6 && x5 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && ~x4 && x20 && ~x9 && ~x8 && x10 && ~x11 && x7 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && ~x4 && x20 && ~x9 && ~x8 && x10 && ~x11 && ~x7 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && ~x4 && x20 && ~x9 && ~x8 && ~x10 && x12 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && ~x4 && x20 && ~x9 && ~x8 && ~x10 && ~x12 && x7 && x6 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && ~x4 && x20 && ~x9 && ~x8 && ~x10 && ~x12 && x7 && ~x6 && x5 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && ~x4 && x20 && ~x9 && ~x8 && ~x10 && ~x12 && x7 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && ~x4 && x20 && ~x9 && ~x8 && ~x10 && ~x12 && ~x7 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && ~x4 && ~x20 && x6 )
						begin
							y26 = 1'b1;	
							nx_state = s413;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x21 && ~x4 && ~x20 && ~x6 )
						begin
							y30 = 1'b1;	
							nx_state = s416;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && ~x65 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && ~x65 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && ~x65 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && ~x65 && x22 && ~x23 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && ~x65 && ~x22 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && x63 && x66 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x66 && x65 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x66 && x65 && ~x15 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x66 && x65 && ~x15 && ~x8 && x9 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x66 && x65 && ~x15 && ~x8 && ~x9 && x10 && x6 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x66 && x65 && ~x15 && ~x8 && ~x9 && x10 && ~x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x66 && x65 && ~x15 && ~x8 && ~x9 && ~x10 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x66 && x65 && ~x15 && ~x8 && ~x9 && ~x10 && ~x11 )
						nx_state = s16;
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x66 && ~x65 && x23 && x22 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	y26 = 1'b1;	
							nx_state = s418;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x66 && ~x65 && x23 && ~x22 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	y26 = 1'b1;	
							nx_state = s419;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x66 && ~x65 && ~x23 && x22 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	y26 = 1'b1;	
							nx_state = s419;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x66 && ~x65 && ~x23 && ~x22 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	y26 = 1'b1;	
							nx_state = s418;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x63 && x67 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s420;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x63 && ~x67 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && x66 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && x66 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && x66 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && x66 && x22 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && x66 && ~x22 && x3 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && x66 && ~x22 && ~x3 && x19 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x69 && ~x70 && x65 && x67 && x66 && ~x22 && ~x3 && x19 && x15 && ~x8 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && x65 && x67 && x66 && ~x22 && ~x3 && x19 && ~x15 && x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s126;
						end
					else if( x69 && ~x70 && x65 && x67 && x66 && ~x22 && ~x3 && x19 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( x69 && ~x70 && x65 && x67 && x66 && ~x22 && ~x3 && ~x19 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x66 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && x68 && x20 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && x68 && x20 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && x68 && x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && x68 && x20 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && x68 && ~x20 && x21 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && x68 && ~x20 && ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && x68 && ~x20 && ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && x68 && ~x20 && ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && x68 && ~x20 && ~x21 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && x60 && x61 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && x60 && x61 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && x60 && x61 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && x60 && x61 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && x60 && ~x61 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && x60 && ~x61 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && x60 && ~x61 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && x60 && ~x61 && ~x18 )
						nx_state = s118;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && x62 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && ~x62 && ~x18 )
						nx_state = s118;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && ~x60 && ~x61 )
						nx_state = s47;
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && x21 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && x19 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && x19 && ~x18 )
						nx_state = s16;
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && ~x19 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							nx_state = s165;
						end
					else if( x69 && ~x70 && ~x65 && x68 && x21 && x6 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x65 && x68 && x21 && x6 && ~x18 )
						nx_state = s16;
					else if( x69 && ~x70 && ~x65 && x68 && x21 && ~x6 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && ~x65 && x68 && ~x21 && x4 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x65 && x68 && ~x21 && x4 && ~x18 )
						nx_state = s16;
					else if( x69 && ~x70 && ~x65 && x68 && ~x21 && ~x4 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x68 && x62 && ~x61 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && x63 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && ~x63 && x64 && x16 && x8 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && ~x63 && x64 && x16 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && ~x63 && x64 && ~x16 && x4 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && ~x63 && x64 && ~x16 && ~x4 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s299;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && ~x63 && ~x64 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x69 && x70 && x10 && x6 && x7 && x2 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s201;
						end
					else if( ~x69 && x70 && x10 && x6 && x7 && x2 && ~x3 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( ~x69 && x70 && x10 && x6 && x7 && x2 && ~x3 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x69 && x70 && x10 && x6 && x7 && ~x2 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && x10 && x6 && ~x7 && x8 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && x70 && x10 && x6 && ~x7 && ~x8 && x2 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s201;
						end
					else if( ~x69 && x70 && x10 && x6 && ~x7 && ~x8 && x2 && ~x3 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( ~x69 && x70 && x10 && x6 && ~x7 && ~x8 && x2 && ~x3 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x69 && x70 && x10 && x6 && ~x7 && ~x8 && ~x2 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && x10 && ~x6 && x2 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && x70 && x10 && ~x6 && ~x2 && x64 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( ~x69 && x70 && x10 && ~x6 && ~x2 && ~x64 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x10 && x11 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && x70 && ~x10 && x11 && ~x5 && x6 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x70 && ~x10 && x11 && ~x5 && ~x6 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && x70 && ~x10 && ~x11 && x64 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( ~x69 && x70 && ~x10 && ~x11 && ~x64 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x44 && x45 && x46 && x37 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x46 && ~x37 && x9 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x46 && ~x37 && ~x9 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x46 && x10 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x44 && x45 && ~x46 && ~x10 && x11 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x46 && ~x10 && x11 && ~x5 && x6 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x46 && ~x10 && x11 && ~x5 && ~x6 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x46 && ~x10 && ~x11 && x1 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x44 && x45 && ~x46 && ~x10 && ~x11 && ~x1 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x69 && ~x70 && ~x44 && x46 && x11 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && ~x70 && ~x44 && x46 && ~x11 && x9 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && ~x70 && ~x44 && x46 && ~x11 && ~x9 && x7 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x44 && x46 && ~x11 && ~x9 && ~x7 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x46 && x10 && x1 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x44 && ~x46 && x10 && ~x1 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x46 && ~x10 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x46 && ~x10 && ~x5 && x6 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x46 && ~x10 && ~x5 && ~x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else nx_state = s16;
				s17 : if( x69 && x70 && x62 && x66 && x18 && x17 && x19 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y17 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s389;
						end
					else if( x69 && x70 && x62 && x66 && x18 && x17 && ~x19 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x70 && x62 && x66 && x18 && ~x17 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x70 && x62 && x66 && ~x18 && x17 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && x70 && x62 && x66 && ~x18 && ~x17 && x19 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && x70 && x62 && x66 && ~x18 && ~x17 && ~x19 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x70 && x62 && ~x66 && x3 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s230;
						end
					else if( x69 && x70 && x62 && ~x66 && x3 && ~x2 )
						nx_state = s17;
					else if( x69 && x70 && x62 && ~x66 && ~x3 && x4 && x2 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	
							nx_state = s231;
						end
					else if( x69 && x70 && x62 && ~x66 && ~x3 && x4 && ~x2 )
						nx_state = s17;
					else if( x69 && x70 && x62 && ~x66 && ~x3 && ~x4 && x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x70 && x62 && ~x66 && ~x3 && ~x4 && ~x2 )
						nx_state = s17;
					else if( x69 && x70 && ~x62 && x65 && x63 && x66 && x67 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && x70 && ~x62 && x65 && x63 && x66 && ~x67 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x70 && ~x62 && x65 && x63 && ~x66 && x15 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s6;
						end
					else if( x69 && x70 && ~x62 && x65 && x63 && ~x66 && ~x15 && x3 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s230;
						end
					else if( x69 && x70 && ~x62 && x65 && x63 && ~x66 && ~x15 && x3 && ~x2 )
						nx_state = s17;
					else if( x69 && x70 && ~x62 && x65 && x63 && ~x66 && ~x15 && ~x3 && x4 && x2 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	
							nx_state = s231;
						end
					else if( x69 && x70 && ~x62 && x65 && x63 && ~x66 && ~x15 && ~x3 && x4 && ~x2 )
						nx_state = s17;
					else if( x69 && x70 && ~x62 && x65 && x63 && ~x66 && ~x15 && ~x3 && ~x4 && x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x70 && ~x62 && x65 && x63 && ~x66 && ~x15 && ~x3 && ~x4 && ~x2 )
						nx_state = s17;
					else if( x69 && x70 && ~x62 && x65 && ~x63 && x66 && x64 && x67 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x70 && ~x62 && x65 && ~x63 && x66 && x64 && ~x67 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x70 && ~x62 && x65 && ~x63 && x66 && ~x64 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x70 && ~x62 && x65 && ~x63 && ~x66 && x64 && x67 && x21 && x20 )
						begin
							y60 = 1'b1;	
							nx_state = s424;
						end
					else if( x69 && x70 && ~x62 && x65 && ~x63 && ~x66 && x64 && x67 && x21 && ~x20 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x70 && ~x62 && x65 && ~x63 && ~x66 && x64 && x67 && ~x21 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x70 && ~x62 && x65 && ~x63 && ~x66 && x64 && ~x67 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y62 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s425;
						end
					else if( x69 && x70 && ~x62 && x65 && ~x63 && ~x66 && ~x64 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s328;
						end
					else if( x69 && x70 && ~x62 && ~x65 && x63 && x66 && x67 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s328;
						end
					else if( x69 && x70 && ~x62 && ~x65 && x63 && x66 && ~x67 && x3 && x5 && x7 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s426;
						end
					else if( x69 && x70 && ~x62 && ~x65 && x63 && x66 && ~x67 && x3 && x5 && ~x7 && x1 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && x70 && ~x62 && ~x65 && x63 && x66 && ~x67 && x3 && x5 && ~x7 && x1 && ~x2 )
						nx_state = s17;
					else if( x69 && x70 && ~x62 && ~x65 && x63 && x66 && ~x67 && x3 && x5 && ~x7 && ~x1 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x69 && x70 && ~x62 && ~x65 && x63 && x66 && ~x67 && x3 && ~x5 && x6 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	
							nx_state = s427;
						end
					else if( x69 && x70 && ~x62 && ~x65 && x63 && x66 && ~x67 && x3 && ~x5 && ~x6 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s426;
						end
					else if( x69 && x70 && ~x62 && ~x65 && x63 && x66 && ~x67 && ~x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x70 && ~x62 && ~x65 && x63 && ~x66 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s328;
						end
					else if( x69 && x70 && ~x62 && ~x65 && ~x63 && x64 && x66 && x67 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s328;
						end
					else if( x69 && x70 && ~x62 && ~x65 && ~x63 && x64 && x66 && ~x67 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x70 && ~x62 && ~x65 && ~x63 && x64 && ~x66 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s328;
						end
					else if( x69 && x70 && ~x62 && ~x65 && ~x63 && ~x64 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s328;
						end
					else if( x69 && ~x70 && x65 && x21 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && x65 && ~x21 && x22 && x23 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && ~x70 && x65 && ~x21 && x22 && ~x23 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x70 && x65 && ~x21 && ~x22 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && x64 && x63 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && x64 && ~x63 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x64 && x63 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x64 && ~x63 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && x21 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s362;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x24 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && x10 && x26 && x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && x10 && x26 && ~x12 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && x10 && ~x26 && x12 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s304;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && x10 && ~x26 && ~x12 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && x11 && x26 && x12 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s304;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && x11 && x26 && ~x12 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && x11 && ~x26 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && x11 && ~x26 && ~x12 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s300;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && x12 && x13 && x26 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && x12 && x13 && ~x26 )
						begin
							y8 = 1'b1;	
							nx_state = s373;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && x12 && ~x13 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && x12 && ~x13 && x19 && ~x14 && x26 )
						nx_state = s17;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && x12 && ~x13 && x19 && ~x14 && ~x26 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && x12 && ~x13 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && ~x12 && x14 && x26 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && ~x12 && x14 && ~x26 )
						begin
							y8 = 1'b1;	
							nx_state = s373;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && ~x12 && ~x14 && x19 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && ~x12 && ~x14 && x19 && ~x13 && x26 )
						nx_state = s17;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && ~x12 && ~x14 && x19 && ~x13 && ~x26 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && ~x12 && ~x14 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && x10 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && x10 && ~x3 && x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && x10 && ~x3 && ~x1 && x11 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s309;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && x10 && ~x3 && ~x1 && ~x11 && x12 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s430;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && x10 && ~x3 && ~x1 && ~x11 && ~x12 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && ~x10 && x11 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && ~x10 && x11 && ~x12 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && ~x10 && ~x11 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && ~x10 && ~x11 && ~x3 && x12 && x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && ~x10 && ~x11 && ~x3 && x12 && ~x1 )
						begin
							y6 = 1'b1;	
							nx_state = s431;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && ~x10 && ~x11 && ~x3 && ~x12 && x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s432;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && ~x10 && ~x11 && ~x3 && ~x12 && ~x1 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && x10 && x5 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s369;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && x10 && ~x5 && x2 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s258;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && x10 && ~x5 && ~x2 && x11 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s433;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && x10 && ~x5 && ~x2 && ~x11 && x12 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s433;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && x10 && ~x5 && ~x2 && ~x11 && ~x12 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s309;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && ~x10 && x11 && x12 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && ~x10 && x11 && ~x12 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s433;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && ~x10 && ~x11 && x5 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s369;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && ~x10 && ~x11 && ~x5 && x2 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s258;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && ~x10 && ~x11 && ~x5 && ~x2 && x12 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s433;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && ~x10 && ~x11 && ~x5 && ~x2 && ~x12 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && x10 && x12 && x8 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && x10 && x12 && ~x8 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && x10 && x12 && ~x8 && ~x3 && x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && x10 && x12 && ~x8 && ~x3 && ~x1 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && x10 && ~x12 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && x12 && x7 && x11 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && x12 && x7 && x11 && ~x3 && x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && x12 && x7 && x11 && ~x3 && ~x1 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && x12 && x7 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && x12 && ~x7 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && x12 && ~x7 && ~x3 && x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && x12 && ~x7 && ~x3 && ~x1 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && ~x12 && x11 && x9 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && ~x12 && x11 && ~x9 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && ~x12 && x11 && ~x9 && ~x3 && x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && ~x12 && x11 && ~x9 && ~x3 && ~x1 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && ~x12 && ~x11 && x8 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && ~x12 && ~x11 && x8 && ~x3 && x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && ~x12 && ~x11 && x8 && ~x3 && ~x1 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && ~x12 && ~x11 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && ~x16 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && ~x16 && ~x3 && x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && ~x16 && ~x3 && ~x1 )
						begin
							y6 = 1'b1;	
							nx_state = s368;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && x5 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s369;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && x10 && x8 && x2 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s258;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && x10 && x8 && ~x2 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && x10 && ~x8 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && x10 && ~x8 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && x10 && ~x8 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && x10 && ~x8 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && ~x10 && x11 && x2 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s258;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && ~x10 && x11 && ~x2 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && ~x10 && ~x11 && x7 && x2 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s258;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && ~x10 && ~x11 && x7 && ~x2 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && ~x10 && ~x11 && ~x7 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && ~x10 && ~x11 && ~x7 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && ~x10 && ~x11 && ~x7 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && ~x10 && ~x11 && ~x7 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && x10 && x2 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s35;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && x10 && ~x2 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s258;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && x11 && x9 && x2 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s258;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && x11 && x9 && ~x2 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && x11 && ~x9 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && x11 && ~x9 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && x11 && ~x9 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && x11 && ~x9 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && ~x11 && x8 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && ~x11 && x8 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && ~x11 && x8 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && ~x11 && x8 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && ~x11 && ~x8 && x2 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s258;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && ~x11 && ~x8 && ~x2 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && ~x16 && x2 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s258;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && ~x16 && ~x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s101;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && ~x25 && x26 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x24 && ~x25 && ~x26 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s435;
						end
					else if( ~x69 && x70 && x15 && x62 && x16 && x1 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s436;
						end
					else if( ~x69 && x70 && x15 && x62 && x16 && ~x1 && x5 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s195;
						end
					else if( ~x69 && x70 && x15 && x62 && x16 && ~x1 && ~x5 && x6 && x2 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else if( ~x69 && x70 && x15 && x62 && x16 && ~x1 && ~x5 && x6 && x2 && ~x3 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && x15 && x62 && x16 && ~x1 && ~x5 && x6 && ~x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && x15 && x62 && x16 && ~x1 && ~x5 && ~x6 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && x70 && x15 && x62 && ~x16 && x7 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && x70 && x15 && x62 && ~x16 && ~x7 && x9 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && x70 && x15 && x62 && ~x16 && ~x7 && ~x9 && x10 && x6 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && x70 && x15 && x62 && ~x16 && ~x7 && ~x9 && x10 && ~x6 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s438;
						end
					else if( ~x69 && x70 && x15 && x62 && ~x16 && ~x7 && ~x9 && ~x10 && x11 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s436;
						end
					else if( ~x69 && x70 && x15 && x62 && ~x16 && ~x7 && ~x9 && ~x10 && ~x11 )
						nx_state = s17;
					else if( ~x69 && x70 && x15 && ~x62 && x63 && x64 && x16 && x32 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && x15 && ~x62 && x63 && x64 && x16 && ~x32 && x36 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x69 && x70 && x15 && ~x62 && x63 && x64 && x16 && ~x32 && ~x36 && x6 && x2 && x3 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s440;
						end
					else if( ~x69 && x70 && x15 && ~x62 && x63 && x64 && x16 && ~x32 && ~x36 && x6 && x2 && ~x3 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x69 && x70 && x15 && ~x62 && x63 && x64 && x16 && ~x32 && ~x36 && x6 && ~x2 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x69 && x70 && x15 && ~x62 && x63 && x64 && x16 && ~x32 && ~x36 && ~x6 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s441;
						end
					else if( ~x69 && x70 && x15 && ~x62 && x63 && x64 && ~x16 && x7 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s441;
						end
					else if( ~x69 && x70 && x15 && ~x62 && x63 && x64 && ~x16 && ~x7 && x9 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s441;
						end
					else if( ~x69 && x70 && x15 && ~x62 && x63 && x64 && ~x16 && ~x7 && ~x9 && x41 && x37 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && x70 && x15 && ~x62 && x63 && x64 && ~x16 && ~x7 && ~x9 && x41 && ~x37 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s442;
						end
					else if( ~x69 && x70 && x15 && ~x62 && x63 && x64 && ~x16 && ~x7 && ~x9 && ~x41 && x42 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && x15 && ~x62 && x63 && x64 && ~x16 && ~x7 && ~x9 && ~x41 && ~x42 )
						nx_state = s17;
					else if( ~x69 && x70 && x15 && ~x62 && x63 && ~x64 && x19 && x13 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s443;
						end
					else if( ~x69 && x70 && x15 && ~x62 && x63 && ~x64 && x19 && ~x13 && x32 && x18 && x12 )
						nx_state = s17;
					else if( ~x69 && x70 && x15 && ~x62 && x63 && ~x64 && x19 && ~x13 && x32 && x18 && ~x12 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x69 && x70 && x15 && ~x62 && x63 && ~x64 && x19 && ~x13 && x32 && ~x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && x70 && x15 && ~x62 && x63 && ~x64 && x19 && ~x13 && ~x32 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && x70 && x15 && ~x62 && x63 && ~x64 && ~x19 )
						nx_state = s1;
					else if( ~x69 && x70 && x15 && ~x62 && ~x63 && x16 && x1 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && x15 && ~x62 && ~x63 && x16 && ~x1 && x5 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x69 && x70 && x15 && ~x62 && ~x63 && x16 && ~x1 && ~x5 && x6 && x2 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s445;
						end
					else if( ~x69 && x70 && x15 && ~x62 && ~x63 && x16 && ~x1 && ~x5 && x6 && x2 && ~x3 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x69 && x70 && x15 && ~x62 && ~x63 && x16 && ~x1 && ~x5 && x6 && ~x2 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x69 && x70 && x15 && ~x62 && ~x63 && x16 && ~x1 && ~x5 && ~x6 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s441;
						end
					else if( ~x69 && x70 && x15 && ~x62 && ~x63 && ~x16 && x7 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s441;
						end
					else if( ~x69 && x70 && x15 && ~x62 && ~x63 && ~x16 && ~x7 && x9 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s441;
						end
					else if( ~x69 && x70 && x15 && ~x62 && ~x63 && ~x16 && ~x7 && ~x9 && x10 && x6 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && x70 && x15 && ~x62 && ~x63 && ~x16 && ~x7 && ~x9 && x10 && ~x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s446;
						end
					else if( ~x69 && x70 && x15 && ~x62 && ~x63 && ~x16 && ~x7 && ~x9 && ~x10 && x11 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && x15 && ~x62 && ~x63 && ~x16 && ~x7 && ~x9 && ~x10 && ~x11 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && x16 && x4 && x5 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( ~x69 && x70 && ~x15 && x62 && x16 && x4 && x5 && ~x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x69 && x70 && ~x15 && x62 && x16 && x4 && ~x5 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s436;
						end
					else if( ~x69 && x70 && ~x15 && x62 && x16 && ~x4 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s436;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && x3 && x11 && x2 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s447;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && x3 && x11 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && x3 && ~x11 && x4 && x12 && x13 && x2 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s448;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && x3 && ~x11 && x4 && x12 && x13 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && x3 && ~x11 && x4 && x12 && ~x13 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && x3 && ~x11 && x4 && ~x12 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && x3 && ~x11 && ~x4 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && x4 && x11 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s449;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && x4 && x11 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && x4 && ~x11 && x12 && x13 && x14 && x2 )
						begin
							y13 = 1'b1;	
							nx_state = s450;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && x4 && ~x11 && x12 && x13 && x14 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && x4 && ~x11 && x12 && x13 && ~x14 && x2 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s451;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && x4 && ~x11 && x12 && x13 && ~x14 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && x4 && ~x11 && x12 && ~x13 && x2 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s195;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && x4 && ~x11 && x12 && ~x13 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && x4 && ~x11 && ~x12 && x2 )
						begin
							y10 = 1'b1;	
							nx_state = s193;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && x4 && ~x11 && ~x12 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && x5 && x6 && x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s436;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && x5 && x6 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && x7 && x8 && x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s436;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && x7 && x8 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && x7 && ~x8 && x2 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && x7 && ~x8 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && x8 && x2 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && x8 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && ~x8 && x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s436;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && ~x8 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && x7 && x9 && x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s436;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && x7 && x9 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && x7 && ~x9 && x2 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && x7 && ~x9 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && x9 && x2 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && x9 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && ~x9 && x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s436;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && ~x9 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && x10 && x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s436;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && x10 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && ~x10 && x2 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && ~x10 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && x10 && x2 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && x10 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && ~x10 && x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s436;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && ~x10 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && x47 && x35 && x5 && x33 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && x47 && x35 && x5 && ~x33 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && x47 && x35 && x5 && ~x33 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && x47 && x35 && ~x5 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && x47 && ~x35 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && x34 && x42 && x2 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y12 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s452;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && x34 && x42 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && x34 && ~x42 && x3 && x4 && x12 && x13 && x2 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s453;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && x34 && ~x42 && x3 && x4 && x12 && x13 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && x34 && ~x42 && x3 && x4 && x12 && ~x13 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && x34 && ~x42 && x3 && x4 && ~x12 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && x34 && ~x42 && x3 && ~x4 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && x34 && ~x42 && ~x3 && x4 && x12 && x13 && x2 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && x34 && ~x42 && ~x3 && x4 && x12 && x13 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && x34 && ~x42 && ~x3 && x4 && x12 && ~x13 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && x34 && ~x42 && ~x3 && x4 && ~x12 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && x34 && ~x42 && ~x3 && ~x4 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && ~x34 && x33 && x35 && x11 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y29 = 1'b1;	
							nx_state = s288;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && ~x34 && x33 && x35 && ~x11 && x43 && x44 && x14 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && ~x34 && x33 && x35 && ~x11 && x43 && x44 && ~x14 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s322;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && ~x34 && x33 && x35 && ~x11 && x43 && ~x44 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && ~x34 && x33 && x35 && ~x11 && ~x43 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && ~x34 && x33 && ~x35 && x36 && x37 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && ~x34 && x33 && ~x35 && x36 && ~x37 && x38 && x39 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && ~x34 && x33 && ~x35 && x36 && ~x37 && x38 && ~x39 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s440;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && ~x34 && x33 && ~x35 && x36 && ~x37 && ~x38 && x8 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s440;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && ~x34 && x33 && ~x35 && x36 && ~x37 && ~x38 && ~x8 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && ~x34 && x33 && ~x35 && ~x36 && x6 && x7 && x9 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && ~x34 && x33 && ~x35 && ~x36 && x6 && x7 && ~x9 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s440;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && ~x34 && x33 && ~x35 && ~x36 && x6 && ~x7 && x40 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s440;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && ~x34 && x33 && ~x35 && ~x36 && x6 && ~x7 && ~x40 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && ~x34 && x33 && ~x35 && ~x36 && ~x6 && x38 && x41 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && ~x34 && x33 && ~x35 && ~x36 && ~x6 && x38 && ~x41 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s440;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && ~x34 && x33 && ~x35 && ~x36 && ~x6 && ~x38 && x10 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s440;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && ~x34 && x33 && ~x35 && ~x36 && ~x6 && ~x38 && ~x10 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 && ~x34 && ~x33 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && ~x64 && x17 && x19 && x10 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && ~x64 && x17 && x19 && ~x10 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && ~x64 && x17 && ~x19 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && ~x64 && ~x17 && x20 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && ~x64 && ~x17 && ~x20 && x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && ~x64 && ~x17 && ~x20 && ~x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && x16 && x4 && x5 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && x16 && x4 && x5 && ~x2 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && x16 && x4 && x5 && ~x2 && ~x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && x16 && x4 && ~x5 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && x16 && ~x4 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && x3 && x11 && x2 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s447;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && x3 && x11 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && x3 && ~x11 && x4 && x12 && x13 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s455;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && x3 && ~x11 && x4 && x12 && x13 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && x3 && ~x11 && x4 && x12 && ~x13 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && x3 && ~x11 && x4 && ~x12 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && x3 && ~x11 && ~x4 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && x4 && x11 && x2 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s456;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && x4 && x11 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && x4 && ~x11 && x12 && x13 && x14 && x2 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && x4 && ~x11 && x12 && x13 && x14 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && x4 && ~x11 && x12 && x13 && ~x14 && x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s326;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && x4 && ~x11 && x12 && x13 && ~x14 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && x4 && ~x11 && x12 && ~x13 && x2 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && x4 && ~x11 && x12 && ~x13 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && x4 && ~x11 && ~x12 && x2 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && x4 && ~x11 && ~x12 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && x5 && x6 && x2 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && x5 && x6 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && x7 && x8 && x2 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && x7 && x8 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && x7 && ~x8 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s445;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && x7 && ~x8 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && x8 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s445;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && x8 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && ~x8 && x2 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && ~x8 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && x7 && x9 && x2 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && x7 && x9 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && x7 && ~x9 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s445;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && x7 && ~x9 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && x9 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s445;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && x9 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && ~x9 && x2 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && ~x9 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && x10 && x2 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && x10 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && ~x10 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s445;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && ~x10 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && x10 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s445;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && x10 && ~x2 )
						nx_state = s17;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && ~x10 && x2 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && ~x10 && ~x2 )
						nx_state = s17;
					else if( ~x69 && ~x70 && x44 && x45 && x46 && x29 && x41 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x46 && x29 && ~x41 )
						nx_state = s17;
					else if( ~x69 && ~x70 && x44 && x45 && x46 && ~x29 && x14 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x44 && x45 && x46 && ~x29 && ~x14 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x46 && x11 && x10 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x44 && x45 && ~x46 && x11 && ~x10 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x46 && ~x11 && x10 && x12 && x4 && x1 )
						nx_state = s17;
					else if( ~x69 && ~x70 && x44 && x45 && ~x46 && ~x11 && x10 && x12 && x4 && ~x1 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x46 && ~x11 && x10 && x12 && ~x4 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x46 && ~x11 && x10 && ~x12 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x46 && ~x11 && ~x10 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x46 && x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x46 && ~x2 )
						nx_state = s17;
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x46 && x47 && x19 && x13 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s443;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x46 && x47 && x19 && ~x13 && x21 && x18 && x12 )
						nx_state = s17;
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x46 && x47 && x19 && ~x13 && x21 && x18 && ~x12 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x46 && x47 && x19 && ~x13 && x21 && ~x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x46 && x47 && x19 && ~x13 && ~x21 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x46 && x47 && ~x19 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x46 && ~x47 && x12 && x15 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x46 && ~x47 && x12 && ~x15 )
						nx_state = s17;
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x46 && ~x47 && ~x12 && x3 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x46 && ~x47 && ~x12 && ~x3 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && ~x44 && x45 && x46 && x47 && x1 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x44 && x45 && x46 && x47 && ~x1 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x44 && x45 && x46 && ~x47 && x10 && x2 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && ~x70 && ~x44 && x45 && x46 && ~x47 && x10 && ~x2 )
						nx_state = s17;
					else if( ~x69 && ~x70 && ~x44 && x45 && x46 && ~x47 && ~x10 && x3 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x44 && x45 && x46 && ~x47 && ~x10 && ~x3 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && ~x44 && x45 && ~x46 && x10 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( ~x69 && ~x70 && ~x44 && x45 && ~x46 && ~x10 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x45 && x3 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x44 && ~x45 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else nx_state = s17;
				s18 : if( x70 && x62 && x65 && x4 && x5 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s18;
						end
					else if( x70 && x62 && x65 && x4 && x5 && ~x1 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( x70 && x62 && x65 && x4 && ~x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x70 && x62 && x65 && ~x4 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( x70 && x62 && ~x65 && x3 && x1 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	
							nx_state = s457;
						end
					else if( x70 && x62 && ~x65 && x3 && ~x1 && x4 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	
							nx_state = s457;
						end
					else if( x70 && x62 && ~x65 && x3 && ~x1 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s18;
						end
					else if( x70 && x62 && ~x65 && ~x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( x70 && ~x62 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x21 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x22 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( ~x70 && ~x21 && ~x22 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s269;
						end
					else nx_state = s18;
				s19 : if( x65 && x6 && x4 && x5 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s18;
						end
					else if( x65 && x6 && x4 && x5 && ~x1 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( x65 && x6 && x4 && ~x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x65 && x6 && ~x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( x65 && ~x6 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y8 = 1'b1;	
							nx_state = s2;
						end
					else if( ~x65 && ~x5 && x2 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s459;
						end
					else if( ~x65 && ~x5 && x2 && ~x1 )
						begin
							y3 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							nx_state = s460;
						end
					else if( ~x65 && ~x5 && ~x2 && x1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s461;
						end
					else if( ~x65 && ~x5 && ~x2 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y8 = 1'b1;	
							nx_state = s2;
						end
					else nx_state = s19;
				s20 : if( x65 && x4 && x5 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s18;
						end
					else if( x65 && x4 && x5 && ~x1 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( x65 && x4 && ~x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x65 && ~x4 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && x17 && x18 && x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	
							nx_state = s20;
						end
					else if( ~x65 && x17 && x18 && ~x1 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && x17 && x18 && ~x1 && ~x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x65 && x17 && ~x18 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x65 && ~x17 && x18 && x2 && x19 && x4 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x65 && ~x17 && x18 && x2 && x19 && ~x4 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && ~x17 && x18 && x2 && ~x19 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && ~x17 && x18 && ~x2 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && ~x17 && ~x18 && x19 && x2 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && ~x17 && ~x18 && x19 && ~x2 )
						nx_state = s1;
					else if( ~x65 && ~x17 && ~x18 && ~x19 && x1 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x65 && ~x17 && ~x18 && ~x19 && x1 && ~x3 && x4 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( ~x65 && ~x17 && ~x18 && ~x19 && x1 && ~x3 && ~x4 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && ~x17 && ~x18 && ~x19 && ~x1 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else nx_state = s20;
				s21 : if( x69 && x70 && x62 && x64 )
						begin
							y3 = 1'b1;	
							nx_state = s462;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x3 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && ~x3 && x4 && x5 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s18;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && ~x3 && x4 && x5 && ~x1 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && ~x3 && x4 && ~x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && ~x3 && ~x4 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && x66 && x4 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && x66 && x4 && ~x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && x66 && ~x4 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s18;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && ~x3 && x1 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s46;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && ~x3 && x1 && ~x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && ~x3 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( x69 && x70 && ~x62 && x65 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y14 = 1'b1;	
							y16 = 1'b1;	y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s463;
						end
					else if( x69 && x70 && ~x62 && ~x65 )
						begin
							y14 = 1'b1;	
							nx_state = s124;
						end
					else if( x69 && ~x70 && x65 && x66 && x67 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && x21 && x20 )
						begin
							y9 = 1'b1;	y24 = 1'b1;	
							nx_state = s464;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && x21 && ~x20 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x67 && ~x21 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && x65 && ~x66 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( x69 && ~x70 && ~x65 && x20 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && ~x65 && ~x20 && x21 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y21 = 1'b1;	
							nx_state = s121;
						end
					else if( x69 && ~x70 && ~x65 && ~x20 && ~x21 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( ~x69 && x7 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s206;
						end
					else if( ~x69 && ~x7 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else nx_state = s21;
				s22 : if( x62 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s466;
						end
					else if( ~x62 && x21 && x20 )
						begin
							y7 = 1'b1;	y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s467;
						end
					else if( ~x62 && x21 && ~x20 )
						begin
							y28 = 1'b1;	
							nx_state = s468;
						end
					else if( ~x62 && ~x21 && x20 )
						begin
							y28 = 1'b1;	
							nx_state = s469;
						end
					else if( ~x62 && ~x21 && ~x20 )
						begin
							y7 = 1'b1;	y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s467;
						end
					else nx_state = s22;
				s23 : if( x33 && x32 && x10 && x11 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s470;
						end
					else if( x33 && x32 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s470;
						end
					else if( x33 && x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x33 && x32 && ~x10 )
						nx_state = s1;
					else if( x33 && ~x32 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s471;
						end
					else if( ~x33 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s471;
						end
					else nx_state = s23;
				s24 : if( x13 && x10 && x11 && x12 && x4 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s27;
						end
					else if( x13 && x10 && x11 && x12 && ~x4 )
						nx_state = s24;
					else if( x13 && x10 && x11 && ~x12 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x13 && x10 && x11 && ~x12 && ~x3 && x2 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s30;
						end
					else if( x13 && x10 && x11 && ~x12 && ~x3 && ~x2 )
						nx_state = s24;
					else if( x13 && x10 && ~x11 && x12 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x13 && x10 && ~x11 && x12 && ~x3 && x2 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s30;
						end
					else if( x13 && x10 && ~x11 && x12 && ~x3 && ~x2 )
						nx_state = s24;
					else if( x13 && x10 && ~x11 && ~x12 && x14 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x13 && x10 && ~x11 && ~x12 && x14 && ~x3 && x2 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s30;
						end
					else if( x13 && x10 && ~x11 && ~x12 && x14 && ~x3 && ~x2 )
						nx_state = s24;
					else if( x13 && x10 && ~x11 && ~x12 && ~x14 )
						begin
							y16 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							nx_state = s472;
						end
					else if( x13 && ~x10 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x13 && ~x10 && ~x3 && x2 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s30;
						end
					else if( x13 && ~x10 && ~x3 && ~x2 )
						nx_state = s24;
					else if( ~x13 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( ~x13 && ~x3 && x2 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s30;
						end
					else if( ~x13 && ~x3 && ~x2 )
						nx_state = s24;
					else nx_state = s24;
				s25 : if( x10 && x12 && x4 && x11 && x3 && x13 )
						begin
							y16 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							nx_state = s472;
						end
					else if( x10 && x12 && x4 && x11 && x3 && ~x13 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s473;
						end
					else if( x10 && x12 && x4 && x11 && ~x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x10 && x12 && x4 && ~x11 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x10 && x12 && ~x4 )
						nx_state = s25;
					else if( x10 && ~x12 && x13 && x11 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s24;
						end
					else if( x10 && ~x12 && x13 && ~x11 && x14 && x4 && x3 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s30;
						end
					else if( x10 && ~x12 && x13 && ~x11 && x14 && x4 && ~x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x10 && ~x12 && x13 && ~x11 && x14 && ~x4 )
						nx_state = s25;
					else if( x10 && ~x12 && x13 && ~x11 && ~x14 )
						nx_state = s1;
					else if( x10 && ~x12 && ~x13 && x14 && x4 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x10 && ~x12 && ~x13 && x14 && ~x4 )
						nx_state = s25;
					else if( x10 && ~x12 && ~x13 && ~x14 )
						nx_state = s1;
					else if( ~x10 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s24;
						end
					else nx_state = s25;
				s26 : if( x11 && x12 && x2 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	
							nx_state = s474;
						end
					else if( x11 && x12 && ~x2 )
						nx_state = s26;
					else if( x11 && ~x12 && x3 )
						nx_state = s1;
					else if( x11 && ~x12 && ~x3 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( ~x11 && x3 )
						nx_state = s1;
					else if( ~x11 && ~x3 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else nx_state = s26;
				s27 : if( x12 )
						begin
							y15 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s475;
						end
					else if( ~x12 && x11 && x13 && x7 )
						nx_state = s1;
					else if( ~x12 && x11 && x13 && ~x7 )
						begin
							y15 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s475;
						end
					else if( ~x12 && x11 && ~x13 )
						begin
							y15 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s475;
						end
					else if( ~x12 && ~x11 && x14 )
						begin
							y15 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s475;
						end
					else if( ~x12 && ~x11 && ~x14 && x7 )
						nx_state = s1;
					else if( ~x12 && ~x11 && ~x14 && ~x7 )
						begin
							y15 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s475;
						end
					else nx_state = s27;
				s28 : if( x12 && x11 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x12 && x11 && ~x3 && x2 )
						nx_state = s1;
					else if( x12 && x11 && ~x3 && ~x2 )
						nx_state = s28;
					else if( x12 && ~x11 && x10 )
						begin
							y15 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s475;
						end
					else if( x12 && ~x11 && ~x10 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x12 && ~x11 && ~x10 && ~x3 && x2 )
						nx_state = s1;
					else if( x12 && ~x11 && ~x10 && ~x3 && ~x2 )
						nx_state = s28;
					else if( ~x12 && x13 && x11 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( ~x12 && x13 && x11 && ~x3 && x2 )
						nx_state = s1;
					else if( ~x12 && x13 && x11 && ~x3 && ~x2 )
						nx_state = s28;
					else if( ~x12 && x13 && ~x11 && x14 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( ~x12 && x13 && ~x11 && x14 && ~x3 && x2 )
						nx_state = s1;
					else if( ~x12 && x13 && ~x11 && x14 && ~x3 && ~x2 )
						nx_state = s28;
					else if( ~x12 && x13 && ~x11 && ~x14 && x10 && x5 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	
							nx_state = s474;
						end
					else if( ~x12 && x13 && ~x11 && ~x14 && x10 && ~x5 && x1 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s476;
						end
					else if( ~x12 && x13 && ~x11 && ~x14 && x10 && ~x5 && ~x1 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( ~x12 && x13 && ~x11 && ~x14 && ~x10 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( ~x12 && x13 && ~x11 && ~x14 && ~x10 && ~x3 && x2 )
						nx_state = s1;
					else if( ~x12 && x13 && ~x11 && ~x14 && ~x10 && ~x3 && ~x2 )
						nx_state = s28;
					else if( ~x12 && ~x13 && x14 && x10 )
						begin
							y15 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s475;
						end
					else if( ~x12 && ~x13 && x14 && ~x10 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( ~x12 && ~x13 && x14 && ~x10 && ~x3 && x2 )
						nx_state = s1;
					else if( ~x12 && ~x13 && x14 && ~x10 && ~x3 && ~x2 )
						nx_state = s28;
					else if( ~x12 && ~x13 && ~x14 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( ~x12 && ~x13 && ~x14 && ~x3 && x2 )
						nx_state = s1;
					else if( ~x12 && ~x13 && ~x14 && ~x3 && ~x2 )
						nx_state = s28;
					else nx_state = s28;
				s29 : if( x12 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s28;
						end
					else if( ~x12 && x10 && x13 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x12 && x10 && x13 && ~x11 && x14 && x6 && x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x12 && x10 && x13 && ~x11 && x14 && x6 && ~x2 )
						nx_state = s29;
					else if( ~x12 && x10 && x13 && ~x11 && x14 && ~x6 && x2 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x12 && x10 && x13 && ~x11 && x14 && ~x6 && ~x2 )
						nx_state = s29;
					else if( ~x12 && x10 && x13 && ~x11 && ~x14 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s28;
						end
					else if( ~x12 && x10 && ~x13 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s28;
						end
					else if( ~x12 && ~x10 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s28;
						end
					else nx_state = s29;
				s30 : if( x10 && x12 )
						begin
							y16 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							nx_state = s472;
						end
					else if( x10 && ~x12 && x11 && x13 )
						begin
							y16 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							nx_state = s472;
						end
					else if( x10 && ~x12 && x11 && ~x13 && x14 )
						begin
							y16 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							nx_state = s472;
						end
					else if( x10 && ~x12 && x11 && ~x13 && ~x14 && x1 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s33;
						end
					else if( x10 && ~x12 && x11 && ~x13 && ~x14 && ~x1 && x2 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x10 && ~x12 && x11 && ~x13 && ~x14 && ~x1 && ~x2 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s476;
						end
					else if( x10 && ~x12 && ~x11 && x13 && x14 && x6 && x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x10 && ~x12 && ~x11 && x13 && x14 && x6 && ~x2 )
						nx_state = s30;
					else if( x10 && ~x12 && ~x11 && x13 && x14 && ~x6 && x2 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x10 && ~x12 && ~x11 && x13 && x14 && ~x6 && ~x2 )
						nx_state = s30;
					else if( x10 && ~x12 && ~x11 && x13 && ~x14 )
						begin
							y16 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							nx_state = s472;
						end
					else if( x10 && ~x12 && ~x11 && ~x13 )
						begin
							y16 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							nx_state = s472;
						end
					else if( ~x10 )
						begin
							y16 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							nx_state = s472;
						end
					else nx_state = s30;
				s31 : if( x62 && x10 && x12 )
						nx_state = s1;
					else if( x62 && x10 && ~x12 && x13 && x11 && x4 && x2 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s33;
						end
					else if( x62 && x10 && ~x12 && x13 && x11 && x4 && ~x2 )
						nx_state = s31;
					else if( x62 && x10 && ~x12 && x13 && x11 && ~x4 && x2 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s30;
						end
					else if( x62 && x10 && ~x12 && x13 && x11 && ~x4 && ~x2 )
						nx_state = s31;
					else if( x62 && x10 && ~x12 && x13 && ~x11 && x14 )
						nx_state = s1;
					else if( x62 && x10 && ~x12 && x13 && ~x11 && ~x14 && x1 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s24;
						end
					else if( x62 && x10 && ~x12 && x13 && ~x11 && ~x14 && ~x1 )
						begin
							y16 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							nx_state = s472;
						end
					else if( x62 && x10 && ~x12 && ~x13 && x14 )
						nx_state = s1;
					else if( x62 && x10 && ~x12 && ~x13 && ~x14 && x4 && x2 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s33;
						end
					else if( x62 && x10 && ~x12 && ~x13 && ~x14 && x4 && ~x2 )
						nx_state = s31;
					else if( x62 && x10 && ~x12 && ~x13 && ~x14 && ~x4 && x2 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s30;
						end
					else if( x62 && x10 && ~x12 && ~x13 && ~x14 && ~x4 && ~x2 )
						nx_state = s31;
					else if( x62 && ~x10 && x4 && x2 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s33;
						end
					else if( x62 && ~x10 && x4 && ~x2 )
						nx_state = s31;
					else if( x62 && ~x10 && ~x4 && x2 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s30;
						end
					else if( x62 && ~x10 && ~x4 && ~x2 )
						nx_state = s31;
					else if( ~x62 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x62 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x62 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x62 && ~x14 )
						nx_state = s1;
					else nx_state = s31;
				s32 : if( x10 && x12 && x11 && x13 && x3 && x6 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s24;
						end
					else if( x10 && x12 && x11 && x13 && x3 && ~x6 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x10 && x12 && x11 && x13 && ~x3 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x10 && x12 && x11 && ~x13 && x5 )
						begin
							y5 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s26;
						end
					else if( x10 && x12 && x11 && ~x13 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x10 && x12 && ~x11 && x5 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s28;
						end
					else if( x10 && x12 && ~x11 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x10 && ~x12 && x13 && x11 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s31;
						end
					else if( x10 && ~x12 && x13 && ~x11 && x14 && x5 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s29;
						end
					else if( x10 && ~x12 && x13 && ~x11 && x14 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x10 && ~x12 && x13 && ~x11 && ~x14 && x8 && x1 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s28;
						end
					else if( x10 && ~x12 && x13 && ~x11 && ~x14 && x8 && ~x1 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x10 && ~x12 && x13 && ~x11 && ~x14 && ~x8 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s28;
						end
					else if( x10 && ~x12 && ~x13 && x14 && x5 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s28;
						end
					else if( x10 && ~x12 && ~x13 && x14 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x10 && ~x12 && ~x13 && ~x14 && x1 )
						begin
							y5 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s26;
						end
					else if( x10 && ~x12 && ~x13 && ~x14 && ~x1 && x3 )
						nx_state = s1;
					else if( x10 && ~x12 && ~x13 && ~x14 && ~x1 && ~x3 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( ~x10 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s31;
						end
					else nx_state = s32;
				s33 : if( x12 && x11 && x10 && x13 && x2 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s476;
						end
					else if( x12 && x11 && x10 && x13 && ~x2 )
						nx_state = s33;
					else if( x12 && x11 && x10 && ~x13 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s476;
						end
					else if( x12 && x11 && ~x10 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s476;
						end
					else if( x12 && ~x11 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s476;
						end
					else if( ~x12 && x14 && x11 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s476;
						end
					else if( ~x12 && x14 && ~x11 && x10 && x13 && x2 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s476;
						end
					else if( ~x12 && x14 && ~x11 && x10 && x13 && ~x2 )
						nx_state = s33;
					else if( ~x12 && x14 && ~x11 && x10 && ~x13 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s476;
						end
					else if( ~x12 && x14 && ~x11 && ~x10 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s476;
						end
					else if( ~x12 && ~x14 && x13 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s476;
						end
					else if( ~x12 && ~x14 && ~x13 && x10 && x2 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( ~x12 && ~x14 && ~x13 && x10 && ~x2 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s476;
						end
					else if( ~x12 && ~x14 && ~x13 && ~x10 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s476;
						end
					else nx_state = s33;
				s34 : if( x69 && x70 && x62 && x4 && x5 && x1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s477;
						end
					else if( x69 && x70 && x62 && x4 && x5 && ~x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s60;
						end
					else if( x69 && x70 && x62 && x4 && ~x5 && x1 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( x69 && x70 && x62 && x4 && ~x5 && ~x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x69 && x70 && x62 && ~x4 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s479;
						end
					else if( x69 && x70 && ~x62 && x64 && x63 && x16 && x15 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( x69 && x70 && ~x62 && x64 && x63 && x16 && ~x15 && x4 && x5 && x1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s477;
						end
					else if( x69 && x70 && ~x62 && x64 && x63 && x16 && ~x15 && x4 && x5 && ~x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s60;
						end
					else if( x69 && x70 && ~x62 && x64 && x63 && x16 && ~x15 && x4 && ~x5 && x1 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( x69 && x70 && ~x62 && x64 && x63 && x16 && ~x15 && x4 && ~x5 && ~x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x69 && x70 && ~x62 && x64 && x63 && x16 && ~x15 && ~x4 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( x69 && x70 && ~x62 && x64 && x63 && ~x16 && x15 && x3 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( x69 && x70 && ~x62 && x64 && x63 && ~x16 && x15 && x3 && ~x2 )
						nx_state = s34;
					else if( x69 && x70 && ~x62 && x64 && x63 && ~x16 && x15 && ~x3 && x4 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s60;
						end
					else if( x69 && x70 && ~x62 && x64 && x63 && ~x16 && x15 && ~x3 && x4 && ~x2 )
						nx_state = s34;
					else if( x69 && x70 && ~x62 && x64 && x63 && ~x16 && x15 && ~x3 && ~x4 && x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( x69 && x70 && ~x62 && x64 && x63 && ~x16 && x15 && ~x3 && ~x4 && ~x2 )
						nx_state = s34;
					else if( x69 && x70 && ~x62 && x64 && x63 && ~x16 && ~x15 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s477;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && x66 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && x66 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && x66 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && x66 && ~x14 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x67 && x21 && x20 )
						begin
							y60 = 1'b1;	
							nx_state = s424;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x67 && x21 && ~x20 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && x67 && ~x21 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x65 && ~x66 && ~x67 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s481;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && ~x65 && x67 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s482;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && ~x65 && ~x67 && x18 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && ~x65 && ~x67 && ~x18 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && ~x65 && ~x67 && ~x18 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && ~x65 && ~x67 && ~x18 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && ~x65 && ~x67 && ~x18 && ~x9 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && x63 && x65 )
						begin
							y63 = 1'b1;	
							nx_state = s483;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x65 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x65 && ~x7 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x63 && x65 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x63 && x65 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x63 && x65 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && ~x63 && x65 && ~x23 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && ~x63 && ~x65 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x63 && ~x65 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x63 && ~x65 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && ~x63 && ~x65 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x67 && x65 && x22 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	
							nx_state = s486;
						end
					else if( x69 && ~x70 && x66 && x67 && x65 && ~x22 && x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && x66 && x67 && x65 && ~x22 && ~x23 && x18 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x66 && x67 && x65 && ~x22 && ~x23 && x18 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x66 && x67 && x65 && ~x22 && ~x23 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x67 && x65 && ~x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && x15 && x64 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && x15 && x64 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && x15 && ~x64 && x16 && x8 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && x15 && ~x64 && x16 && x8 && ~x14 && x7 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s296;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && x15 && ~x64 && x16 && x8 && ~x14 && ~x7 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && x15 && ~x64 && x16 && x8 && ~x14 && ~x7 && ~x12 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && x15 && ~x64 && x16 && ~x8 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && x15 && ~x64 && x16 && ~x8 && ~x14 && x7 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s297;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && x15 && ~x64 && x16 && ~x8 && ~x14 && ~x7 && x13 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && x15 && ~x64 && x16 && ~x8 && ~x14 && ~x7 && ~x13 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && x15 && ~x64 && ~x16 && x7 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s298;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && x15 && ~x64 && ~x16 && ~x7 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && x15 && ~x64 && ~x16 && ~x7 && ~x3 && x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && x15 && ~x64 && ~x16 && ~x7 && ~x3 && ~x5 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && x15 && ~x64 && ~x16 && ~x7 && ~x3 && ~x5 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && x16 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && x8 && x7 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && x8 && x7 && ~x3 && x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && x8 && x7 && ~x3 && ~x5 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && x8 && ~x7 && x9 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && x8 && ~x7 && x9 && ~x3 && x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && x8 && ~x7 && x9 && ~x3 && ~x5 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && x8 && ~x7 && ~x9 && x3 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && x8 && ~x7 && ~x9 && ~x3 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && ~x8 && x7 && x11 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && ~x8 && x7 && x11 && ~x3 && x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && ~x8 && x7 && x11 && ~x3 && ~x5 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && ~x8 && x7 && ~x11 && x3 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && ~x8 && x7 && ~x11 && ~x3 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && ~x8 && ~x7 && x10 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && ~x8 && ~x7 && x10 && ~x3 && x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && ~x8 && ~x7 && x10 && ~x3 && ~x5 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && ~x8 && ~x7 && ~x10 && x3 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && ~x8 && ~x7 && ~x10 && ~x3 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && ~x16 && x64 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s299;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && ~x16 && ~x64 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && ~x16 && ~x64 && ~x3 && x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && x63 && ~x15 && ~x16 && ~x64 && ~x3 && ~x5 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y28 = 1'b1;	
							nx_state = s299;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x63 && x64 && x19 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x63 && x64 && x19 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x63 && x64 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x63 && x64 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x67 && ~x65 && ~x63 && ~x64 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x61 && x60 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x61 && x60 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x61 && x60 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x61 && x60 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x61 && ~x60 && x62 && x11 && x13 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x61 && ~x60 && x62 && x11 && x13 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x61 && ~x60 && x62 && x11 && x13 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x61 && ~x60 && x62 && x11 && x13 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x61 && ~x60 && x62 && x11 && ~x13 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x61 && ~x60 && x62 && ~x11 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x61 && ~x60 && x62 && ~x11 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x61 && ~x60 && x62 && ~x11 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x61 && ~x60 && x62 && ~x11 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x61 && ~x60 && ~x62 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x69 && ~x70 && x66 && ~x67 && x65 && x61 && ~x60 && ~x62 && ~x7 )
						nx_state = s118;
					else if( x69 && ~x70 && x66 && ~x67 && x65 && ~x61 && x60 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x69 && ~x70 && x66 && ~x67 && x65 && ~x61 && x60 && ~x7 )
						nx_state = s118;
					else if( x69 && ~x70 && x66 && ~x67 && x65 && ~x61 && ~x60 && x62 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x69 && ~x70 && x66 && ~x67 && x65 && ~x61 && ~x60 && ~x62 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s487;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && x21 && x68 && x9 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && x21 && x68 && x9 && ~x8 && x7 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && x21 && x68 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && x21 && x68 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && x21 && ~x68 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && x21 && ~x68 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && x21 && ~x68 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && x21 && ~x68 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && x5 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && x17 && x10 && x15 && x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s334;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && x17 && x10 && x15 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && x17 && x10 && ~x15 && x16 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && x17 && x10 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && x17 && ~x10 && x6 )
						begin
							y13 = 1'b1;	y16 = 1'b1;	
							nx_state = s335;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && x17 && ~x10 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && ~x17 && x18 && x6 && x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && ~x17 && x18 && x6 && ~x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && ~x17 && x18 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && ~x17 && ~x18 && x6 && x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && ~x17 && ~x18 && x6 && ~x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s107;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && ~x17 && ~x18 && ~x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && x23 && x18 && x15 && x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && x23 && x18 && x15 && ~x10 && x12 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && x23 && x18 && x15 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s366;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && x23 && x18 && ~x15 && x16 && x10 && x12 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && x23 && x18 && ~x15 && x16 && x10 && ~x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && x23 && x18 && ~x15 && x16 && ~x10 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && x23 && x18 && ~x15 && ~x16 )
						nx_state = s47;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && x23 && ~x18 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && ~x23 && x18 && x14 )
						nx_state = s47;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s47;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && ~x23 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && x10 && x15 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && x10 && ~x15 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && ~x10 && x15 && x6 && x14 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && ~x10 && x15 && x6 && ~x14 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s488;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && ~x10 && x15 && ~x6 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && ~x10 && x15 && ~x6 && x4 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && ~x10 && x15 && ~x6 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && ~x10 && ~x15 && x5 && x14 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s253;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && ~x10 && ~x15 && x5 && ~x14 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s488;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && ~x10 && ~x15 && ~x5 && x4 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && ~x10 && ~x15 && ~x5 && x4 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && ~x10 && ~x15 && ~x5 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && x14 && x10 )
						begin
							y13 = 1'b1;	y16 = 1'b1;	
							nx_state = s489;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && x14 && ~x10 && x15 )
						begin
							y13 = 1'b1;	y16 = 1'b1;	
							nx_state = s335;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && x14 && ~x10 && ~x15 )
						begin
							y12 = 1'b1;	
							nx_state = s490;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && ~x14 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && ~x14 && ~x2 && x15 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && ~x14 && ~x2 && x15 && ~x3 && x10 )
						begin
							y12 = 1'b1;	
							nx_state = s244;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && ~x14 && ~x2 && x15 && ~x3 && ~x10 )
						begin
							y12 = 1'b1;	
							nx_state = s491;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && ~x14 && ~x2 && ~x15 && x10 && x3 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	
							nx_state = s268;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && ~x14 && ~x2 && ~x15 && x10 && ~x3 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && ~x14 && ~x2 && ~x15 && ~x10 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && ~x14 && ~x2 && ~x15 && ~x10 && ~x3 )
						begin
							y14 = 1'b1;	y16 = 1'b1;	
							nx_state = s492;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && x10 && x15 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && x10 && x15 && ~x3 )
						begin
							y12 = 1'b1;	
							nx_state = s490;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && x10 && ~x15 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && x15 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && x15 && ~x3 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && x13 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && x13 && ~x3 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && ~x13 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && ~x13 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && ~x13 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && ~x13 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && x12 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && x12 && ~x3 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && ~x12 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && ~x12 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && ~x12 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && x11 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && x11 && ~x3 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && ~x11 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && ~x11 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && ~x11 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && ~x17 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && ~x17 && ~x3 && x10 )
						begin
							y12 = 1'b1;	
							nx_state = s493;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && ~x17 && ~x3 && ~x10 )
						begin
							y12 = 1'b1;	
							nx_state = s245;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && ~x68 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && ~x68 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && ~x68 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && ~x68 && x23 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x67 && ~x65 && ~x21 && ~x22 && ~x68 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x15 && x9 && x21 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x15 && x9 && ~x21 && x23 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x15 && x9 && ~x21 && ~x23 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s494;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x15 && ~x9 && x21 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x15 && ~x9 && ~x21 && x23 && x6 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x15 && ~x9 && ~x21 && x23 && ~x6 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x15 && ~x9 && ~x21 && ~x23 && x6 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x15 && ~x9 && ~x21 && ~x23 && ~x6 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s494;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && x21 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s333;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && x23 && x9 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && x23 && ~x9 && x12 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && x23 && ~x9 && ~x12 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && x23 && ~x9 && ~x12 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && x23 && ~x9 && ~x12 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && x23 && ~x9 && ~x12 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && ~x23 && x9 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s494;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && ~x23 && ~x9 && x12 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s494;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && ~x23 && ~x9 && ~x12 && x18 && x14 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && ~x23 && ~x9 && ~x12 && x18 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && ~x23 && ~x9 && ~x12 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && ~x23 && ~x9 && ~x12 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && x23 && x9 && x10 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && x23 && x9 && ~x10 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && x23 && x9 && ~x10 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && x23 && x9 && ~x10 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && x23 && x9 && ~x10 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && x23 && ~x9 && x11 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && x23 && ~x9 && ~x11 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && x23 && ~x9 && ~x11 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && x23 && ~x9 && ~x11 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && x23 && ~x9 && ~x11 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && ~x23 && x9 && x10 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s494;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && ~x23 && x9 && ~x10 && x18 && x14 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && ~x23 && x9 && ~x10 && x18 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && ~x23 && x9 && ~x10 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && ~x23 && x9 && ~x10 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && ~x23 && ~x9 && x11 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s494;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && ~x23 && ~x9 && ~x11 && x18 && x14 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && ~x23 && ~x9 && ~x11 && x18 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && ~x23 && ~x9 && ~x11 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && ~x23 && ~x9 && ~x11 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && ~x16 && x23 && x6 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s495;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && ~x16 && x23 && ~x6 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && ~x16 && ~x23 && x6 )
						begin
							y31 = 1'b1;	
							nx_state = s164;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x15 && ~x21 && ~x16 && ~x23 && ~x6 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s494;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x24 && x26 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x24 && x26 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x24 && x26 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x24 && x26 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x24 && ~x26 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x24 && x25 && x26 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x24 && x25 && x26 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x24 && x25 && x26 && x19 && ~x14 && ~x13 )
						nx_state = s34;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x24 && x25 && x26 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x24 && x25 && ~x26 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x24 && ~x25 && x26 && x16 && x10 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x24 && ~x25 && x26 && x16 && ~x10 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x24 && ~x25 && x26 && x16 && ~x10 && ~x11 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x24 && ~x25 && x26 && x16 && ~x10 && ~x11 && ~x12 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x24 && ~x25 && x26 && ~x16 && x17 && x10 && x12 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s497;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x24 && ~x25 && x26 && ~x16 && x17 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x24 && ~x25 && x26 && ~x16 && x17 && ~x10 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s497;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x24 && ~x25 && x26 && ~x16 && ~x17 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x24 && ~x25 && ~x26 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x69 && x70 && x63 && x55 && x10 && x39 && x46 && x51 && x36 )
						nx_state = s34;
					else if( ~x69 && x70 && x63 && x55 && x10 && x39 && x46 && x51 && ~x36 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s498;
						end
					else if( ~x69 && x70 && x63 && x55 && x10 && x39 && x46 && ~x51 && x36 )
						nx_state = s34;
					else if( ~x69 && x70 && x63 && x55 && x10 && x39 && x46 && ~x51 && ~x36 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && x70 && x63 && x55 && x10 && x39 && ~x46 && x36 )
						nx_state = s34;
					else if( ~x69 && x70 && x63 && x55 && x10 && x39 && ~x46 && ~x36 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && x70 && x63 && x55 && x10 && ~x39 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( ~x69 && x70 && x63 && x55 && ~x10 && x42 && x34 && x8 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && x70 && x63 && x55 && ~x10 && x42 && x34 && ~x8 && x36 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s498;
						end
					else if( ~x69 && x70 && x63 && x55 && ~x10 && x42 && x34 && ~x8 && ~x36 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( ~x69 && x70 && x63 && x55 && ~x10 && x42 && ~x34 && x32 && x7 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && x70 && x63 && x55 && ~x10 && x42 && ~x34 && x32 && ~x7 && x54 && x36 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s498;
						end
					else if( ~x69 && x70 && x63 && x55 && ~x10 && x42 && ~x34 && x32 && ~x7 && x54 && ~x36 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( ~x69 && x70 && x63 && x55 && ~x10 && x42 && ~x34 && x32 && ~x7 && ~x54 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && x70 && x63 && x55 && ~x10 && x42 && ~x34 && ~x32 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x69 && x70 && x63 && x55 && ~x10 && ~x42 && x43 && x20 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && x70 && x63 && x55 && ~x10 && ~x42 && x43 && ~x20 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( ~x69 && x70 && x63 && x55 && ~x10 && ~x42 && x43 && ~x20 && ~x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s503;
						end
					else if( ~x69 && x70 && x63 && x55 && ~x10 && ~x42 && ~x43 && x13 && x32 && x3 && x6 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s504;
						end
					else if( ~x69 && x70 && x63 && x55 && ~x10 && ~x42 && ~x43 && x13 && x32 && x3 && ~x6 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( ~x69 && x70 && x63 && x55 && ~x10 && ~x42 && ~x43 && x13 && x32 && ~x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( ~x69 && x70 && x63 && x55 && ~x10 && ~x42 && ~x43 && x13 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && x70 && x63 && x55 && ~x10 && ~x42 && ~x43 && ~x13 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && x70 && x63 && ~x55 && x41 && x11 && x1 && x33 && x34 && x35 )
						nx_state = s34;
					else if( ~x69 && x70 && x63 && ~x55 && x41 && x11 && x1 && x33 && x34 && ~x35 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( ~x69 && x70 && x63 && ~x55 && x41 && x11 && x1 && x33 && ~x34 && x4 && x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && x70 && x63 && ~x55 && x41 && x11 && x1 && x33 && ~x34 && x4 && ~x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x69 && x70 && x63 && ~x55 && x41 && x11 && x1 && x33 && ~x34 && ~x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s503;
						end
					else if( ~x69 && x70 && x63 && ~x55 && x41 && x11 && x1 && ~x33 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && x70 && x63 && ~x55 && x41 && x11 && ~x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( ~x69 && x70 && x63 && ~x55 && x41 && ~x11 && x12 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && x70 && x63 && ~x55 && x41 && ~x11 && ~x12 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s504;
						end
					else if( ~x69 && x70 && x63 && ~x55 && ~x41 && x32 && x42 )
						begin
							y23 = 1'b1;	y25 = 1'b1;	y32 = 1'b1;	
							nx_state = s505;
						end
					else if( ~x69 && x70 && x63 && ~x55 && ~x41 && x32 && ~x42 && x43 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s503;
						end
					else if( ~x69 && x70 && x63 && ~x55 && ~x41 && x32 && ~x42 && ~x43 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y33 = 1'b1;	
							nx_state = s506;
						end
					else if( ~x69 && x70 && x63 && ~x55 && ~x41 && ~x32 && x11 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s503;
						end
					else if( ~x69 && x70 && x63 && ~x55 && ~x41 && ~x32 && x11 && ~x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( ~x69 && x70 && x63 && ~x55 && ~x41 && ~x32 && ~x11 && x12 && x35 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( ~x69 && x70 && x63 && ~x55 && ~x41 && ~x32 && ~x11 && x12 && ~x35 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( ~x69 && x70 && x63 && ~x55 && ~x41 && ~x32 && ~x11 && ~x12 && x33 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( ~x69 && x70 && x63 && ~x55 && ~x41 && ~x32 && ~x11 && ~x12 && ~x33 && x40 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( ~x69 && x70 && x63 && ~x55 && ~x41 && ~x32 && ~x11 && ~x12 && ~x33 && ~x40 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( ~x69 && x70 && ~x63 && x10 && x64 && x40 && x39 && x46 && x51 && x36 )
						nx_state = s34;
					else if( ~x69 && x70 && ~x63 && x10 && x64 && x40 && x39 && x46 && x51 && ~x36 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s507;
						end
					else if( ~x69 && x70 && ~x63 && x10 && x64 && x40 && x39 && x46 && ~x51 && x36 )
						nx_state = s34;
					else if( ~x69 && x70 && ~x63 && x10 && x64 && x40 && x39 && x46 && ~x51 && ~x36 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && x70 && ~x63 && x10 && x64 && x40 && x39 && ~x46 && x36 )
						nx_state = s34;
					else if( ~x69 && x70 && ~x63 && x10 && x64 && x40 && x39 && ~x46 && ~x36 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && x70 && ~x63 && x10 && x64 && x40 && ~x39 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x69 && x70 && ~x63 && x10 && x64 && ~x40 && x11 && x1 && x2 && x4 && x5 && x3 )
						nx_state = s34;
					else if( ~x69 && x70 && ~x63 && x10 && x64 && ~x40 && x11 && x1 && x2 && x4 && x5 && ~x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && x70 && ~x63 && x10 && x64 && ~x40 && x11 && x1 && x2 && x4 && ~x5 && x3 )
						nx_state = s34;
					else if( ~x69 && x70 && ~x63 && x10 && x64 && ~x40 && x11 && x1 && x2 && x4 && ~x5 && ~x3 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x69 && x70 && ~x63 && x10 && x64 && ~x40 && x11 && x1 && x2 && ~x4 && x3 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x70 && ~x63 && x10 && x64 && ~x40 && x11 && x1 && x2 && ~x4 && ~x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x69 && x70 && ~x63 && x10 && x64 && ~x40 && x11 && x1 && ~x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && x70 && ~x63 && x10 && x64 && ~x40 && x11 && ~x1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && x70 && ~x63 && x10 && x64 && ~x40 && ~x11 && x12 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && x70 && ~x63 && x10 && x64 && ~x40 && ~x11 && ~x12 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s510;
						end
					else if( ~x69 && x70 && ~x63 && x10 && ~x64 && x44 && x39 && x46 && x51 && x36 )
						nx_state = s34;
					else if( ~x69 && x70 && ~x63 && x10 && ~x64 && x44 && x39 && x46 && x51 && ~x36 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s511;
						end
					else if( ~x69 && x70 && ~x63 && x10 && ~x64 && x44 && x39 && x46 && ~x51 && x36 )
						nx_state = s34;
					else if( ~x69 && x70 && ~x63 && x10 && ~x64 && x44 && x39 && x46 && ~x51 && ~x36 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else if( ~x69 && x70 && ~x63 && x10 && ~x64 && x44 && x39 && ~x46 && x36 )
						nx_state = s34;
					else if( ~x69 && x70 && ~x63 && x10 && ~x64 && x44 && x39 && ~x46 && ~x36 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s513;
						end
					else if( ~x69 && x70 && ~x63 && x10 && ~x64 && x44 && ~x39 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x69 && x70 && ~x63 && x10 && ~x64 && ~x44 && x11 && x36 && x34 && x4 && x5 && x3 )
						nx_state = s34;
					else if( ~x69 && x70 && ~x63 && x10 && ~x64 && ~x44 && x11 && x36 && x34 && x4 && x5 && ~x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else if( ~x69 && x70 && ~x63 && x10 && ~x64 && ~x44 && x11 && x36 && x34 && x4 && ~x5 && x3 )
						nx_state = s34;
					else if( ~x69 && x70 && ~x63 && x10 && ~x64 && ~x44 && x11 && x36 && x34 && x4 && ~x5 && ~x3 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x69 && x70 && ~x63 && x10 && ~x64 && ~x44 && x11 && x36 && x34 && ~x4 && x3 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x70 && ~x63 && x10 && ~x64 && ~x44 && x11 && x36 && x34 && ~x4 && ~x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x69 && x70 && ~x63 && x10 && ~x64 && ~x44 && x11 && x36 && ~x34 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s513;
						end
					else if( ~x69 && x70 && ~x63 && x10 && ~x64 && ~x44 && x11 && ~x36 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && x70 && ~x63 && x10 && ~x64 && ~x44 && ~x11 && x12 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s513;
						end
					else if( ~x69 && x70 && ~x63 && x10 && ~x64 && ~x44 && ~x11 && ~x12 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s510;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && x64 && x40 && x34 && x8 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && x64 && x40 && x34 && ~x8 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s507;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && x64 && x40 && x34 && ~x8 && ~x5 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && x64 && x40 && ~x34 && x32 && x7 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && x64 && x40 && ~x34 && x32 && ~x7 && x45 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s507;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && x64 && x40 && ~x34 && x32 && ~x7 && x45 && ~x5 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && x64 && x40 && ~x34 && x32 && ~x7 && ~x45 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && x64 && x40 && ~x34 && ~x32 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && x64 && ~x40 && x1 )
						begin
							y16 = 1'b1;	y25 = 1'b1;	y27 = 1'b1;	
							nx_state = s514;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && x64 && ~x40 && ~x1 && x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && x64 && ~x40 && ~x1 && ~x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && ~x64 && x44 && x34 && x8 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && ~x64 && x44 && x34 && ~x8 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s511;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && ~x64 && x44 && x34 && ~x8 && ~x5 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && ~x64 && x44 && ~x34 && x32 && x7 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && ~x64 && x44 && ~x34 && x32 && ~x7 && x54 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s511;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && ~x64 && x44 && ~x34 && x32 && ~x7 && x54 && ~x5 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && ~x64 && x44 && ~x34 && x32 && ~x7 && ~x54 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s513;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && ~x64 && x44 && ~x34 && ~x32 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && ~x64 && ~x44 && x37 )
						begin
							y16 = 1'b1;	y25 = 1'b1;	y27 = 1'b1;	
							nx_state = s514;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && ~x64 && ~x44 && ~x37 && x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && x11 && ~x64 && ~x44 && ~x37 && ~x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && x12 && x64 && x40 && x20 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && x12 && x64 && x40 && ~x20 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && x12 && x64 && x40 && ~x20 && ~x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && x12 && x64 && ~x40 && x1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && x12 && x64 && ~x40 && ~x1 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && x12 && x64 && ~x40 && ~x1 && ~x4 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && x12 && ~x64 && x44 && x20 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s513;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && x12 && ~x64 && x44 && ~x20 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && x12 && ~x64 && x44 && ~x20 && ~x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && x12 && ~x64 && ~x44 && x37 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && x12 && ~x64 && ~x44 && ~x37 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && x12 && ~x64 && ~x44 && ~x37 && ~x4 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && ~x12 && x64 && x40 && x13 && x1 && x3 && x6 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s510;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && ~x12 && x64 && x40 && x13 && x1 && x3 && ~x6 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && ~x12 && x64 && x40 && x13 && x1 && ~x3 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && ~x12 && x64 && x40 && x13 && ~x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && ~x12 && x64 && x40 && ~x13 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && ~x12 && x64 && ~x40 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s449;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && ~x12 && x64 && ~x40 && ~x1 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && ~x12 && x64 && ~x40 && ~x1 && ~x2 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && ~x12 && x64 && ~x40 && ~x1 && ~x2 && ~x9 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && ~x12 && ~x64 && x44 && x13 && x37 && x41 && x6 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s510;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && ~x12 && ~x64 && x44 && x13 && x37 && x41 && ~x6 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && ~x12 && ~x64 && x44 && x13 && x37 && ~x41 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && ~x12 && ~x64 && x44 && x13 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s513;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && ~x12 && ~x64 && x44 && ~x13 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && ~x12 && ~x64 && ~x44 && x37 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s449;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && ~x12 && ~x64 && ~x44 && ~x37 && x34 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && ~x12 && ~x64 && ~x44 && ~x37 && ~x34 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && x70 && ~x63 && ~x10 && ~x11 && ~x12 && ~x64 && ~x44 && ~x37 && ~x34 && ~x9 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && ~x70 && x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							nx_state = s38;
						end
					else if( ~x69 && ~x70 && ~x3 && x7 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x3 && ~x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							nx_state = s38;
						end
					else nx_state = s34;
				s35 : if( x70 && x62 && x4 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( x70 && x62 && x4 && ~x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x70 && x62 && ~x4 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x70 && ~x62 && x63 && x9 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && x63 && ~x9 )
						nx_state = s35;
					else if( x70 && ~x62 && ~x63 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x70 && ~x62 && ~x63 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x70 && ~x62 && ~x63 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x65 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x4 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x24 && x26 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x65 && x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && ~x65 && x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && ~x65 && x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x24 && x25 && x26 )
						begin
							y11 = 1'b1;	y16 = 1'b1;	y25 = 1'b1;	
							nx_state = s515;
						end
					else if( ~x70 && ~x65 && ~x24 && x25 && ~x26 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && ~x65 && ~x24 && ~x25 && x26 && x3 && x16 && x11 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s122;
						end
					else if( ~x70 && ~x65 && ~x24 && ~x25 && x26 && x3 && x16 && ~x11 && x12 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s122;
						end
					else if( ~x70 && ~x65 && ~x24 && ~x25 && x26 && x3 && x16 && ~x11 && ~x12 && x10 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && ~x65 && ~x24 && ~x25 && x26 && x3 && x16 && ~x11 && ~x12 && ~x10 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s126;
						end
					else if( ~x70 && ~x65 && ~x24 && ~x25 && x26 && x3 && ~x16 && x17 && x10 && x12 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( ~x70 && ~x65 && ~x24 && ~x25 && x26 && x3 && ~x16 && x17 && x10 && ~x12 )
						begin
							y17 = 1'b1;	
							nx_state = s98;
						end
					else if( ~x70 && ~x65 && ~x24 && ~x25 && x26 && x3 && ~x16 && x17 && ~x10 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( ~x70 && ~x65 && ~x24 && ~x25 && x26 && x3 && ~x16 && ~x17 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s122;
						end
					else if( ~x70 && ~x65 && ~x24 && ~x25 && x26 && ~x3 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && ~x65 && ~x24 && ~x25 && ~x26 && x4 && x15 && x11 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( ~x70 && ~x65 && ~x24 && ~x25 && ~x26 && x4 && x15 && ~x11 && x12 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( ~x70 && ~x65 && ~x24 && ~x25 && ~x26 && x4 && x15 && ~x11 && ~x12 && x10 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && ~x65 && ~x24 && ~x25 && ~x26 && x4 && x15 && ~x11 && ~x12 && ~x10 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s126;
						end
					else if( ~x70 && ~x65 && ~x24 && ~x25 && ~x26 && x4 && ~x15 && x16 && x10 && x12 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x70 && ~x65 && ~x24 && ~x25 && ~x26 && x4 && ~x15 && x16 && x10 && ~x12 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s370;
						end
					else if( ~x70 && ~x65 && ~x24 && ~x25 && ~x26 && x4 && ~x15 && x16 && ~x10 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x70 && ~x65 && ~x24 && ~x25 && ~x26 && x4 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( ~x70 && ~x65 && ~x24 && ~x25 && ~x26 && ~x4 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s304;
						end
					else nx_state = s35;
				s36 : if( x69 && x65 && x70 && x62 && x64 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && x65 && x70 && x62 && ~x64 && x66 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && x65 && x70 && x62 && ~x64 && x66 && ~x6 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x65 && x70 && x62 && ~x64 && ~x66 && x67 )
						nx_state = s1;
					else if( x69 && x65 && x70 && x62 && ~x64 && ~x66 && ~x67 && x4 && x5 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s18;
						end
					else if( x69 && x65 && x70 && x62 && ~x64 && ~x66 && ~x67 && x4 && x5 && ~x1 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( x69 && x65 && x70 && x62 && ~x64 && ~x66 && ~x67 && x4 && ~x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x65 && x70 && x62 && ~x64 && ~x66 && ~x67 && ~x4 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( x69 && x65 && x70 && ~x62 && x63 && x66 && x7 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x69 && x65 && x70 && ~x62 && x63 && x66 && ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && x70 && ~x62 && x63 && ~x66 && x67 && x15 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	
							nx_state = s231;
						end
					else if( x69 && x65 && x70 && ~x62 && x63 && ~x66 && x67 && ~x15 )
						nx_state = s1;
					else if( x69 && x65 && x70 && ~x62 && x63 && ~x66 && ~x67 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && x67 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && x22 && x21 && x10 && x14 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && x22 && x21 && x10 && ~x14 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && x22 && x21 && ~x10 && x11 && x14 && x8 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && x22 && x21 && ~x10 && x11 && x14 && ~x8 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && x22 && x21 && ~x10 && x11 && x14 && ~x8 && x6 && ~x7 )
						nx_state = s1;
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && x22 && x21 && ~x10 && x11 && x14 && ~x8 && ~x6 )
						nx_state = s1;
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && x22 && x21 && ~x10 && x11 && ~x14 && x7 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && x22 && x21 && ~x10 && x11 && ~x14 && ~x7 && x6 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && x22 && x21 && ~x10 && x11 && ~x14 && ~x7 && x6 && ~x8 )
						nx_state = s1;
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && x22 && x21 && ~x10 && x11 && ~x14 && ~x7 && ~x6 )
						nx_state = s1;
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && x22 && x21 && ~x10 && ~x11 && x14 )
						begin
							y60 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y67 = 1'b1;	y68 = 1'b1;	
							nx_state = s516;
						end
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && x22 && x21 && ~x10 && ~x11 && ~x14 )
						begin
							y58 = 1'b1;	y59 = 1'b1;	y60 = 1'b1;	
							y62 = 1'b1;	
							nx_state = s516;
						end
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && x22 && ~x21 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && x22 && ~x21 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && x22 && ~x21 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && x22 && ~x21 && ~x6 )
						nx_state = s1;
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && ~x22 && x12 && x21 && x11 )
						begin
							y7 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y93 = 1'b1;	
							nx_state = s516;
						end
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && ~x22 && x12 && x21 && ~x11 )
						begin
							y7 = 1'b1;	y62 = 1'b1;	y74 = 1'b1;	
							y110 = 1'b1;	
							nx_state = s517;
						end
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && ~x22 && x12 && ~x21 && x10 )
						begin
							y7 = 1'b1;	y62 = 1'b1;	y90 = 1'b1;	
							y92 = 1'b1;	
							nx_state = s516;
						end
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && ~x22 && x12 && ~x21 && ~x10 )
						begin
							y7 = 1'b1;	y62 = 1'b1;	y92 = 1'b1;	
							y93 = 1'b1;	y97 = 1'b1;	
							nx_state = s516;
						end
					else if( x69 && x65 && x70 && ~x62 && ~x63 && x64 && ~x67 && ~x22 && ~x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y62 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s518;
						end
					else if( x69 && x65 && x70 && ~x62 && ~x63 && ~x64 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x65 && ~x70 && x21 && x18 && x20 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x65 && ~x70 && x21 && x18 && ~x20 )
						nx_state = s36;
					else if( x69 && x65 && ~x70 && x21 && ~x18 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && x65 && ~x70 && ~x21 && x22 && x15 && x9 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && x65 && ~x70 && ~x21 && x22 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && x65 && ~x70 && ~x21 && x22 && ~x15 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s495;
						end
					else if( x69 && x65 && ~x70 && ~x21 && ~x22 && x23 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && x65 && ~x70 && ~x21 && ~x22 && x23 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && x65 && ~x70 && ~x21 && ~x22 && x23 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && x65 && ~x70 && ~x21 && ~x22 && x23 && ~x20 )
						nx_state = s1;
					else if( x69 && x65 && ~x70 && ~x21 && ~x22 && ~x23 && x18 && x14 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && x65 && ~x70 && ~x21 && ~x22 && ~x23 && x18 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && x65 && ~x70 && ~x21 && ~x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && x65 && ~x70 && ~x21 && ~x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && x62 && x64 && x12 && x9 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x65 && x70 && x62 && x64 && x12 && ~x9 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x69 && ~x65 && x70 && x62 && x64 && x12 && ~x9 && ~x3 && x1 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x65 && x70 && x62 && x64 && x12 && ~x9 && ~x3 && ~x1 && x7 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	
							nx_state = s474;
						end
					else if( x69 && ~x65 && x70 && x62 && x64 && x12 && ~x9 && ~x3 && ~x1 && ~x7 )
						nx_state = s36;
					else if( x69 && ~x65 && x70 && x62 && x64 && ~x12 && x10 && x13 && x11 && x4 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s476;
						end
					else if( x69 && ~x65 && x70 && x62 && x64 && ~x12 && x10 && x13 && x11 && ~x4 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x65 && x70 && x62 && x64 && ~x12 && x10 && x13 && ~x11 && x14 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s27;
						end
					else if( x69 && ~x65 && x70 && x62 && x64 && ~x12 && x10 && x13 && ~x11 && ~x14 && x9 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x65 && x70 && x62 && x64 && ~x12 && x10 && x13 && ~x11 && ~x14 && ~x9 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x69 && ~x65 && x70 && x62 && x64 && ~x12 && x10 && x13 && ~x11 && ~x14 && ~x9 && ~x3 && x1 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x65 && x70 && x62 && x64 && ~x12 && x10 && x13 && ~x11 && ~x14 && ~x9 && ~x3 && ~x1 && x7 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	
							nx_state = s474;
						end
					else if( x69 && ~x65 && x70 && x62 && x64 && ~x12 && x10 && x13 && ~x11 && ~x14 && ~x9 && ~x3 && ~x1 && ~x7 )
						nx_state = s36;
					else if( x69 && ~x65 && x70 && x62 && x64 && ~x12 && x10 && ~x13 && x9 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x65 && x70 && x62 && x64 && ~x12 && x10 && ~x13 && ~x9 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x69 && ~x65 && x70 && x62 && x64 && ~x12 && x10 && ~x13 && ~x9 && ~x3 && x1 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x65 && x70 && x62 && x64 && ~x12 && x10 && ~x13 && ~x9 && ~x3 && ~x1 && x7 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	
							nx_state = s474;
						end
					else if( x69 && ~x65 && x70 && x62 && x64 && ~x12 && x10 && ~x13 && ~x9 && ~x3 && ~x1 && ~x7 )
						nx_state = s36;
					else if( x69 && ~x65 && x70 && x62 && x64 && ~x12 && ~x10 && x9 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x65 && x70 && x62 && x64 && ~x12 && ~x10 && ~x9 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x69 && ~x65 && x70 && x62 && x64 && ~x12 && ~x10 && ~x9 && ~x3 && x1 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x65 && x70 && x62 && x64 && ~x12 && ~x10 && ~x9 && ~x3 && ~x1 && x7 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	
							nx_state = s474;
						end
					else if( x69 && ~x65 && x70 && x62 && x64 && ~x12 && ~x10 && ~x9 && ~x3 && ~x1 && ~x7 )
						nx_state = s36;
					else if( x69 && ~x65 && x70 && x62 && ~x64 && x66 && x1 && x2 && x3 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x69 && ~x65 && x70 && x62 && ~x64 && x66 && x1 && x2 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x69 && ~x65 && x70 && x62 && ~x64 && x66 && x1 && ~x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x69 && ~x65 && x70 && x62 && ~x64 && x66 && ~x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x65 && x70 && x62 && ~x64 && ~x66 && x17 && x18 && x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	
							nx_state = s20;
						end
					else if( x69 && ~x65 && x70 && x62 && ~x64 && ~x66 && x17 && x18 && ~x1 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x65 && x70 && x62 && ~x64 && ~x66 && x17 && x18 && ~x1 && ~x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && ~x65 && x70 && x62 && ~x64 && ~x66 && x17 && ~x18 && x7 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x65 && x70 && x62 && ~x64 && ~x66 && x17 && ~x18 && ~x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x65 && x70 && x62 && ~x64 && ~x66 && ~x17 && x18 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x65 && x70 && x62 && ~x64 && ~x66 && ~x17 && x18 && ~x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( x69 && ~x65 && x70 && x62 && ~x64 && ~x66 && ~x17 && ~x18 && x19 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && x62 && ~x64 && ~x66 && ~x17 && ~x18 && ~x19 && x1 && x2 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x65 && x70 && x62 && ~x64 && ~x66 && ~x17 && ~x18 && ~x19 && x1 && ~x2 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && x62 && ~x64 && ~x66 && ~x17 && ~x18 && ~x19 && ~x1 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && x66 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && x66 && ~x8 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s35;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && x22 && x16 && x23 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s442;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && x22 && x16 && ~x23 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && x22 && x16 && ~x23 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && x22 && x16 && ~x23 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && x22 && x16 && ~x23 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && x22 && x16 && ~x23 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && x22 && ~x16 && x23 )
						begin
							y3 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s520;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && x22 && ~x16 && ~x23 )
						begin
							y3 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s521;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && x9 && x8 && x10 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y5 = 1'b1;	
							y22 = 1'b1;	y23 = 1'b1;	
							nx_state = s72;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && x9 && x8 && ~x10 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && x9 && ~x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && x10 && x8 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && x10 && x8 && ~x13 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && x10 && x8 && ~x13 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && x10 && x8 && ~x13 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && x10 && x8 && ~x13 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && x10 && x8 && ~x13 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && x10 && ~x8 && x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && x10 && ~x8 && ~x3 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && x10 && ~x8 && ~x3 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && x10 && ~x8 && ~x3 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && x10 && ~x8 && ~x3 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && x10 && ~x8 && ~x3 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && ~x10 && x8 && x1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && ~x10 && x8 && ~x1 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && ~x10 && x8 && ~x1 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && ~x10 && x8 && ~x1 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && ~x10 && x8 && ~x1 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && ~x10 && x8 && ~x1 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && ~x10 && ~x8 && x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && ~x10 && ~x8 && ~x15 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && ~x10 && ~x8 && ~x15 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && ~x10 && ~x8 && ~x15 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && ~x10 && ~x8 && ~x15 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && x7 && ~x9 && ~x10 && ~x8 && ~x15 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && x23 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s523;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && x16 && ~x23 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s442;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && ~x16 && x23 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s524;
						end
					else if( x69 && ~x65 && x70 && ~x62 && x63 && ~x66 && ~x22 && ~x16 && ~x23 )
						begin
							y3 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s520;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && x4 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && x5 && x18 && x19 && x12 )
						begin
							y54 = 1'b1;	
							nx_state = s525;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && x5 && x18 && x19 && ~x12 )
						begin
							y55 = 1'b1;	
							nx_state = s526;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && x5 && x18 && ~x19 && x12 && x6 )
						begin
							y16 = 1'b1;	y50 = 1'b1;	
							nx_state = s527;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && x5 && x18 && ~x19 && x12 && ~x6 && x16 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && x5 && x18 && ~x19 && x12 && ~x6 && ~x16 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && x5 && x18 && ~x19 && x12 && ~x6 && ~x16 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && x5 && x18 && ~x19 && x12 && ~x6 && ~x16 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && x5 && x18 && ~x19 && x12 && ~x6 && ~x16 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && x5 && x18 && ~x19 && ~x12 && x6 )
						begin
							y12 = 1'b1;	y48 = 1'b1;	
							nx_state = s529;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && x5 && x18 && ~x19 && ~x12 && ~x6 && x15 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && x5 && x18 && ~x19 && ~x12 && ~x6 && ~x15 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && x5 && x18 && ~x19 && ~x12 && ~x6 && ~x15 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && x5 && x18 && ~x19 && ~x12 && ~x6 && ~x15 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && x5 && x18 && ~x19 && ~x12 && ~x6 && ~x15 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && x5 && ~x18 && x19 )
						begin
							y27 = 1'b1;	y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s284;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && x5 && ~x18 && ~x19 && x6 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && x5 && ~x18 && ~x19 && ~x6 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && x19 && x6 && x12 && x11 )
						begin
							y46 = 1'b1;	
							nx_state = s531;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && x19 && x6 && x12 && ~x11 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && x19 && x6 && x12 && ~x11 && x9 && ~x10 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && x19 && x6 && x12 && ~x11 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && x19 && x6 && ~x12 && x10 )
						begin
							y46 = 1'b1;	
							nx_state = s531;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && x19 && x6 && ~x12 && ~x10 && x9 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && x19 && x6 && ~x12 && ~x10 && x9 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && x19 && x6 && ~x12 && ~x10 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && x19 && ~x6 && x12 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && x19 && ~x6 && ~x12 )
						begin
							y56 = 1'b1;	y57 = 1'b1;	
							nx_state = s284;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && ~x19 && x6 && x12 && x14 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && ~x19 && x6 && x12 && ~x14 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && ~x19 && x6 && x12 && ~x14 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && ~x19 && x6 && x12 && ~x14 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && ~x19 && x6 && x12 && ~x14 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && ~x19 && x6 && ~x12 && x13 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && ~x19 && x6 && ~x12 && ~x13 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && ~x19 && x6 && ~x12 && ~x13 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && ~x19 && x6 && ~x12 && ~x13 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && ~x19 && x6 && ~x12 && ~x13 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && x18 && ~x19 && ~x6 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && ~x18 && x19 && x12 && x6 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && ~x18 && x19 && x12 && ~x6 )
						begin
							y38 = 1'b1;	
							nx_state = s532;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && ~x18 && x19 && ~x12 && x6 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && ~x18 && x19 && ~x12 && ~x6 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && x8 && ~x5 && ~x18 && ~x19 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && x64 && ~x4 && ~x8 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && ~x64 && x21 && x22 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && ~x64 && x21 && ~x22 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && ~x64 && x21 && ~x22 && ~x23 )
						nx_state = s1;
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && ~x64 && ~x21 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( x69 && ~x65 && x70 && ~x62 && ~x63 && ~x64 && ~x21 && ~x23 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && x68 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && x68 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && x68 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && x68 && x21 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && x68 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && x68 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && x68 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && x68 && ~x21 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && x14 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && x14 && ~x8 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && ~x14 && x7 && x8 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s296;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && ~x14 && x7 && ~x8 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s297;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && ~x14 && ~x7 && x8 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && x17 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && x17 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && ~x14 && ~x7 && ~x8 && x13 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && x17 && x12 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && x17 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && x2 && x8 && x7 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && x2 && x8 && ~x7 && x9 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && x2 && x8 && ~x7 && ~x9 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && x2 && ~x8 && x7 && x11 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && x2 && ~x8 && x7 && ~x11 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && x2 && ~x8 && ~x7 && x10 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && x2 && ~x8 && ~x7 && ~x10 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && x7 && x8 && x1 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && x7 && x8 && ~x1 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && x7 && ~x8 && x11 && x1 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && x7 && ~x8 && x11 && ~x1 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && x7 && ~x8 && ~x11 && x17 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && x7 && ~x8 && ~x11 && x17 && ~x13 && x12 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && x7 && ~x8 && ~x11 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && x7 && ~x8 && ~x11 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && x8 && x9 && x1 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && x8 && x9 && ~x1 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && x8 && ~x9 && x17 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && x8 && ~x9 && x17 && ~x13 && x12 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && x8 && ~x9 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && x8 && ~x9 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && ~x8 && x10 && x1 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && ~x8 && x10 && ~x1 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && ~x8 && ~x10 && x17 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && ~x8 && ~x10 && x17 && ~x13 && x12 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && ~x8 && ~x10 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && ~x8 && ~x10 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && ~x16 && x15 && x7 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s298;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && ~x16 && x15 && ~x7 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && ~x16 && x15 && ~x7 && ~x2 && x1 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && ~x16 && x15 && ~x7 && ~x2 && ~x1 && x8 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && ~x16 && x15 && ~x7 && ~x2 && ~x1 && ~x8 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && ~x16 && ~x15 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && ~x16 && ~x15 && ~x2 && x1 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && x64 && ~x16 && ~x15 && ~x2 && ~x1 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y28 = 1'b1;	
							nx_state = s299;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && x63 && ~x64 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && x16 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && x16 && ~x8 && x6 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && x16 && ~x8 && ~x6 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && x8 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && x8 && ~x7 && x9 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && x8 && ~x7 && ~x9 && x19 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && x8 && ~x7 && ~x9 && x19 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && x8 && ~x7 && ~x9 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && x8 && ~x7 && ~x9 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && ~x8 && x7 && x11 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && ~x8 && x7 && ~x11 && x19 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && ~x8 && x7 && ~x11 && x19 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && ~x8 && x7 && ~x11 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && ~x8 && x7 && ~x11 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && ~x8 && ~x7 && x10 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && ~x8 && ~x7 && ~x10 && x19 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && ~x8 && ~x7 && ~x10 && x19 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && ~x8 && ~x7 && ~x10 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && ~x8 && ~x7 && ~x10 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && ~x4 && x6 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y28 = 1'b1;	
							nx_state = s299;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && ~x4 && ~x6 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && ~x64 && x19 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && ~x64 && x19 && ~x13 && x12 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && ~x64 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && x66 && ~x68 && ~x63 && ~x64 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && x24 && x26 && x16 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && x24 && x26 && ~x16 && x17 && x13 && x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && x24 && x26 && ~x16 && x17 && x13 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s497;
						end
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && x24 && x26 && ~x16 && x17 && x13 && ~x11 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && x24 && x26 && ~x16 && x17 && ~x13 && x11 )
						begin
							y17 = 1'b1;	
							nx_state = s98;
						end
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && x24 && x26 && ~x16 && x17 && ~x13 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && x24 && x26 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s35;
						end
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && x24 && ~x26 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && ~x24 && x25 && x26 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && ~x24 && x25 && x26 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && ~x24 && x25 && x26 && x19 && ~x14 && ~x13 )
						nx_state = s36;
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && ~x24 && x25 && x26 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && ~x24 && x25 && ~x26 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && ~x24 && ~x25 && x26 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && ~x24 && ~x25 && ~x26 && x15 && x12 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && ~x24 && ~x25 && ~x26 && x15 && ~x12 && x11 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && ~x24 && ~x25 && ~x26 && x15 && ~x12 && ~x11 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && ~x24 && ~x25 && ~x26 && x15 && ~x12 && ~x11 && ~x10 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && ~x24 && ~x25 && ~x26 && ~x15 && x16 && x10 && x12 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s122;
						end
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && ~x24 && ~x25 && ~x26 && ~x15 && x16 && x10 && ~x12 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && ~x24 && ~x25 && ~x26 && ~x15 && x16 && ~x10 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s122;
						end
					else if( x69 && ~x65 && ~x70 && x67 && ~x66 && ~x24 && ~x25 && ~x26 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x65 && ~x70 && ~x67 && x66 && x21 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && ~x67 && x66 && ~x21 && x22 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x69 && ~x65 && ~x70 && ~x67 && x66 && ~x21 && x22 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x69 && ~x65 && ~x70 && ~x67 && x66 && ~x21 && x22 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && ~x67 && x66 && ~x21 && x22 && ~x7 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && ~x67 && x66 && ~x21 && ~x22 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x65 && ~x70 && ~x67 && x66 && ~x21 && ~x22 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x65 && ~x70 && ~x67 && x66 && ~x21 && ~x22 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && ~x67 && ~x66 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x69 && ~x65 && ~x70 && ~x67 && ~x66 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x69 && ~x65 && ~x70 && ~x67 && ~x66 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x70 && ~x67 && ~x66 && ~x3 )
						nx_state = s1;
					else if( ~x69 && x45 && x44 && x31 && x19 && x10 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s387;
						end
					else if( ~x69 && x45 && x44 && x31 && x19 && ~x10 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x69 && x45 && x44 && x31 && ~x19 )
						nx_state = s36;
					else if( ~x69 && x45 && x44 && ~x31 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x69 && x45 && ~x44 && x46 && x47 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && x45 && ~x44 && x46 && ~x47 && x10 && x6 && x2 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s387;
						end
					else if( ~x69 && x45 && ~x44 && x46 && ~x47 && x10 && x6 && ~x2 )
						nx_state = s36;
					else if( ~x69 && x45 && ~x44 && x46 && ~x47 && x10 && ~x6 && x2 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x69 && x45 && ~x44 && x46 && ~x47 && x10 && ~x6 && ~x2 )
						nx_state = s36;
					else if( ~x69 && x45 && ~x44 && x46 && ~x47 && ~x10 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x69 && x45 && ~x44 && ~x46 && x12 && x9 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && x45 && ~x44 && ~x46 && x12 && ~x9 && x7 )
						nx_state = s1;
					else if( ~x69 && x45 && ~x44 && ~x46 && x12 && ~x9 && ~x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( ~x69 && x45 && ~x44 && ~x46 && ~x12 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && ~x45 && x44 && x46 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x69 && ~x45 && x44 && ~x46 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && ~x45 && ~x44 && x46 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && ~x45 && ~x44 && ~x46 && x11 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && ~x45 && ~x44 && ~x46 && ~x11 && x9 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && ~x45 && ~x44 && ~x46 && ~x11 && ~x9 && x7 )
						nx_state = s1;
					else if( ~x69 && ~x45 && ~x44 && ~x46 && ~x11 && ~x9 && ~x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else nx_state = s36;
				s37 : if( x1 && x2 && x3 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x1 && x2 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x1 && ~x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else nx_state = s37;
				s38 : if( x69 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s534;
						end
					else if( ~x69 && x3 && x4 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && x3 && ~x4 )
						nx_state = s38;
					else if( ~x69 && ~x3 )
						nx_state = s1;
					else nx_state = s38;
				s39 : if( x62 && x65 && x20 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y20 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s535;
						end
					else if( x62 && x65 && ~x20 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s536;
						end
					else if( x62 && ~x65 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s537;
						end
					else if( ~x62 && x21 && x20 )
						begin
							y28 = 1'b1;	
							nx_state = s539;
						end
					else if( ~x62 && x21 && ~x20 )
						begin
							y7 = 1'b1;	y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s538;
						end
					else if( ~x62 && ~x21 )
						begin
							y28 = 1'b1;	
							nx_state = s539;
						end
					else nx_state = s39;
				s40 : if( x69 && x62 && x13 && x10 && x3 && x5 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( x69 && x62 && x13 && x10 && x3 && ~x5 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && x62 && x13 && x10 && ~x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && x62 && x13 && ~x10 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && x62 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && x62 && ~x13 && ~x12 && x10 && x5 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && x62 && ~x13 && ~x12 && x10 && ~x5 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && x62 && ~x13 && ~x12 && ~x10 && x5 && x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s540;
						end
					else if( x69 && x62 && ~x13 && ~x12 && ~x10 && x5 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x69 && x62 && ~x13 && ~x12 && ~x10 && x5 && ~x3 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && x62 && ~x13 && ~x12 && ~x10 && ~x5 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && ~x62 && x17 && x18 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x1 && x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x1 && ~x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && ~x62 && x17 && ~x18 && x7 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s541;
						end
					else if( x69 && ~x62 && x17 && ~x18 && ~x7 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s542;
						end
					else if( x69 && ~x62 && ~x17 && x15 && x18 && x5 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && ~x62 && ~x17 && x15 && x18 && ~x5 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && ~x62 && ~x17 && x15 && ~x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && ~x62 && ~x17 && ~x15 && x5 && x18 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && ~x62 && ~x17 && ~x15 && x5 && ~x18 && x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && ~x62 && ~x17 && ~x15 && x5 && ~x18 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x69 && ~x62 && ~x17 && ~x15 && x5 && ~x18 && ~x3 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && ~x62 && ~x17 && ~x15 && ~x5 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x69 && x18 && x17 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( ~x69 && x18 && x17 && ~x1 && x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x18 && x17 && ~x1 && ~x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x69 && x18 && ~x17 && x19 && x5 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x18 && ~x17 && x19 && ~x5 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s543;
						end
					else if( ~x69 && x18 && ~x17 && ~x19 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x69 && ~x18 && x17 && x7 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s541;
						end
					else if( ~x69 && ~x18 && x17 && ~x7 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s542;
						end
					else if( ~x69 && ~x18 && ~x17 && x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( ~x69 && ~x18 && ~x17 && ~x19 && x5 && x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x69 && ~x18 && ~x17 && ~x19 && x5 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && ~x18 && ~x17 && ~x19 && x5 && ~x3 && ~x4 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s543;
						end
					else if( ~x69 && ~x18 && ~x17 && ~x19 && ~x5 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else nx_state = s40;
				s41 : if( x69 && x62 && x13 && x10 && x17 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x69 && x62 && x13 && x10 && ~x17 && x15 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && x62 && x13 && x10 && ~x17 && ~x15 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && x62 && x13 && ~x10 && x3 && x15 )
						nx_state = s41;
					else if( x69 && x62 && x13 && ~x10 && x3 && ~x15 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && x62 && x13 && ~x10 && ~x3 && x4 && x5 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && x62 && x13 && ~x10 && ~x3 && x4 && ~x5 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && x62 && x13 && ~x10 && ~x3 && ~x4 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && x62 && ~x13 && x12 && x4 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && x62 && ~x13 && x12 && ~x4 )
						nx_state = s1;
					else if( x69 && x62 && ~x13 && ~x12 && x10 && x11 )
						nx_state = s1;
					else if( x69 && x62 && ~x13 && ~x12 && x10 && ~x11 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s544;
						end
					else if( x69 && x62 && ~x13 && ~x12 && ~x10 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && x17 && x18 && x6 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s540;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x6 && x8 && x4 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x6 && x8 && ~x4 && x1 && x3 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x6 && x8 && ~x4 && x1 && ~x3 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x6 && x8 && ~x4 && ~x1 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x6 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x62 && x17 && ~x18 && x12 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s45;
						end
					else if( x69 && ~x62 && x17 && ~x18 && ~x12 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && ~x62 && ~x17 && x15 && x18 && x9 )
						nx_state = s1;
					else if( x69 && ~x62 && ~x17 && x15 && x18 && ~x9 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s544;
						end
					else if( x69 && ~x62 && ~x17 && x15 && ~x18 && x2 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && ~x17 && x15 && ~x18 && ~x2 )
						nx_state = s1;
					else if( x69 && ~x62 && ~x17 && ~x15 && x18 && x4 && x5 && x3 )
						nx_state = s41;
					else if( x69 && ~x62 && ~x17 && ~x15 && x18 && x4 && x5 && ~x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && ~x17 && ~x15 && x18 && x4 && ~x5 && x3 )
						nx_state = s41;
					else if( x69 && ~x62 && ~x17 && ~x15 && x18 && x4 && ~x5 && ~x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && ~x62 && ~x17 && ~x15 && x18 && ~x4 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && ~x62 && ~x17 && ~x15 && x18 && ~x4 && ~x3 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && ~x62 && ~x17 && ~x15 && ~x18 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x63 && x11 && x43 && x41 && x13 && x3 && x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s99;
						end
					else if( ~x69 && x63 && x11 && x43 && x41 && x13 && x3 && ~x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x63 && x11 && x43 && x41 && x13 && ~x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x63 && x11 && x43 && x41 && ~x13 && x5 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s181;
						end
					else if( ~x69 && x63 && x11 && x43 && x41 && ~x13 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x63 && x11 && x43 && ~x41 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x69 && x63 && x11 && ~x43 && x44 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x69 && x63 && x11 && ~x43 && ~x44 && x10 && x45 && x5 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s183;
						end
					else if( ~x69 && x63 && x11 && ~x43 && ~x44 && x10 && x45 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x63 && x11 && ~x43 && ~x44 && x10 && ~x45 && x32 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s181;
						end
					else if( ~x69 && x63 && x11 && ~x43 && ~x44 && x10 && ~x45 && ~x32 && x3 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x63 && x11 && ~x43 && ~x44 && x10 && ~x45 && ~x32 && x3 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x69 && x63 && x11 && ~x43 && ~x44 && x10 && ~x45 && ~x32 && x3 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x69 && x63 && x11 && ~x43 && ~x44 && x10 && ~x45 && ~x32 && x3 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x63 && x11 && ~x43 && ~x44 && x10 && ~x45 && ~x32 && x3 && x15 && ~x47 && ~x1 )
						nx_state = s41;
					else if( ~x69 && x63 && x11 && ~x43 && ~x44 && x10 && ~x45 && ~x32 && x3 && ~x15 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x63 && x11 && ~x43 && ~x44 && x10 && ~x45 && ~x32 && ~x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x63 && x11 && ~x43 && ~x44 && ~x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x69 && x63 && ~x11 && x41 && x12 && x5 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s183;
						end
					else if( ~x69 && x63 && ~x11 && x41 && x12 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x63 && ~x11 && x41 && ~x12 && x13 && x45 && x36 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x63 && ~x11 && x41 && ~x12 && x13 && x45 && ~x36 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x63 && ~x11 && x41 && ~x12 && x13 && ~x45 && x39 && x1 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s183;
						end
					else if( ~x69 && x63 && ~x11 && x41 && ~x12 && x13 && ~x45 && x39 && ~x1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x63 && ~x11 && x41 && ~x12 && x13 && ~x45 && ~x39 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s183;
						end
					else if( ~x69 && x63 && ~x11 && x41 && ~x12 && ~x13 && x45 && x5 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s183;
						end
					else if( ~x69 && x63 && ~x11 && x41 && ~x12 && ~x13 && x45 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x63 && ~x11 && x41 && ~x12 && ~x13 && ~x45 && x32 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s181;
						end
					else if( ~x69 && x63 && ~x11 && x41 && ~x12 && ~x13 && ~x45 && ~x32 && x3 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x63 && ~x11 && x41 && ~x12 && ~x13 && ~x45 && ~x32 && x3 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x69 && x63 && ~x11 && x41 && ~x12 && ~x13 && ~x45 && ~x32 && x3 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x69 && x63 && ~x11 && x41 && ~x12 && ~x13 && ~x45 && ~x32 && x3 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x63 && ~x11 && x41 && ~x12 && ~x13 && ~x45 && ~x32 && x3 && x15 && ~x47 && ~x1 )
						nx_state = s41;
					else if( ~x69 && x63 && ~x11 && x41 && ~x12 && ~x13 && ~x45 && ~x32 && x3 && ~x15 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x63 && ~x11 && x41 && ~x12 && ~x13 && ~x45 && ~x32 && ~x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x63 && ~x11 && ~x41 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x69 && ~x63 && x18 && x17 && x6 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s546;
						end
					else if( ~x69 && ~x63 && x18 && x17 && ~x6 && x8 && x4 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( ~x69 && ~x63 && x18 && x17 && ~x6 && x8 && ~x4 && x40 && x31 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && ~x63 && x18 && x17 && ~x6 && x8 && ~x4 && x40 && ~x31 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x69 && ~x63 && x18 && x17 && ~x6 && x8 && ~x4 && ~x40 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s543;
						end
					else if( ~x69 && ~x63 && x18 && x17 && ~x6 && ~x8 && x15 && x16 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x69 && ~x63 && x18 && x17 && ~x6 && ~x8 && x15 && x16 && ~x5 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x69 && ~x63 && x18 && x17 && ~x6 && ~x8 && x15 && ~x16 && x1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x63 && x18 && x17 && ~x6 && ~x8 && x15 && ~x16 && ~x1 )
						nx_state = s41;
					else if( ~x69 && ~x63 && x18 && x17 && ~x6 && ~x8 && ~x15 && x16 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x63 && x18 && x17 && ~x6 && ~x8 && ~x15 && ~x16 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x69 && ~x63 && x18 && x17 && ~x6 && ~x8 && ~x15 && ~x16 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x63 && x18 && ~x17 && x19 && x9 && x15 && x16 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x69 && ~x63 && x18 && ~x17 && x19 && x9 && x15 && x16 && ~x5 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x69 && ~x63 && x18 && ~x17 && x19 && x9 && x15 && x16 && ~x5 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x69 && ~x63 && x18 && ~x17 && x19 && x9 && x15 && ~x16 && x1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x63 && x18 && ~x17 && x19 && x9 && x15 && ~x16 && ~x1 )
						nx_state = s41;
					else if( ~x69 && ~x63 && x18 && ~x17 && x19 && x9 && ~x15 && x16 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x63 && x18 && ~x17 && x19 && x9 && ~x15 && ~x16 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x69 && ~x63 && x18 && ~x17 && x19 && x9 && ~x15 && ~x16 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x63 && x18 && ~x17 && x19 && ~x9 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s544;
						end
					else if( ~x69 && ~x63 && x18 && ~x17 && ~x19 && x4 && x5 && x3 )
						nx_state = s41;
					else if( ~x69 && ~x63 && x18 && ~x17 && ~x19 && x4 && x5 && ~x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && ~x63 && x18 && ~x17 && ~x19 && x4 && ~x5 && x3 )
						nx_state = s41;
					else if( ~x69 && ~x63 && x18 && ~x17 && ~x19 && x4 && ~x5 && ~x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x69 && ~x63 && x18 && ~x17 && ~x19 && ~x4 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( ~x69 && ~x63 && x18 && ~x17 && ~x19 && ~x4 && ~x3 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( ~x69 && ~x63 && ~x18 && x17 && x12 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s45;
						end
					else if( ~x69 && ~x63 && ~x18 && x17 && ~x12 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( ~x69 && ~x63 && ~x18 && ~x17 && x19 && x35 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && ~x63 && ~x18 && ~x17 && x19 && ~x35 && x15 && x16 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x69 && ~x63 && ~x18 && ~x17 && x19 && ~x35 && x15 && x16 && ~x5 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x69 && ~x63 && ~x18 && ~x17 && x19 && ~x35 && x15 && x16 && ~x5 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x69 && ~x63 && ~x18 && ~x17 && x19 && ~x35 && x15 && ~x16 && x1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x63 && ~x18 && ~x17 && x19 && ~x35 && x15 && ~x16 && ~x1 )
						nx_state = s41;
					else if( ~x69 && ~x63 && ~x18 && ~x17 && x19 && ~x35 && ~x15 && x16 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x63 && ~x18 && ~x17 && x19 && ~x35 && ~x15 && ~x16 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x69 && ~x63 && ~x18 && ~x17 && x19 && ~x35 && ~x15 && ~x16 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x63 && ~x18 && ~x17 && ~x19 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else nx_state = s41;
				s42 : if( x69 && x62 && x13 && x10 && x9 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && x62 && x13 && x10 && ~x9 && x17 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && x62 && x13 && x10 && ~x9 && ~x17 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && x62 && x13 && ~x10 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && x62 && ~x13 && x12 && x4 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && x62 && ~x13 && x12 && ~x4 )
						nx_state = s1;
					else if( x69 && x62 && ~x13 && ~x12 && x10 && x2 && x16 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( x69 && x62 && ~x13 && ~x12 && x10 && x2 && ~x16 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && x62 && ~x13 && ~x12 && x10 && ~x2 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && x62 && ~x13 && ~x12 && ~x10 && x18 && x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s540;
						end
					else if( x69 && x62 && ~x13 && ~x12 && ~x10 && x18 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x69 && x62 && ~x13 && ~x12 && ~x10 && x18 && ~x3 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && x62 && ~x13 && ~x12 && ~x10 && ~x18 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && x17 && x18 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x1 && x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x1 && ~x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && ~x62 && x17 && ~x18 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && ~x62 && ~x17 && x15 && x18 && x2 && x4 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( x69 && ~x62 && ~x17 && x15 && x18 && x2 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && ~x62 && ~x17 && x15 && x18 && ~x2 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && ~x17 && x15 && ~x18 && x2 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && ~x17 && x15 && ~x18 && ~x2 )
						nx_state = s1;
					else if( x69 && ~x62 && ~x17 && ~x15 && x1 && x18 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && ~x17 && ~x15 && x1 && ~x18 && x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && ~x62 && ~x17 && ~x15 && x1 && ~x18 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x69 && ~x62 && ~x17 && ~x15 && x1 && ~x18 && ~x3 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && ~x62 && ~x17 && ~x15 && ~x1 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x17 && x18 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( ~x69 && x17 && x18 && ~x1 && x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x17 && x18 && ~x1 && ~x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x69 && x17 && ~x18 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && ~x17 && x19 && x18 && x39 && x4 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x69 && ~x17 && x19 && x18 && x39 && ~x4 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s543;
						end
					else if( ~x69 && ~x17 && x19 && x18 && ~x39 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && ~x17 && x19 && ~x18 && x35 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && ~x17 && x19 && ~x18 && ~x35 && x15 && x16 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x69 && ~x17 && x19 && ~x18 && ~x35 && x15 && x16 && ~x5 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x69 && ~x17 && x19 && ~x18 && ~x35 && x15 && x16 && ~x5 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x69 && ~x17 && x19 && ~x18 && ~x35 && x15 && ~x16 && x1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x17 && x19 && ~x18 && ~x35 && x15 && ~x16 && ~x1 )
						nx_state = s42;
					else if( ~x69 && ~x17 && x19 && ~x18 && ~x35 && ~x15 && x16 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x17 && x19 && ~x18 && ~x35 && ~x15 && ~x16 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x69 && ~x17 && x19 && ~x18 && ~x35 && ~x15 && ~x16 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x17 && ~x19 && x18 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && ~x17 && ~x19 && ~x18 && x40 && x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x69 && ~x17 && ~x19 && ~x18 && x40 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && ~x17 && ~x19 && ~x18 && x40 && ~x3 && ~x4 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s543;
						end
					else if( ~x69 && ~x17 && ~x19 && ~x18 && ~x40 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else nx_state = s42;
				s43 : if( x69 && x62 && x13 && x10 && x6 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && x62 && x13 && x10 && ~x6 && x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && x62 && x13 && x10 && ~x6 && ~x4 )
						nx_state = s1;
					else if( x69 && x62 && x13 && ~x10 )
						nx_state = s1;
					else if( x69 && x62 && ~x13 && x12 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && x62 && ~x13 && ~x12 && x10 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s541;
						end
					else if( x69 && x62 && ~x13 && ~x12 && ~x10 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && ~x62 && x17 && x18 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s551;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x7 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s542;
						end
					else if( x69 && ~x62 && x17 && ~x18 )
						nx_state = s43;
					else if( x69 && ~x62 && ~x17 && x18 && x15 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s541;
						end
					else if( x69 && ~x62 && ~x17 && x18 && ~x15 )
						nx_state = s1;
					else if( x69 && ~x62 && ~x17 && ~x18 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x69 && x63 && x42 && x43 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s183;
						end
					else if( ~x69 && x63 && x42 && ~x43 && x44 && x10 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x69 && x63 && x42 && ~x43 && x44 && ~x10 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s183;
						end
					else if( ~x69 && x63 && x42 && ~x43 && ~x44 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s183;
						end
					else if( ~x69 && x63 && ~x42 && x12 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s183;
						end
					else if( ~x69 && x63 && ~x42 && ~x12 && x13 && x14 && x41 && x37 && x2 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x63 && ~x42 && ~x12 && x13 && x14 && x41 && x37 && ~x2 )
						nx_state = s43;
					else if( ~x69 && x63 && ~x42 && ~x12 && x13 && x14 && x41 && ~x37 && x2 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x69 && x63 && ~x42 && ~x12 && x13 && x14 && x41 && ~x37 && ~x2 )
						nx_state = s43;
					else if( ~x69 && x63 && ~x42 && ~x12 && x13 && x14 && ~x41 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s183;
						end
					else if( ~x69 && x63 && ~x42 && ~x12 && x13 && ~x14 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s183;
						end
					else if( ~x69 && x63 && ~x42 && ~x12 && ~x13 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s183;
						end
					else if( ~x69 && ~x63 && x18 && x17 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s551;
						end
					else if( ~x69 && ~x63 && x18 && x17 && ~x7 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s542;
						end
					else if( ~x69 && ~x63 && x18 && ~x17 && x19 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s541;
						end
					else if( ~x69 && ~x63 && x18 && ~x17 && ~x19 && x15 && x16 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x69 && ~x63 && x18 && ~x17 && ~x19 && x15 && x16 && ~x5 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x69 && ~x63 && x18 && ~x17 && ~x19 && x15 && x16 && ~x5 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x69 && ~x63 && x18 && ~x17 && ~x19 && x15 && ~x16 && x1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x63 && x18 && ~x17 && ~x19 && x15 && ~x16 && ~x1 )
						nx_state = s43;
					else if( ~x69 && ~x63 && x18 && ~x17 && ~x19 && ~x15 && x16 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x63 && x18 && ~x17 && ~x19 && ~x15 && ~x16 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x69 && ~x63 && x18 && ~x17 && ~x19 && ~x15 && ~x16 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x63 && ~x18 && x17 )
						nx_state = s43;
					else if( ~x69 && ~x63 && ~x18 && ~x17 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s543;
						end
					else nx_state = s43;
				s44 : if( x69 && x62 && x13 && x10 && x7 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && x62 && x13 && x10 && ~x7 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && x62 && x13 && ~x10 )
						nx_state = s1;
					else if( x69 && x62 && ~x13 && x12 && x15 && x9 )
						nx_state = s44;
					else if( x69 && x62 && ~x13 && x12 && x15 && ~x9 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && x62 && ~x13 && x12 && ~x15 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && x62 && ~x13 && ~x12 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && x17 && x18 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s544;
						end
					else if( x69 && ~x62 && x17 && ~x18 && x14 && x5 )
						nx_state = s44;
					else if( x69 && ~x62 && x17 && ~x18 && x14 && ~x5 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && ~x62 && x17 && ~x18 && ~x14 && x5 )
						nx_state = s44;
					else if( x69 && ~x62 && x17 && ~x18 && ~x14 && ~x5 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( x69 && ~x62 && ~x17 && x15 && x18 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && ~x17 && x15 && ~x18 && x4 && x1 )
						nx_state = s44;
					else if( x69 && ~x62 && ~x17 && x15 && ~x18 && x4 && ~x1 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && ~x62 && ~x17 && x15 && ~x18 && ~x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && ~x62 && ~x17 && ~x15 && x18 )
						nx_state = s1;
					else if( x69 && ~x62 && ~x17 && ~x15 && ~x18 )
						nx_state = s44;
					else if( ~x69 && x18 && x17 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s544;
						end
					else if( ~x69 && x18 && ~x17 && x19 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x18 && ~x17 && ~x19 && x15 && x16 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x69 && x18 && ~x17 && ~x19 && x15 && x16 && ~x5 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x69 && x18 && ~x17 && ~x19 && x15 && x16 && ~x5 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x69 && x18 && ~x17 && ~x19 && x15 && ~x16 && x1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && x18 && ~x17 && ~x19 && x15 && ~x16 && ~x1 )
						nx_state = s44;
					else if( ~x69 && x18 && ~x17 && ~x19 && ~x15 && x16 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && x18 && ~x17 && ~x19 && ~x15 && ~x16 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x69 && x18 && ~x17 && ~x19 && ~x15 && ~x16 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x18 && x17 && x14 && x5 )
						nx_state = s44;
					else if( ~x69 && ~x18 && x17 && x14 && ~x5 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( ~x69 && ~x18 && x17 && ~x14 && x5 )
						nx_state = s44;
					else if( ~x69 && ~x18 && x17 && ~x14 && ~x5 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x69 && ~x18 && ~x17 && x4 && x19 && x1 )
						nx_state = s44;
					else if( ~x69 && ~x18 && ~x17 && x4 && x19 && ~x1 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s543;
						end
					else if( ~x69 && ~x18 && ~x17 && x4 && ~x19 )
						nx_state = s44;
					else if( ~x69 && ~x18 && ~x17 && ~x4 && x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( ~x69 && ~x18 && ~x17 && ~x4 && ~x19 )
						nx_state = s44;
					else nx_state = s44;
				s45 : if( x69 && x62 && x13 && x10 && x9 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && x62 && x13 && x10 && ~x9 && x17 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && x62 && x13 && x10 && ~x9 && ~x17 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && x62 && x13 && ~x10 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && x62 && ~x13 && x12 && x1 && x2 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && x62 && ~x13 && x12 && x1 && ~x2 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && x62 && ~x13 && x12 && x1 && ~x2 && ~x3 )
						nx_state = s45;
					else if( x69 && x62 && ~x13 && x12 && ~x1 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && x62 && ~x13 && ~x12 && x1 && x5 && x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s540;
						end
					else if( x69 && x62 && ~x13 && ~x12 && x1 && x5 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x69 && x62 && ~x13 && ~x12 && x1 && x5 && ~x3 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && x62 && ~x13 && ~x12 && x1 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && x62 && ~x13 && ~x12 && ~x1 && x2 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && x62 && ~x13 && ~x12 && ~x1 && ~x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && ~x62 && x17 && x18 && x4 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x4 && x1 && x3 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x4 && x1 && ~x3 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x4 && ~x1 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && ~x62 && x17 && ~x18 && x11 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s45;
						end
					else if( x69 && ~x62 && x17 && ~x18 && ~x11 && x16 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && ~x62 && x17 && ~x18 && ~x11 && ~x16 )
						nx_state = s1;
					else if( x69 && ~x62 && ~x17 && x18 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 && x15 && x1 && x2 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 && x15 && x1 && ~x2 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 && x15 && x1 && ~x2 && ~x3 )
						nx_state = s45;
					else if( x69 && ~x62 && ~x17 && ~x18 && x15 && ~x1 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 && ~x15 && x2 && x1 && x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 && ~x15 && x2 && x1 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 && ~x15 && x2 && x1 && ~x3 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 && ~x15 && x2 && ~x1 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 && ~x15 && ~x2 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 && ~x15 && ~x2 && ~x1 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x18 && x17 && x4 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( ~x69 && x18 && x17 && ~x4 && x40 && x31 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x18 && x17 && ~x4 && x40 && ~x31 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x69 && x18 && x17 && ~x4 && ~x40 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s543;
						end
					else if( ~x69 && x18 && ~x17 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( ~x69 && ~x18 && x17 && x11 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s45;
						end
					else if( ~x69 && ~x18 && x17 && ~x11 && x16 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( ~x69 && ~x18 && x17 && ~x11 && ~x16 && x15 && x1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x18 && x17 && ~x11 && ~x16 && x15 && ~x1 )
						nx_state = s45;
					else if( ~x69 && ~x18 && x17 && ~x11 && ~x16 && ~x15 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x69 && ~x18 && x17 && ~x11 && ~x16 && ~x15 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x18 && ~x17 && x19 && x1 && x39 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( ~x69 && ~x18 && ~x17 && x19 && x1 && ~x39 && x31 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && ~x18 && ~x17 && x19 && x1 && ~x39 && ~x31 )
						nx_state = s45;
					else if( ~x69 && ~x18 && ~x17 && x19 && ~x1 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x69 && ~x18 && ~x17 && ~x19 && x1 && x39 && x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x69 && ~x18 && ~x17 && ~x19 && x1 && x39 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && ~x18 && ~x17 && ~x19 && x1 && x39 && ~x3 && ~x4 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s543;
						end
					else if( ~x69 && ~x18 && ~x17 && ~x19 && x1 && ~x39 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( ~x69 && ~x18 && ~x17 && ~x19 && ~x1 && x2 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( ~x69 && ~x18 && ~x17 && ~x19 && ~x1 && ~x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else nx_state = s45;
				s46 : if( x2 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s46;
						end
					else if( x2 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s19;
						end
					else if( ~x2 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y8 = 1'b1;	
							nx_state = s552;
						end
					else if( ~x2 && ~x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s57;
						end
					else nx_state = s46;
				s47 : if( x70 && x62 )
						nx_state = s1;
					else if( x70 && ~x62 && x7 && x9 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x70 && ~x62 && x7 && ~x9 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x70 && ~x62 && x7 && ~x9 && ~x8 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x7 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && x60 && x61 && x15 && x2 && x12 && x7 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && x15 && x2 && x12 && ~x7 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s553;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && x15 && x2 && ~x12 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && x15 && x2 && ~x12 && ~x7 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && x15 && ~x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && x16 && x7 && x12 && x2 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s554;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && x16 && x7 && x12 && ~x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && x16 && x7 && ~x12 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && x12 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && x12 && ~x9 && x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && x12 && ~x9 && ~x11 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && x12 && ~x9 && ~x11 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && x12 && ~x9 && ~x11 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && x12 && ~x9 && ~x11 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && ~x12 && x11 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && ~x12 && x11 && ~x10 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && ~x12 && x11 && ~x10 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && ~x12 && x11 && ~x10 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && ~x12 && x11 && ~x10 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && ~x12 && ~x11 && x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && ~x12 && ~x11 && ~x8 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && ~x12 && ~x11 && ~x8 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && ~x12 && ~x11 && ~x8 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && ~x12 && ~x11 && ~x8 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && ~x16 && x2 && x7 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s555;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && ~x16 && x2 && ~x7 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x70 && x66 && x65 && x60 && x61 && ~x15 && ~x16 && ~x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x70 && x66 && x65 && x60 && ~x61 && x11 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && x60 && ~x61 && ~x11 && x7 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && x60 && ~x61 && ~x11 && ~x7 && x16 && x15 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x66 && x65 && x60 && ~x61 && ~x11 && ~x7 && x16 && x15 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x66 && x65 && x60 && ~x61 && ~x11 && ~x7 && x16 && x15 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( ~x70 && x66 && x65 && x60 && ~x61 && ~x11 && ~x7 && x16 && x15 && ~x18 )
						nx_state = s118;
					else if( ~x70 && x66 && x65 && x60 && ~x61 && ~x11 && ~x7 && x16 && ~x15 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && x60 && ~x61 && ~x11 && ~x7 && ~x16 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x60 && x61 && x62 && x16 && x11 && x12 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x70 && x66 && x65 && ~x60 && x61 && x62 && x16 && x11 && ~x12 && x13 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x70 && x66 && x65 && ~x60 && x61 && x62 && x16 && x11 && ~x12 && ~x13 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( ~x70 && x66 && x65 && ~x60 && x61 && x62 && x16 && ~x11 && x13 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x70 && x66 && x65 && ~x60 && x61 && x62 && x16 && ~x11 && ~x13 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x70 && x66 && x65 && ~x60 && x61 && x62 && ~x16 && x17 && x11 && x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s487;
						end
					else if( ~x70 && x66 && x65 && ~x60 && x61 && x62 && ~x16 && x17 && x11 && ~x13 && x2 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x70 && x66 && x65 && ~x60 && x61 && x62 && ~x16 && x17 && x11 && ~x13 && ~x2 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x70 && x66 && x65 && ~x60 && x61 && x62 && ~x16 && x17 && ~x11 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s487;
						end
					else if( ~x70 && x66 && x65 && ~x60 && x61 && x62 && ~x16 && ~x17 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && x66 && x65 && ~x60 && x61 && ~x62 && x11 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x60 && x61 && ~x62 && ~x11 && x7 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x60 && x61 && ~x62 && ~x11 && ~x7 && x16 && x15 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x66 && x65 && ~x60 && x61 && ~x62 && ~x11 && ~x7 && x16 && x15 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x66 && x65 && ~x60 && x61 && ~x62 && ~x11 && ~x7 && x16 && x15 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( ~x70 && x66 && x65 && ~x60 && x61 && ~x62 && ~x11 && ~x7 && x16 && x15 && ~x18 )
						nx_state = s118;
					else if( ~x70 && x66 && x65 && ~x60 && x61 && ~x62 && ~x11 && ~x7 && x16 && ~x15 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x60 && x61 && ~x62 && ~x11 && ~x7 && ~x16 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x60 && ~x61 && x62 && x18 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x66 && x65 && ~x60 && ~x61 && x62 && x18 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x66 && x65 && ~x60 && ~x61 && x62 && x18 && ~x13 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x60 && ~x61 && x62 && ~x18 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x60 && ~x61 && ~x62 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x66 && x65 && ~x60 && ~x61 && ~x62 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x66 && x65 && ~x60 && ~x61 && ~x62 && x19 && ~x13 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x60 && ~x61 && ~x62 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x65 && x21 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x65 && ~x21 && x22 && x23 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && x66 && ~x65 && ~x21 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x65 && ~x21 && ~x22 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x70 && x66 && ~x65 && ~x21 && ~x22 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x70 && x66 && ~x65 && ~x21 && ~x22 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x65 && ~x21 && ~x22 && x23 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x65 && ~x21 && ~x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x66 && x65 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && ~x66 && x65 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && ~x66 && x65 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && ~x66 && x65 && ~x4 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && x67 && x20 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && x67 && ~x20 && x21 )
						nx_state = s118;
					else if( ~x70 && ~x66 && ~x65 && x67 && ~x20 && ~x21 && x18 && x15 && x8 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x66 && ~x65 && x67 && ~x20 && ~x21 && x18 && x15 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s556;
						end
					else if( ~x70 && ~x66 && ~x65 && x67 && ~x20 && ~x21 && x18 && ~x15 && x16 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x70 && ~x66 && ~x65 && x67 && ~x20 && ~x21 && x18 && ~x15 && ~x16 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x70 && ~x66 && ~x65 && x67 && ~x20 && ~x21 && ~x18 )
						nx_state = s118;
					else if( ~x70 && ~x66 && ~x65 && ~x67 && x21 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && x3 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y9 = 1'b1;	
							nx_state = s173;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && x3 && ~x2 )
						nx_state = s47;
					else if( ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x3 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && x2 && x11 )
						nx_state = s47;
					else if( ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && x2 && ~x11 )
						nx_state = s47;
					else if( ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else nx_state = s47;
				s48 : if( x70 && x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s557;
						end
					else if( x70 && ~x3 && x2 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s46;
						end
					else if( x70 && ~x3 && x2 && ~x1 )
						begin
							y3 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							nx_state = s460;
						end
					else if( x70 && ~x3 && ~x2 && x1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( x70 && ~x3 && ~x2 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( ~x70 && x67 && x22 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x67 && x22 && ~x4 && x20 && x15 && x8 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x67 && x22 && ~x4 && x20 && x15 && ~x8 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && x67 && x22 && ~x4 && x20 && ~x15 && x16 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( ~x70 && x67 && x22 && ~x4 && x20 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( ~x70 && x67 && x22 && ~x4 && ~x20 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s558;
						end
					else if( ~x70 && x67 && ~x22 && x23 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x67 && ~x22 && ~x23 )
						nx_state = s1;
					else if( ~x70 && ~x67 && x61 && x60 && x3 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s559;
						end
					else if( ~x70 && ~x67 && x61 && x60 && ~x3 && x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s117;
						end
					else if( ~x70 && ~x67 && x61 && x60 && ~x3 && ~x18 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x70 && ~x67 && x61 && ~x60 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && ~x67 && x61 && ~x60 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && ~x67 && x61 && ~x60 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( ~x70 && ~x67 && x61 && ~x60 && x62 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x67 && x61 && ~x60 && ~x62 && x19 && x15 )
						nx_state = s143;
					else if( ~x70 && ~x67 && x61 && ~x60 && ~x62 && x19 && ~x15 && x16 )
						begin
							y12 = 1'b1;	
							nx_state = s244;
						end
					else if( ~x70 && ~x67 && x61 && ~x60 && ~x62 && x19 && ~x15 && ~x16 )
						nx_state = s143;
					else if( ~x70 && ~x67 && x61 && ~x60 && ~x62 && ~x19 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y24 = 1'b1;	
							nx_state = s136;
						end
					else if( ~x70 && ~x67 && ~x61 && x60 && x19 && x15 )
						nx_state = s143;
					else if( ~x70 && ~x67 && ~x61 && x60 && x19 && ~x15 && x16 )
						begin
							y12 = 1'b1;	
							nx_state = s244;
						end
					else if( ~x70 && ~x67 && ~x61 && x60 && x19 && ~x15 && ~x16 )
						nx_state = s143;
					else if( ~x70 && ~x67 && ~x61 && x60 && ~x19 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y24 = 1'b1;	
							nx_state = s136;
						end
					else if( ~x70 && ~x67 && ~x61 && ~x60 && x62 )
						nx_state = s1;
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && x18 && x15 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && x18 && x15 && ~x7 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && x18 && x15 && ~x7 && ~x11 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && x4 )
						nx_state = s47;
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && ~x4 && x11 && x9 )
						nx_state = s47;
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && ~x4 && x11 && ~x9 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && ~x4 && x11 && ~x9 && ~x7 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s559;
						end
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && ~x4 && ~x11 && x9 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && ~x4 && ~x11 && x9 && ~x7 && x10 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && ~x4 && ~x11 && x9 && ~x7 && ~x10 )
						nx_state = s47;
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && x7 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && x7 && ~x8 )
						nx_state = s47;
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && ~x7 && x12 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && ~x7 && ~x12 )
						nx_state = s47;
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && ~x18 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y24 = 1'b1;	
							nx_state = s136;
						end
					else nx_state = s48;
				s49 : if( x69 && x70 && x62 && x64 && x12 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x69 && x70 && x62 && x64 && ~x12 && x10 && x13 && x11 && x5 && x6 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s27;
						end
					else if( x69 && x70 && x62 && x64 && ~x12 && x10 && x13 && x11 && x5 && ~x6 && x7 )
						nx_state = s1;
					else if( x69 && x70 && x62 && x64 && ~x12 && x10 && x13 && x11 && x5 && ~x6 && ~x7 )
						begin
							y15 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s475;
						end
					else if( x69 && x70 && x62 && x64 && ~x12 && x10 && x13 && x11 && ~x5 && x4 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s476;
						end
					else if( x69 && x70 && x62 && x64 && ~x12 && x10 && x13 && x11 && ~x5 && ~x4 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && x70 && x62 && x64 && ~x12 && x10 && x13 && ~x11 && x14 && x4 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s27;
						end
					else if( x69 && x70 && x62 && x64 && ~x12 && x10 && x13 && ~x11 && x14 && ~x4 )
						nx_state = s49;
					else if( x69 && x70 && x62 && x64 && ~x12 && x10 && x13 && ~x11 && ~x14 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x69 && x70 && x62 && x64 && ~x12 && x10 && ~x13 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x69 && x70 && x62 && x64 && ~x12 && ~x10 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x6 && x3 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x6 && ~x3 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s18;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x6 && ~x3 && ~x1 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && ~x6 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && x66 && x5 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x64 && ~x65 && x66 && ~x5 && x1 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s35;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && x66 && ~x5 && ~x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && x18 && x17 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && x18 && x17 && ~x6 && x8 && x4 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s320;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && x18 && x17 && ~x6 && x8 && ~x4 && x1 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && x18 && x17 && ~x6 && x8 && ~x4 && x1 && ~x3 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && x18 && x17 && ~x6 && x8 && ~x4 && ~x1 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && x18 && x17 && ~x6 && ~x8 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && x18 && ~x17 && x19 && x9 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && x18 && ~x17 && x19 && ~x9 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && x18 && ~x17 && ~x19 && x4 && x5 && x3 )
						nx_state = s49;
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && x18 && ~x17 && ~x19 && x4 && x5 && ~x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && x18 && ~x17 && ~x19 && x4 && ~x5 && x3 )
						nx_state = s49;
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && x18 && ~x17 && ~x19 && x4 && ~x5 && ~x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && x18 && ~x17 && ~x19 && ~x4 && x3 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	
							nx_state = s20;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && x18 && ~x17 && ~x19 && ~x4 && ~x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && ~x18 && x17 && x12 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && ~x18 && x17 && ~x12 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && ~x18 && ~x17 && x19 && x2 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && ~x18 && ~x17 && x19 && ~x2 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x66 && ~x18 && ~x17 && ~x19 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && x70 && ~x62 && x66 && x12 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s560;
						end
					else if( x69 && x70 && ~x62 && x66 && x12 && ~x4 && x5 )
						begin
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s561;
						end
					else if( x69 && x70 && ~x62 && x66 && x12 && ~x4 && ~x5 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else if( x69 && x70 && ~x62 && x66 && ~x12 && x4 && x5 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && x70 && ~x62 && x66 && ~x12 && x4 && ~x5 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && x70 && ~x62 && x66 && ~x12 && ~x4 )
						begin
							y5 = 1'b1;	
							nx_state = s562;
						end
					else if( x69 && x70 && ~x62 && ~x66 && x20 && x21 && x12 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && ~x66 && x20 && x21 && x12 && ~x8 && x7 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && ~x66 && x20 && x21 && x12 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x66 && x20 && x21 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x66 && x20 && ~x21 && x7 && x6 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && ~x66 && x20 && ~x21 && x7 && ~x6 && x5 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && ~x66 && x20 && ~x21 && x7 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x66 && x20 && ~x21 && ~x7 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x66 && ~x20 && x6 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x69 && x70 && ~x62 && ~x66 && ~x20 && x6 && ~x7 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x69 && x70 && ~x62 && ~x66 && ~x20 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x66 && ~x20 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x66 && x68 && x21 && x20 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( x69 && ~x70 && x65 && x66 && x68 && x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x65 && x66 && x68 && x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x65 && x66 && x68 && x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x66 && x68 && x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x66 && x68 && ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && x66 && x68 && ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && x66 && x68 && ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x66 && x68 && ~x21 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && x7 && x12 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && x7 && ~x12 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s251;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && ~x7 && x12 && x14 && x11 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s564;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && ~x7 && x12 && x14 && ~x11 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && ~x7 && x12 && ~x14 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && ~x7 && x12 && ~x14 && x19 && ~x13 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && ~x7 && x12 && ~x14 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && ~x7 && ~x12 && x13 && x11 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s565;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && ~x7 && ~x12 && x13 && ~x11 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && ~x7 && ~x12 && ~x13 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && ~x7 && ~x12 && ~x13 && x19 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && ~x7 && ~x12 && ~x13 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && x11 && x7 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && x11 && ~x7 && x12 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && x11 && ~x7 && ~x12 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s555;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && ~x11 && x1 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && ~x11 && ~x1 && x12 && x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && ~x11 && ~x1 && x12 && ~x3 && x7 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && ~x11 && ~x1 && x12 && ~x3 && ~x7 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s555;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && ~x11 && ~x1 && ~x12 && x7 && x3 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s566;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && ~x11 && ~x1 && ~x12 && x7 && ~x3 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && ~x11 && ~x1 && ~x12 && ~x7 && x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && ~x11 && ~x1 && ~x12 && ~x7 && ~x3 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && x1 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && x7 && x12 && x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && x7 && x12 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s555;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && x7 && ~x12 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && x12 && x11 && x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && x12 && x11 && ~x3 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && x12 && ~x11 && x9 && x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && x12 && ~x11 && x9 && ~x3 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && x12 && ~x11 && ~x9 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && x12 && ~x11 && ~x9 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && x12 && ~x11 && ~x9 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && x12 && ~x11 && ~x9 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && x11 && x10 && x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && x11 && x10 && ~x3 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && x11 && ~x10 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && x11 && ~x10 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && x11 && ~x10 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && x11 && ~x10 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && ~x11 && x8 && x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && ~x11 && x8 && ~x3 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && ~x11 && ~x8 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && ~x11 && ~x8 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && ~x11 && ~x8 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && ~x11 && ~x8 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && ~x16 && x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && ~x16 && ~x3 && x7 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s555;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && ~x16 && ~x3 && ~x7 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s567;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && ~x60 && x62 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && ~x60 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && ~x60 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && ~x60 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( x69 && ~x70 && x65 && x66 && ~x68 && x61 && ~x60 && ~x62 && ~x18 )
						nx_state = s118;
					else if( x69 && ~x70 && x65 && x66 && ~x68 && ~x61 && x60 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && ~x61 && x60 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && ~x61 && x60 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( x69 && ~x70 && x65 && x66 && ~x68 && ~x61 && x60 && ~x18 )
						nx_state = s118;
					else if( x69 && ~x70 && x65 && x66 && ~x68 && ~x61 && ~x60 && x62 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x68 && ~x61 && ~x60 && ~x62 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x65 && ~x66 && x68 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && x65 && ~x66 && x68 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && x65 && ~x66 && x68 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && x68 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x23 && x22 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x23 && x22 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x23 && x22 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x23 && ~x22 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x23 && ~x22 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x23 && ~x22 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x23 && ~x22 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && ~x23 && x18 && x14 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && ~x23 && x18 && x14 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && ~x23 && x18 && ~x14 && x13 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && ~x23 && x18 && ~x14 && x13 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && ~x23 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x67 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && x67 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && x67 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x67 && x20 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x67 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && x21 && x68 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && x21 && x68 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && x21 && x68 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && x21 && x68 && ~x3 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && x21 && ~x68 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s174;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && x12 && x17 )
						begin
							y8 = 1'b1;	
							nx_state = s568;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && x12 && ~x17 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	
							nx_state = s569;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && ~x12 && x17 && x8 && x16 )
						begin
							y8 = 1'b1;	y22 = 1'b1;	
							nx_state = s570;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && ~x12 && x17 && x8 && ~x16 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s571;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && ~x12 && x17 && ~x8 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && ~x12 && x17 && ~x8 && x6 && ~x7 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && ~x12 && x17 && ~x8 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && ~x12 && ~x17 && x7 && x16 )
						begin
							y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s572;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && ~x12 && ~x17 && x7 && ~x16 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s571;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && ~x12 && ~x17 && ~x7 && x6 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && ~x12 && ~x17 && ~x7 && x6 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && ~x12 && ~x17 && ~x7 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && ~x19 && x16 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s573;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && ~x19 && x16 && ~x12 && x17 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s175;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && ~x19 && x16 && ~x12 && ~x17 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s379;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && ~x19 && ~x16 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && ~x19 && ~x16 && ~x2 && x3 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && ~x19 && ~x16 && ~x2 && ~x3 && x17 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s574;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && ~x19 && ~x16 && ~x2 && ~x3 && x17 && ~x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s574;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && ~x19 && ~x16 && ~x2 && ~x3 && ~x17 && x12 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s377;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && ~x19 && ~x16 && ~x2 && ~x3 && ~x17 && ~x12 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s377;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && x12 && x3 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && x12 && ~x3 && x17 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s379;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && x12 && ~x3 && ~x17 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && x16 && x17 && x3 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && x16 && x17 && ~x3 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s377;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && x16 && ~x17 && x15 && x3 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && x16 && ~x17 && x15 && ~x3 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s377;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && x16 && ~x17 && ~x15 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && x16 && ~x17 && ~x15 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && x16 && ~x17 && ~x15 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && x16 && ~x17 && ~x15 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && x17 && x14 && x3 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && x17 && x14 && ~x3 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s377;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && x17 && ~x14 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && x17 && ~x14 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && x17 && ~x14 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && x17 && ~x14 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && ~x17 && x13 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && ~x17 && x13 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && ~x17 && x13 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && ~x17 && x13 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && ~x17 && ~x13 && x3 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && ~x17 && ~x13 && ~x3 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s377;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && ~x19 && x3 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && ~x19 && ~x3 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s379;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && ~x19 && ~x3 && ~x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s574;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x22 && ~x68 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s358;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && x15 && x17 )
						begin
							y8 = 1'b1;	
							nx_state = s568;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && x15 && ~x17 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	
							nx_state = s569;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && ~x15 && x16 && x17 )
						begin
							y8 = 1'b1;	y22 = 1'b1;	
							nx_state = s570;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && ~x15 && x16 && ~x17 )
						begin
							y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s572;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && ~x15 && ~x16 && x17 && x10 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s377;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && ~x15 && ~x16 && x17 && ~x10 && x9 && x8 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && ~x15 && ~x16 && x17 && ~x10 && x9 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && ~x15 && ~x16 && x17 && ~x10 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && ~x15 && ~x16 && ~x17 && x9 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s377;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && ~x15 && ~x16 && ~x17 && ~x9 && x8 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && ~x15 && ~x16 && ~x17 && ~x9 && x8 && ~x10 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && ~x15 && ~x16 && ~x17 && ~x9 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && ~x19 && x16 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s575;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && ~x19 && ~x16 && x2 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s311;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && ~x19 && ~x16 && ~x2 && x5 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s576;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && ~x19 && ~x16 && ~x2 && ~x5 && x15 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s377;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && ~x19 && ~x16 && ~x2 && ~x5 && ~x15 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s377;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && x2 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s311;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && x15 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s576;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && x16 && x17 && x5 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s576;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && x16 && x17 && ~x5 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s377;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && x16 && ~x17 && x14 && x5 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s576;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && x16 && ~x17 && x14 && ~x5 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s377;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && x16 && ~x17 && ~x14 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && x16 && ~x17 && ~x14 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && x16 && ~x17 && ~x14 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && x16 && ~x17 && ~x14 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && x17 && x13 && x5 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s576;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && x17 && x13 && ~x5 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s377;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && x17 && ~x13 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && x17 && ~x13 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && x17 && ~x13 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && x17 && ~x13 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && ~x17 && x12 && x5 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s576;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && ~x17 && x12 && ~x5 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s377;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && ~x17 && ~x12 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && ~x17 && ~x12 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && ~x17 && ~x12 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && ~x17 && ~x12 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && ~x19 && x5 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s576;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && ~x19 && ~x5 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s575;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x22 && ~x68 )
						nx_state = s1;
					else if( ~x69 && x70 && x10 && x11 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s577;
						end
					else if( ~x69 && x70 && x10 && ~x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x69 && x70 && ~x10 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( ~x69 && x70 && ~x10 && ~x1 && x3 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x10 && ~x1 && ~x3 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s209;
						end
					else if( ~x69 && ~x70 && x45 && x44 && x16 && x22 && x29 && x27 && x15 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( ~x69 && ~x70 && x45 && x44 && x16 && x22 && x29 && x27 && ~x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && x45 && x44 && x16 && x22 && x29 && ~x27 )
						nx_state = s49;
					else if( ~x69 && ~x70 && x45 && x44 && x16 && x22 && ~x29 && x27 && x33 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && x45 && x44 && x16 && x22 && ~x29 && x27 && ~x33 && x18 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x69 && ~x70 && x45 && x44 && x16 && x22 && ~x29 && x27 && ~x33 && ~x18 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && x45 && x44 && x16 && x22 && ~x29 && ~x27 )
						nx_state = s49;
					else if( ~x69 && ~x70 && x45 && x44 && x16 && ~x22 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x45 && x44 && ~x16 && x37 && x21 && x1 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && x45 && x44 && ~x16 && x37 && x21 && ~x1 )
						nx_state = s49;
					else if( ~x69 && ~x70 && x45 && x44 && ~x16 && x37 && ~x21 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x45 && x44 && ~x16 && ~x37 && x25 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x45 && x44 && ~x16 && ~x37 && ~x25 && x5 && x4 )
						begin
							y8 = 1'b1;	y17 = 1'b1;	
							nx_state = s408;
						end
					else if( ~x69 && ~x70 && x45 && x44 && ~x16 && ~x37 && ~x25 && x5 && ~x4 )
						nx_state = s49;
					else if( ~x69 && ~x70 && x45 && x44 && ~x16 && ~x37 && ~x25 && ~x5 && x4 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && x45 && x44 && ~x16 && ~x37 && ~x25 && ~x5 && ~x4 )
						nx_state = s49;
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && x10 && x47 && x7 && x3 && x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && x10 && x47 && x7 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && x10 && x47 && x7 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && x10 && x47 && ~x7 && x9 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && x10 && x47 && ~x7 && ~x9 && x1 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && x10 && x47 && ~x7 && ~x9 && ~x1 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && x10 && ~x47 && x11 && x4 && x12 && x3 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && x10 && ~x47 && x11 && x4 && x12 && ~x3 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && x10 && ~x47 && x11 && x4 && ~x12 && x13 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && x10 && ~x47 && x11 && x4 && ~x12 && ~x13 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && x10 && ~x47 && x11 && x4 && ~x12 && ~x13 && ~x3 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && x10 && ~x47 && x11 && ~x4 )
						nx_state = s49;
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && x10 && ~x47 && ~x11 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && ~x10 && x11 && x47 && x5 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	
							nx_state = s213;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && ~x10 && x11 && x47 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && ~x10 && x11 && ~x47 && x13 && x4 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && ~x10 && x11 && ~x47 && x13 && ~x4 )
						nx_state = s49;
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && ~x10 && x11 && ~x47 && ~x13 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && ~x10 && ~x11 && x47 && x9 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && ~x10 && ~x11 && x47 && ~x9 && x1 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && ~x10 && ~x11 && x47 && ~x9 && ~x1 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && ~x10 && ~x11 && ~x47 && x12 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && ~x10 && ~x11 && ~x47 && ~x12 && x4 && x3 )
						begin
							y8 = 1'b1;	y17 = 1'b1;	
							nx_state = s408;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && ~x10 && ~x11 && ~x47 && ~x12 && x4 && ~x3 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && x46 && ~x10 && ~x11 && ~x47 && ~x12 && ~x4 )
						nx_state = s49;
					else if( ~x69 && ~x70 && x45 && ~x44 && ~x46 && x12 && x10 && x11 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && ~x46 && x12 && x10 && ~x11 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s578;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && ~x46 && x12 && ~x10 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && ~x46 && x12 && ~x10 && ~x1 && x3 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x45 && ~x44 && ~x46 && x12 && ~x10 && ~x1 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && ~x46 && ~x12 && x9 && x5 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && ~x46 && ~x12 && x9 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && ~x46 && ~x12 && ~x9 && x11 && x3 && x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && ~x46 && ~x12 && ~x9 && x11 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && ~x46 && ~x12 && ~x9 && x11 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && ~x46 && ~x12 && ~x9 && ~x11 && x5 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s176;
						end
					else if( ~x69 && ~x70 && x45 && ~x44 && ~x46 && ~x12 && ~x9 && ~x11 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x45 && x46 && x44 && x3 && x5 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x70 && ~x45 && x46 && x44 && x3 && ~x5 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s209;
						end
					else if( ~x69 && ~x70 && ~x45 && x46 && x44 && ~x3 && x10 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x70 && ~x45 && x46 && x44 && ~x3 && ~x10 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x69 && ~x70 && ~x45 && x46 && ~x44 && x47 && x8 && x7 && x3 && x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x69 && ~x70 && ~x45 && x46 && ~x44 && x47 && x8 && x7 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x45 && x46 && ~x44 && x47 && x8 && x7 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x45 && x46 && ~x44 && x47 && x8 && ~x7 && x5 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	
							nx_state = s213;
						end
					else if( ~x69 && ~x70 && ~x45 && x46 && ~x44 && x47 && x8 && ~x7 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x45 && x46 && ~x44 && x47 && ~x8 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && ~x45 && x46 && ~x44 && x47 && ~x8 && ~x1 && x3 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x45 && x46 && ~x44 && x47 && ~x8 && ~x1 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x45 && x46 && ~x44 && ~x47 && x9 && x5 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && ~x70 && ~x45 && x46 && ~x44 && ~x47 && x9 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x45 && x46 && ~x44 && ~x47 && ~x9 && x11 && x3 && x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x69 && ~x70 && ~x45 && x46 && ~x44 && ~x47 && ~x9 && x11 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x45 && x46 && ~x44 && ~x47 && ~x9 && x11 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x45 && x46 && ~x44 && ~x47 && ~x9 && ~x11 && x5 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s176;
						end
					else if( ~x69 && ~x70 && ~x45 && x46 && ~x44 && ~x47 && ~x9 && ~x11 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x46 && x44 && x7 && x9 && x8 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x46 && x44 && x7 && x9 && ~x8 )
						nx_state = s49;
					else if( ~x69 && ~x70 && ~x45 && ~x46 && x44 && x7 && ~x9 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x45 && ~x46 && x44 && ~x7 && x6 && x13 && x4 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s579;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x46 && x44 && ~x7 && x6 && x13 && ~x4 )
						nx_state = s49;
					else if( ~x69 && ~x70 && ~x45 && ~x46 && x44 && ~x7 && x6 && ~x13 && x4 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x46 && x44 && ~x7 && x6 && ~x13 && ~x4 )
						nx_state = s49;
					else if( ~x69 && ~x70 && ~x45 && ~x46 && x44 && ~x7 && ~x6 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x45 && ~x46 && ~x44 && x10 && x11 && x5 && x13 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x46 && ~x44 && x10 && x11 && x5 && ~x13 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s176;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x46 && ~x44 && x10 && x11 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x46 && ~x44 && x10 && ~x11 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x46 && ~x44 && ~x10 && x11 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							nx_state = s214;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x46 && ~x44 && ~x10 && x11 && ~x1 && x3 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x45 && ~x46 && ~x44 && ~x10 && x11 && ~x1 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x46 && ~x44 && ~x10 && ~x11 && x12 && x3 && x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x46 && ~x44 && ~x10 && ~x11 && x12 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x46 && ~x44 && ~x10 && ~x11 && x12 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x46 && ~x44 && ~x10 && ~x11 && ~x12 && x13 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							nx_state = s214;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x46 && ~x44 && ~x10 && ~x11 && ~x12 && x13 && ~x1 && x3 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x45 && ~x46 && ~x44 && ~x10 && ~x11 && ~x12 && x13 && ~x1 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x46 && ~x44 && ~x10 && ~x11 && ~x12 && ~x13 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s578;
						end
					else nx_state = s49;
				s50 : if( x69 && x70 && x62 && x64 )
						begin
							y1 = 1'b1;	y21 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s580;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && x5 && x6 && x30 && x36 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && x5 && x6 && x30 && ~x36 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && x5 && x6 && ~x30 && x31 && x33 && x34 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && x5 && x6 && ~x30 && x31 && x33 && ~x34 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && x5 && x6 && ~x30 && x31 && x33 && ~x34 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && x5 && x6 && ~x30 && x31 && x33 && ~x34 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && x5 && x6 && ~x30 && x31 && x33 && ~x34 && ~x27 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && x5 && x6 && ~x30 && x31 && ~x33 && x35 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && x5 && x6 && ~x30 && x31 && ~x33 && ~x35 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && x5 && x6 && ~x30 && x31 && ~x33 && ~x35 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && x5 && x6 && ~x30 && x31 && ~x33 && ~x35 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && x5 && x6 && ~x30 && x31 && ~x33 && ~x35 && ~x27 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && x5 && x6 && ~x30 && ~x31 && x32 )
						begin
							y1 = 1'b1;	y22 = 1'b1;	y37 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s581;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && x5 && x6 && ~x30 && ~x31 && ~x32 )
						begin
							y1 = 1'b1;	y20 = 1'b1;	y37 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s582;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && x5 && ~x6 && x7 && x23 && x24 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y15 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s583;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && x5 && ~x6 && x7 && x23 && ~x24 )
						begin
							y1 = 1'b1;	y33 = 1'b1;	y37 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s584;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && x5 && ~x6 && x7 && ~x23 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y39 = 1'b1;	
							nx_state = s584;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && x5 && ~x6 && ~x7 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	y33 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s585;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && ~x5 && x8 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	y33 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s585;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && ~x5 && ~x8 && x9 && x25 && x26 )
						begin
							y14 = 1'b1;	y19 = 1'b1;	y33 = 1'b1;	
							y37 = 1'b1;	y39 = 1'b1;	
							nx_state = s584;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && ~x5 && ~x8 && x9 && x25 && ~x26 )
						begin
							y14 = 1'b1;	y18 = 1'b1;	y33 = 1'b1;	
							y37 = 1'b1;	y39 = 1'b1;	
							nx_state = s584;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && ~x5 && ~x8 && x9 && ~x25 )
						begin
							y14 = 1'b1;	y17 = 1'b1;	y35 = 1'b1;	
							y37 = 1'b1;	y39 = 1'b1;	
							nx_state = s584;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && x4 && ~x5 && ~x8 && ~x9 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	y33 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s585;
						end
					else if( x69 && x70 && x62 && ~x64 && x65 && ~x4 )
						begin
							y1 = 1'b1;	y33 = 1'b1;	y37 = 1'b1;	
							y46 = 1'b1;	
							nx_state = s586;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && x17 && x18 && x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && x17 && x18 && ~x7 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s280;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && x17 && ~x18 )
						nx_state = s50;
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x17 && x18 && x19 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s215;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x17 && x18 && ~x19 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x64 && ~x65 && ~x17 && ~x18 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && x67 && x11 && x13 && x14 && x5 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && x67 && x11 && x13 && x14 && ~x5 && x1 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && x67 && x11 && x13 && x14 && ~x5 && ~x1 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && x67 && x11 && x13 && ~x14 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && x67 && x11 && x13 && ~x14 && ~x3 && x2 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x64 && x67 && x11 && x13 && ~x14 && ~x3 && ~x2 )
						nx_state = s50;
					else if( x69 && x70 && ~x62 && x63 && x64 && x67 && x11 && ~x13 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && x67 && x11 && ~x13 && ~x3 && x2 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x64 && x67 && x11 && ~x13 && ~x3 && ~x2 )
						nx_state = s50;
					else if( x69 && x70 && ~x62 && x63 && x64 && x67 && ~x11 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && x67 && ~x11 && ~x3 && x2 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x64 && x67 && ~x11 && ~x3 && ~x2 )
						nx_state = s50;
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && x14 && x13 && x10 && x15 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && x14 && x13 && x10 && x15 && ~x3 && x2 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && x14 && x13 && x10 && x15 && ~x3 && ~x2 )
						nx_state = s50;
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && x14 && x13 && x10 && ~x15 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && x14 && x13 && ~x10 && x15 && x5 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && x14 && x13 && ~x10 && x15 && ~x5 && x1 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && x14 && x13 && ~x10 && x15 && ~x5 && ~x1 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && x14 && x13 && ~x10 && ~x15 && x11 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && x14 && x13 && ~x10 && ~x15 && ~x11 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && x14 && x13 && ~x10 && ~x15 && ~x11 && ~x3 && x2 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && x14 && x13 && ~x10 && ~x15 && ~x11 && ~x3 && ~x2 )
						nx_state = s50;
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && x14 && ~x13 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && x14 && ~x13 && ~x3 && x2 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && x14 && ~x13 && ~x3 && ~x2 )
						nx_state = s50;
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && ~x14 && x9 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && ~x14 && x9 && ~x3 && x2 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && ~x14 && x9 && ~x3 && ~x2 )
						nx_state = s50;
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && ~x14 && ~x9 && x15 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && ~x14 && ~x9 && x15 && ~x3 && x2 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && ~x14 && ~x9 && x15 && ~x3 && ~x2 )
						nx_state = s50;
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && ~x14 && ~x9 && ~x15 && x7 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x67 && ~x14 && ~x9 && ~x15 && ~x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x64 && x66 && x7 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x64 && x66 && ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x64 && ~x66 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y4 = 1'b1;	
							nx_state = s71;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x65 && x66 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x65 && ~x66 && x67 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x65 && ~x66 && ~x67 && x21 && x15 )
						begin
							y44 = 1'b1;	y45 = 1'b1;	
							nx_state = s516;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x65 && ~x66 && ~x67 && x21 && ~x15 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x65 && ~x66 && ~x67 && x21 && ~x15 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x65 && ~x66 && ~x67 && x21 && ~x15 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x65 && ~x66 && ~x67 && x21 && ~x15 && ~x6 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x65 && ~x66 && ~x67 && ~x21 )
						begin
							y4 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y78 = 1'b1;	
							nx_state = s587;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && x19 && x12 )
						begin
							y54 = 1'b1;	
							nx_state = s525;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && x19 && ~x12 )
						begin
							y55 = 1'b1;	
							nx_state = s526;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && x12 && x6 )
						begin
							y16 = 1'b1;	y50 = 1'b1;	
							nx_state = s527;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && x12 && ~x6 && x16 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && x12 && ~x6 && ~x16 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && x12 && ~x6 && ~x16 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && x12 && ~x6 && ~x16 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && x12 && ~x6 && ~x16 && ~x9 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && ~x12 && x6 )
						begin
							y12 = 1'b1;	y48 = 1'b1;	
							nx_state = s529;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && ~x12 && ~x6 && x15 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && ~x12 && ~x6 && ~x15 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && ~x12 && ~x6 && ~x15 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && ~x12 && ~x6 && ~x15 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && ~x12 && ~x6 && ~x15 && ~x9 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && ~x18 && x19 )
						begin
							y27 = 1'b1;	y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s284;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && ~x18 && ~x19 && x6 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && ~x18 && ~x19 && ~x6 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && x19 && x6 && x12 && x11 )
						begin
							y46 = 1'b1;	
							nx_state = s531;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && x19 && x6 && x12 && ~x11 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && x19 && x6 && x12 && ~x11 && x9 && ~x10 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && x19 && x6 && x12 && ~x11 && ~x9 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && x19 && x6 && ~x12 && x10 )
						begin
							y46 = 1'b1;	
							nx_state = s531;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && x19 && x6 && ~x12 && ~x10 && x9 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && x19 && x6 && ~x12 && ~x10 && x9 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && x19 && x6 && ~x12 && ~x10 && ~x9 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && x19 && ~x6 && x12 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && x19 && ~x6 && ~x12 )
						begin
							y56 = 1'b1;	y57 = 1'b1;	
							nx_state = s284;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && x6 && x12 && x14 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && x6 && x12 && ~x14 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && x6 && x12 && ~x14 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && x6 && x12 && ~x14 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && x6 && x12 && ~x14 && ~x9 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && x6 && ~x12 && x13 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && x6 && ~x12 && ~x13 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && x6 && ~x12 && ~x13 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && x6 && ~x12 && ~x13 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && x6 && ~x12 && ~x13 && ~x9 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && ~x6 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && ~x18 && x19 && x12 && x6 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && ~x18 && x19 && x12 && ~x6 )
						begin
							y38 = 1'b1;	
							nx_state = s532;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && ~x18 && x19 && ~x12 && x6 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && ~x18 && x19 && ~x12 && ~x6 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && ~x18 && ~x19 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && x4 && x24 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && x4 && ~x24 && x23 && x9 && x10 && x8 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && x4 && ~x24 && x23 && x9 && x10 && ~x8 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && x4 && ~x24 && x23 && x9 && ~x10 && x8 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && x4 && ~x24 && x23 && x9 && ~x10 && ~x8 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && x4 && ~x24 && x23 && ~x9 && x10 && x8 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && x4 && ~x24 && x23 && ~x9 && x10 && ~x8 )
						begin
							y25 = 1'b1;	
							nx_state = s53;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && x4 && ~x24 && x23 && ~x9 && ~x10 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && x4 && ~x24 && x23 && ~x9 && ~x10 && ~x8 )
						begin
							y23 = 1'b1;	
							nx_state = s588;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && x4 && ~x24 && ~x23 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && x23 && x24 && x6 && x5 && x10 && x11 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && x23 && x24 && x6 && x5 && x10 && ~x11 && x12 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && x23 && x24 && x6 && x5 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && x23 && x24 && x6 && x5 && ~x10 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && x23 && x24 && x6 && ~x5 && x7 && x8 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && x23 && x24 && x6 && ~x5 && x7 && ~x8 && x10 && x11 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && x23 && x24 && x6 && ~x5 && x7 && ~x8 && x10 && ~x11 && x12 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && x23 && x24 && x6 && ~x5 && x7 && ~x8 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && x23 && x24 && x6 && ~x5 && x7 && ~x8 && ~x10 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && x23 && x24 && x6 && ~x5 && ~x7 && x9 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && x23 && x24 && x6 && ~x5 && ~x7 && ~x9 && x10 && x11 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && x23 && x24 && x6 && ~x5 && ~x7 && ~x9 && x10 && ~x11 && x12 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && x23 && x24 && x6 && ~x5 && ~x7 && ~x9 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && x23 && x24 && x6 && ~x5 && ~x7 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && x23 && x24 && ~x6 && x7 && x5 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && x23 && x24 && ~x6 && x7 && ~x5 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && x23 && x24 && ~x6 && ~x7 && x5 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && x23 && x24 && ~x6 && ~x7 && ~x5 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && x23 && ~x24 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && ~x23 && x24 && x8 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && ~x23 && x24 && ~x8 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && ~x23 && ~x24 && x9 && x10 && x8 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && ~x23 && ~x24 && x9 && x10 && ~x8 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && ~x23 && ~x24 && x9 && ~x10 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && ~x23 && ~x24 && x9 && ~x10 && ~x8 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && ~x23 && ~x24 && ~x9 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && ~x23 && ~x24 && ~x9 && x8 && ~x10 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x4 && ~x23 && ~x24 && ~x9 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && ~x67 && x30 && x31 )
						begin
							y33 = 1'b1;	
							nx_state = s589;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && ~x67 && x30 && ~x31 )
						begin
							y24 = 1'b1;	
							nx_state = s590;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && ~x67 && ~x30 )
						begin
							y47 = 1'b1;	y52 = 1'b1;	y61 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s353;
						end
					else if( x69 && ~x70 && x65 && x66 && x22 && x20 && x15 && x8 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && x66 && x22 && x20 && x15 && ~x8 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && x65 && x66 && x22 && x20 && ~x15 && x16 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x69 && ~x70 && x65 && x66 && x22 && x20 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( x69 && ~x70 && x65 && x66 && x22 && ~x20 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s558;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x22 && x23 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x66 && ~x22 && ~x23 && x3 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s558;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x22 && ~x23 && ~x3 && x19 && x15 && x8 )
						begin
							y11 = 1'b1;	
							nx_state = s91;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x22 && ~x23 && ~x3 && x19 && x15 && ~x8 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s591;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x22 && ~x23 && ~x3 && x19 && ~x15 && x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s126;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x22 && ~x23 && ~x3 && x19 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x22 && ~x23 && ~x3 && ~x19 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s592;
						end
					else if( x69 && ~x70 && x65 && ~x66 && x68 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && x21 && x5 )
						begin
							y31 = 1'b1;	
							nx_state = s164;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && x21 && ~x5 && x17 && x15 && x9 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && x21 && ~x5 && x17 && x15 && ~x9 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && x21 && ~x5 && x17 && ~x15 && x16 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && x21 && ~x5 && x17 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s333;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && x21 && ~x5 && ~x17 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s494;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && x15 && x9 && x23 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && x15 && x9 && ~x23 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && x15 && ~x9 && x23 && x6 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && x15 && ~x9 && x23 && ~x6 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && x15 && ~x9 && ~x23 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && x9 && x8 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && x9 && ~x8 && x10 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && x9 && ~x8 && ~x10 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && x9 && ~x8 && ~x10 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && x9 && ~x8 && ~x10 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && x9 && ~x8 && ~x10 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && x9 && ~x8 && ~x10 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && x8 && x12 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && x8 && ~x12 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && x8 && ~x12 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && x8 && ~x12 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && x8 && ~x12 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && x8 && ~x12 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && ~x8 && x11 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && ~x8 && ~x11 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && ~x8 && ~x11 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && ~x8 && ~x11 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && ~x8 && ~x11 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && ~x8 && ~x11 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && ~x16 && x6 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s495;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && ~x16 && ~x6 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && ~x23 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s495;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && ~x22 && x23 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && ~x22 && x23 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && ~x22 && x23 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && ~x22 && x23 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && ~x22 && ~x23 && x18 && x14 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && ~x22 && ~x23 && x18 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && ~x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x68 && ~x21 && ~x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && x62 && x6 && x15 && x8 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s593;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && x62 && x6 && x15 && ~x8 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && x62 && x6 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s593;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && x62 && x6 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s299;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && x62 && ~x6 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s593;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && x63 && x17 && x13 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && x63 && x17 && ~x13 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && x14 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && x14 && ~x8 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && ~x14 && x7 && x8 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s296;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && ~x14 && x7 && ~x8 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s297;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && ~x14 && ~x7 && x8 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && ~x14 && ~x7 && x8 && ~x12 && x19 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && ~x14 && ~x7 && x8 && ~x12 && x19 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && ~x14 && ~x7 && x8 && ~x12 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && ~x14 && ~x7 && ~x8 && x13 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && ~x14 && ~x7 && ~x8 && ~x13 && x19 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && ~x14 && ~x7 && ~x8 && ~x13 && x19 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && ~x14 && ~x7 && ~x8 && ~x13 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && ~x4 && x7 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s298;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && ~x4 && ~x7 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s435;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && ~x4 && ~x7 && ~x3 && x8 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && ~x4 && ~x7 && ~x3 && ~x8 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s435;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && x7 && x11 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && x7 && ~x11 && x8 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && x7 && ~x11 && ~x8 && x19 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && x7 && ~x11 && ~x8 && x19 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && x7 && ~x11 && ~x8 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && x7 && ~x11 && ~x8 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && ~x7 && x8 && x9 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && ~x7 && x8 && ~x9 && x19 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && ~x7 && x8 && ~x9 && x19 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && ~x7 && x8 && ~x9 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && ~x7 && x8 && ~x9 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && ~x7 && ~x8 && x10 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && ~x7 && ~x8 && ~x10 && x19 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && ~x7 && ~x8 && ~x10 && x19 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && ~x7 && ~x8 && ~x10 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && ~x7 && ~x8 && ~x10 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && ~x4 && x15 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && ~x4 && ~x15 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s468;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && ~x64 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && ~x64 && x15 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && ~x64 && ~x15 && x16 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && ~x64 && ~x15 && ~x16 && x14 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s299;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x62 && ~x63 && ~x64 && ~x15 && ~x16 && ~x14 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s295;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && x21 && x68 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && x21 && x68 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && x21 && x68 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && x21 && x68 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && x21 && ~x68 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && x21 && ~x68 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && x21 && ~x68 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && x21 && ~x68 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && x68 && x17 && x10 && x15 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s334;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && x68 && x17 && x10 && ~x15 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && x68 && x17 && ~x10 )
						begin
							y13 = 1'b1;	y16 = 1'b1;	
							nx_state = s335;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && x68 && ~x17 && x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && x68 && ~x17 && ~x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && x23 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && x10 && x12 && x18 && x14 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && x10 && x12 && x18 && ~x14 && x13 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && x10 && x12 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && x10 && x12 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && x10 && ~x12 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && ~x10 && x18 && x14 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && ~x10 && x18 && ~x14 && x13 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && ~x10 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && ~x10 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && ~x22 && x68 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && ~x22 && ~x68 && x23 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s362;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x23 && x15 && x9 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s361;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x23 && x15 && ~x9 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x23 && ~x15 && x16 && x7 && x9 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s274;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x23 && ~x15 && x16 && x7 && ~x9 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s275;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x23 && ~x15 && x16 && ~x7 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s274;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x23 && ~x15 && ~x16 )
						begin
							y14 = 1'b1;	
							nx_state = s366;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && x68 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	
							nx_state = s594;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && x19 && x13 && x20 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && x19 && x13 && x20 && ~x15 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && x19 && x13 && ~x20 )
						begin
							y2 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s385;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && x20 && x14 && x15 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && x20 && x14 && ~x15 )
						begin
							y22 = 1'b1;	y25 = 1'b1;	
							nx_state = s315;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && x20 && ~x14 && x15 && x4 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s595;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && x20 && ~x14 && x15 && ~x4 && x9 && x3 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && x20 && ~x14 && x15 && ~x4 && x9 && ~x3 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && x20 && ~x14 && x15 && ~x4 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && x20 && ~x14 && ~x15 && x3 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s595;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && x20 && ~x14 && ~x15 && ~x3 && x9 && x4 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && x20 && ~x14 && ~x15 && ~x3 && x9 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && x20 && ~x14 && ~x15 && ~x3 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && ~x20 && x14 )
						begin
							y2 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s385;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && ~x20 && ~x14 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s384;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && ~x20 && ~x14 && ~x5 && x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y9 = 1'b1;	
							nx_state = s173;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && ~x20 && ~x14 && ~x5 && ~x6 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && ~x20 && ~x14 && ~x5 && ~x6 && ~x15 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	
							nx_state = s315;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && ~x19 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s384;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && x14 && x18 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							nx_state = s315;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && x14 && ~x18 && x15 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							nx_state = s315;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && x14 && ~x18 && ~x15 && x9 && x3 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && x14 && ~x18 && ~x15 && x9 && ~x3 && x4 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && x14 && ~x18 && ~x15 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && x14 && ~x18 && ~x15 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && ~x14 && x15 && x16 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							nx_state = s315;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && ~x14 && x15 && ~x16 && x9 && x3 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && ~x14 && x15 && ~x16 && x9 && ~x3 && x4 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && ~x14 && x15 && ~x16 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && ~x14 && x15 && ~x16 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && ~x14 && ~x15 && x17 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							nx_state = s315;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && ~x14 && ~x15 && ~x17 && x9 && x3 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && ~x14 && ~x15 && ~x17 && x9 && ~x3 && x4 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && ~x14 && ~x15 && ~x17 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && ~x14 && ~x15 && ~x17 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && ~x20 && x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y9 = 1'b1;	
							nx_state = s173;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && ~x20 && ~x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	y23 = 1'b1;	
							nx_state = s383;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x21 && x68 && x22 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x21 && x68 && x22 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x21 && x68 && x22 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x21 && x68 && x22 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x21 && x68 && ~x22 && x15 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	
							nx_state = s594;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x21 && x68 && ~x22 && ~x15 && x19 && x18 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	
							nx_state = s594;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x21 && x68 && ~x22 && ~x15 && x19 && ~x18 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x21 && x68 && ~x22 && ~x15 && x19 && ~x18 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x21 && x68 && ~x22 && ~x15 && x19 && ~x18 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x21 && x68 && ~x22 && ~x15 && x19 && ~x18 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x21 && x68 && ~x22 && ~x15 && ~x19 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	
							nx_state = s594;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x21 && ~x68 && x22 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s174;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x21 && ~x68 && ~x22 && x9 && x11 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x21 && ~x68 && ~x22 && x9 && ~x11 && x2 )
						nx_state = s50;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x21 && ~x68 && ~x22 && x9 && ~x11 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x21 && ~x68 && ~x22 && ~x9 && x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s174;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x21 && ~x68 && ~x22 && ~x9 && ~x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x69 && x45 && x44 && x17 && x19 && x10 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s387;
						end
					else if( ~x69 && x45 && x44 && x17 && x19 && ~x10 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x69 && x45 && x44 && x17 && ~x19 )
						nx_state = s50;
					else if( ~x69 && x45 && x44 && ~x17 && x20 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x69 && x45 && x44 && ~x17 && ~x20 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && x45 && x44 && ~x17 && ~x20 && ~x2 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && x45 && ~x44 && x46 && x10 && x47 && x7 && x3 && x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x69 && x45 && ~x44 && x46 && x10 && x47 && x7 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && x45 && ~x44 && x46 && x10 && x47 && x7 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && x45 && ~x44 && x46 && x10 && x47 && ~x7 && x9 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && x45 && ~x44 && x46 && x10 && x47 && ~x7 && ~x9 && x1 )
						nx_state = s1;
					else if( ~x69 && x45 && ~x44 && x46 && x10 && x47 && ~x7 && ~x9 && ~x1 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && x45 && ~x44 && x46 && x10 && ~x47 && x6 && x2 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s387;
						end
					else if( ~x69 && x45 && ~x44 && x46 && x10 && ~x47 && x6 && ~x2 )
						nx_state = s50;
					else if( ~x69 && x45 && ~x44 && x46 && x10 && ~x47 && ~x6 && x2 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x69 && x45 && ~x44 && x46 && x10 && ~x47 && ~x6 && ~x2 )
						nx_state = s50;
					else if( ~x69 && x45 && ~x44 && x46 && ~x10 && x47 && x11 && x5 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	
							nx_state = s213;
						end
					else if( ~x69 && x45 && ~x44 && x46 && ~x10 && x47 && x11 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && x45 && ~x44 && x46 && ~x10 && x47 && ~x11 && x9 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && x45 && ~x44 && x46 && ~x10 && x47 && ~x11 && ~x9 && x1 )
						nx_state = s1;
					else if( ~x69 && x45 && ~x44 && x46 && ~x10 && x47 && ~x11 && ~x9 && ~x1 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && x45 && ~x44 && x46 && ~x10 && ~x47 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x69 && x45 && ~x44 && x46 && ~x10 && ~x47 && ~x1 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && x45 && ~x44 && x46 && ~x10 && ~x47 && ~x1 && ~x2 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && x45 && ~x44 && ~x46 && x12 && x10 && x8 && x1 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && x45 && ~x44 && ~x46 && x12 && x10 && x8 && ~x1 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && x45 && ~x44 && ~x46 && x12 && x10 && ~x8 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && x45 && ~x44 && ~x46 && x12 && ~x10 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x69 && x45 && ~x44 && ~x46 && x12 && ~x10 && ~x1 && x3 )
						nx_state = s1;
					else if( ~x69 && x45 && ~x44 && ~x46 && x12 && ~x10 && ~x1 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && x45 && ~x44 && ~x46 && ~x12 && x9 && x5 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && x45 && ~x44 && ~x46 && ~x12 && x9 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && x45 && ~x44 && ~x46 && ~x12 && ~x9 && x10 && x5 && x11 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && x45 && ~x44 && ~x46 && ~x12 && ~x9 && x10 && x5 && ~x11 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							nx_state = s214;
						end
					else if( ~x69 && x45 && ~x44 && ~x46 && ~x12 && ~x9 && x10 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && x45 && ~x44 && ~x46 && ~x12 && ~x9 && ~x10 && x11 && x3 && x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x69 && x45 && ~x44 && ~x46 && ~x12 && ~x9 && ~x10 && x11 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && x45 && ~x44 && ~x46 && ~x12 && ~x9 && ~x10 && x11 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && x45 && ~x44 && ~x46 && ~x12 && ~x9 && ~x10 && ~x11 && x5 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s176;
						end
					else if( ~x69 && x45 && ~x44 && ~x46 && ~x12 && ~x9 && ~x10 && ~x11 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x45 && x44 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x69 && ~x45 && x44 && ~x1 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x45 && x44 && ~x1 && ~x2 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x45 && ~x44 && x46 && x47 && x8 && x7 && x3 && x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x69 && ~x45 && ~x44 && x46 && x47 && x8 && x7 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x45 && ~x44 && x46 && x47 && x8 && x7 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x45 && ~x44 && x46 && x47 && x8 && ~x7 && x5 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	
							nx_state = s213;
						end
					else if( ~x69 && ~x45 && ~x44 && x46 && x47 && x8 && ~x7 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x45 && ~x44 && x46 && x47 && ~x8 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x45 && ~x44 && x46 && x47 && ~x8 && ~x1 && x3 )
						nx_state = s1;
					else if( ~x69 && ~x45 && ~x44 && x46 && x47 && ~x8 && ~x1 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x45 && ~x44 && x46 && ~x47 && x9 && x5 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && ~x45 && ~x44 && x46 && ~x47 && x9 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x45 && ~x44 && x46 && ~x47 && ~x9 && x10 && x5 && x11 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && ~x45 && ~x44 && x46 && ~x47 && ~x9 && x10 && x5 && ~x11 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							nx_state = s214;
						end
					else if( ~x69 && ~x45 && ~x44 && x46 && ~x47 && ~x9 && x10 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x45 && ~x44 && x46 && ~x47 && ~x9 && ~x10 && x11 && x3 && x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x69 && ~x45 && ~x44 && x46 && ~x47 && ~x9 && ~x10 && x11 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x45 && ~x44 && x46 && ~x47 && ~x9 && ~x10 && x11 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x45 && ~x44 && x46 && ~x47 && ~x9 && ~x10 && ~x11 && x5 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s176;
						end
					else if( ~x69 && ~x45 && ~x44 && x46 && ~x47 && ~x9 && ~x10 && ~x11 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x45 && ~x44 && ~x46 && x10 && x11 && x5 && x13 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && ~x45 && ~x44 && ~x46 && x10 && x11 && x5 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							nx_state = s214;
						end
					else if( ~x69 && ~x45 && ~x44 && ~x46 && x10 && x11 && x5 && ~x13 && ~x12 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s176;
						end
					else if( ~x69 && ~x45 && ~x44 && ~x46 && x10 && x11 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x45 && ~x44 && ~x46 && x10 && ~x11 && x8 && x1 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && ~x45 && ~x44 && ~x46 && x10 && ~x11 && x8 && ~x1 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x45 && ~x44 && ~x46 && x10 && ~x11 && ~x8 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && ~x45 && ~x44 && ~x46 && ~x10 && x12 && x11 && x5 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && ~x45 && ~x44 && ~x46 && ~x10 && x12 && x11 && ~x5 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x45 && ~x44 && ~x46 && ~x10 && x12 && ~x11 && x3 && x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x69 && ~x45 && ~x44 && ~x46 && ~x10 && x12 && ~x11 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x45 && ~x44 && ~x46 && ~x10 && x12 && ~x11 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x69 && ~x45 && ~x44 && ~x46 && ~x10 && ~x12 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							nx_state = s214;
						end
					else if( ~x69 && ~x45 && ~x44 && ~x46 && ~x10 && ~x12 && ~x1 && x3 )
						nx_state = s1;
					else if( ~x69 && ~x45 && ~x44 && ~x46 && ~x10 && ~x12 && ~x1 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else nx_state = s50;
				s51 : if( x69 && x70 && x62 && x17 && x18 && x65 && x19 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y17 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s389;
						end
					else if( x69 && x70 && x62 && x17 && x18 && x65 && ~x19 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x70 && x62 && x17 && x18 && ~x65 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x69 && x70 && x62 && x17 && ~x18 && x65 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && x70 && x62 && x17 && ~x18 && ~x65 && x14 && x5 )
						nx_state = s51;
					else if( x69 && x70 && x62 && x17 && ~x18 && ~x65 && x14 && ~x5 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x70 && x62 && x17 && ~x18 && ~x65 && ~x14 && x5 )
						nx_state = s51;
					else if( x69 && x70 && x62 && x17 && ~x18 && ~x65 && ~x14 && ~x5 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && x70 && x62 && ~x17 && x18 && x65 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x70 && x62 && ~x17 && x18 && ~x65 && x19 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && x70 && x62 && ~x17 && x18 && ~x65 && ~x19 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x17 && ~x18 && x19 && x65 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && x70 && x62 && ~x17 && ~x18 && x19 && ~x65 && x4 && x1 )
						nx_state = s51;
					else if( x69 && x70 && x62 && ~x17 && ~x18 && x19 && ~x65 && x4 && ~x1 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && x62 && ~x17 && ~x18 && x19 && ~x65 && ~x4 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	
							nx_state = s20;
						end
					else if( x69 && x70 && x62 && ~x17 && ~x18 && ~x19 && x65 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x70 && x62 && ~x17 && ~x18 && ~x19 && ~x65 )
						nx_state = s51;
					else if( x69 && x70 && ~x62 && x64 && x63 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s596;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x66 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s597;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && ~x66 && x21 && x20 )
						begin
							y4 = 1'b1;	y64 = 1'b1;	
							nx_state = s598;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && ~x66 && x21 && ~x20 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && ~x66 && ~x21 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && x65 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x65 && x4 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x65 && ~x4 && x5 && x7 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s426;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x65 && ~x4 && x5 && ~x7 && x1 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x65 && ~x4 && x5 && ~x7 && x1 && ~x2 && x3 )
						nx_state = s51;
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x65 && ~x4 && x5 && ~x7 && x1 && ~x2 && ~x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x65 && ~x4 && x5 && ~x7 && ~x1 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x65 && ~x4 && ~x5 && x6 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	
							nx_state = s427;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x65 && ~x4 && ~x5 && ~x6 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s426;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x63 && x67 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x63 && ~x67 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x66 && x65 && x67 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x66 && x65 && x67 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x66 && x65 && x67 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && x67 && x22 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && x67 && ~x22 && x18 && x13 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && ~x70 && x66 && x65 && x67 && ~x22 && x18 && x13 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x66 && x65 && x67 && ~x22 && x18 && ~x13 && x12 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && ~x70 && x66 && x65 && x67 && ~x22 && x18 && ~x13 && x12 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x66 && x65 && x67 && ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && x67 && ~x22 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && x20 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && x3 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && x18 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y21 = 1'b1;	
							nx_state = s599;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && x15 && x10 && x11 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s600;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s601;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && x15 && x10 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y13 = 1'b1;	
							nx_state = s600;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s602;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && x10 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && x10 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && x10 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && x10 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && ~x10 && x12 && x11 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s603;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && ~x10 && x12 && ~x11 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && ~x10 && x12 && ~x11 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && ~x10 && x12 && ~x11 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && ~x10 && x12 && ~x11 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && ~x10 && ~x12 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && ~x10 && ~x12 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && ~x10 && ~x12 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && ~x10 && ~x12 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s604;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && ~x21 && x15 && x10 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && ~x21 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s605;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && ~x21 && x15 && x10 && ~x11 && ~x12 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s606;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && ~x21 && x15 && ~x10 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && ~x21 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s600;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && ~x21 && ~x15 && x16 && x10 && x12 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && ~x21 && ~x15 && x16 && x10 && ~x12 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && ~x21 && ~x15 && x16 && ~x10 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && ~x21 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s607;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x21 && x15 && x4 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x21 && x15 && x4 && ~x10 && x12 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x21 && x15 && x4 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x21 && x15 && ~x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x21 && ~x15 && x16 && x10 && x12 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x21 && ~x15 && x16 && x10 && ~x12 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s608;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x21 && ~x15 && x16 && ~x10 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x21 && ~x15 && ~x16 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x21 && ~x15 && ~x16 && ~x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x21 && x22 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x21 && ~x22 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s609;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x21 && ~x22 && ~x23 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x68 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x68 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x68 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && x68 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && x7 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && x7 && ~x9 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && x8 && x9 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s296;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && x8 && ~x9 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s297;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && ~x8 && x9 && x13 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && ~x8 && x9 && ~x13 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && ~x8 && x9 && ~x13 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && ~x8 && x9 && ~x13 && ~x19 && x17 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && ~x8 && x9 && ~x13 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && ~x8 && ~x9 && x14 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && ~x8 && ~x9 && ~x14 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && ~x8 && ~x9 && ~x14 && ~x19 && x17 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && ~x8 && ~x9 && ~x14 && ~x19 && x17 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && ~x8 && ~x9 && ~x14 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && ~x16 && x7 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s406;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && ~x16 && ~x7 && x8 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s406;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && ~x16 && ~x7 && ~x8 && x4 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && ~x16 && ~x7 && ~x8 && ~x4 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && ~x16 && ~x7 && ~x8 && ~x4 && ~x5 && x9 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && ~x16 && ~x7 && ~x8 && ~x4 && ~x5 && ~x9 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && x4 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && x9 && ~x10 && x8 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && x9 && ~x10 && ~x8 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && x9 && ~x10 && ~x8 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && x9 && ~x10 && ~x8 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && x9 && ~x10 && ~x8 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && x9 && ~x10 && ~x8 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && x8 && x12 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && x8 && ~x12 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && x8 && ~x12 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && x8 && ~x12 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && x8 && ~x12 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && x8 && ~x12 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && ~x8 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && ~x8 && ~x11 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && ~x8 && ~x11 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && ~x8 && ~x11 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && ~x8 && ~x11 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && ~x8 && ~x11 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && ~x16 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && ~x16 && ~x5 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s333;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && x2 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x2 && x17 && x15 && x9 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x2 && x17 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x2 && x17 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x2 && x17 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s495;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x2 && ~x17 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x20 && x15 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s556;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x20 && ~x15 )
						begin
							y7 = 1'b1;	y12 = 1'b1;	
							nx_state = s610;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else if( ~x69 && x70 && x26 && x8 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( ~x69 && x70 && x26 && x8 && ~x1 && x14 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( ~x69 && x70 && x26 && x8 && ~x1 && ~x14 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( ~x69 && x70 && x26 && ~x8 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s612;
						end
					else if( ~x69 && x70 && ~x26 && x28 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x26 && ~x28 && x6 && x7 && x5 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s613;
						end
					else if( ~x69 && x70 && ~x26 && ~x28 && x6 && x7 && x5 && ~x3 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && x70 && ~x26 && ~x28 && x6 && x7 && x5 && ~x3 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s614;
						end
					else if( ~x69 && x70 && ~x26 && ~x28 && x6 && x7 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( ~x69 && x70 && ~x26 && ~x28 && x6 && ~x7 && x8 )
						begin
							y10 = 1'b1;	
							nx_state = s405;
						end
					else if( ~x69 && x70 && ~x26 && ~x28 && x6 && ~x7 && ~x8 && x5 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s613;
						end
					else if( ~x69 && x70 && ~x26 && ~x28 && x6 && ~x7 && ~x8 && x5 && ~x3 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && x70 && ~x26 && ~x28 && x6 && ~x7 && ~x8 && x5 && ~x3 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s614;
						end
					else if( ~x69 && x70 && ~x26 && ~x28 && x6 && ~x7 && ~x8 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( ~x69 && x70 && ~x26 && ~x28 && ~x6 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s405;
						end
					else if( ~x69 && x70 && ~x26 && ~x28 && ~x6 && ~x24 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x44 && x45 && x13 && x23 && x42 && x40 )
						begin
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x13 && x23 && x42 && ~x40 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x13 && x23 && ~x42 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x13 && ~x23 )
						begin
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x13 && x28 && x35 && x5 )
						begin
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x13 && x28 && x35 && ~x5 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x13 && x28 && ~x35 && x14 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x44 && x45 && ~x13 && x28 && ~x35 && ~x14 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x13 && ~x28 && x6 && x35 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x13 && ~x28 && x6 && ~x35 && x14 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x44 && x45 && ~x13 && ~x28 && x6 && ~x35 && ~x14 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x13 && ~x28 && ~x6 && x39 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x13 && ~x28 && ~x6 && ~x39 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s387;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x46 && x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							nx_state = s38;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x46 && ~x3 && x5 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x46 && ~x3 && ~x5 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x46 && ~x3 && ~x5 && ~x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x46 && x11 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x46 && ~x11 && x3 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x46 && ~x11 && ~x3 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && ~x44 && x11 && x13 && x5 )
						begin
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x69 && ~x70 && ~x44 && x11 && x13 && ~x5 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && ~x44 && x11 && ~x13 && x10 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x69 && ~x70 && ~x44 && x11 && ~x13 && x10 && ~x5 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && ~x44 && x11 && ~x13 && ~x10 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && ~x44 && x11 && ~x13 && ~x10 && ~x1 && x3 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x44 && x11 && ~x13 && ~x10 && ~x1 && ~x3 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x11 && x10 )
						begin
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x11 && ~x10 && x12 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x11 && ~x10 && x12 && ~x1 && x3 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x44 && ~x11 && ~x10 && x12 && ~x1 && ~x3 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x11 && ~x10 && ~x12 && x13 && x3 && x6 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x11 && ~x10 && ~x12 && x13 && x3 && ~x6 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x11 && ~x10 && ~x12 && x13 && ~x3 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x11 && ~x10 && ~x12 && ~x13 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s387;
						end
					else nx_state = s51;
				s52 : if( 1'b1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s615;
						end
					else nx_state = s52;
				s53 : if( x63 )
						begin
							y26 = 1'b1;	
							nx_state = s262;
						end
					else if( ~x63 && x64 )
						begin
							y26 = 1'b1;	
							nx_state = s262;
						end
					else if( ~x63 && ~x64 && x67 )
						begin
							y26 = 1'b1;	
							nx_state = s262;
						end
					else if( ~x63 && ~x64 && ~x67 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else nx_state = s53;
				s54 : if( 1'b1 )
						begin
							y36 = 1'b1;	
							nx_state = s617;
						end
					else nx_state = s54;
				s55 : if( 1'b1 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							y16 = 1'b1;	y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s618;
						end
					else nx_state = s55;
				s56 : if( 1'b1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y14 = 1'b1;	y38 = 1'b1;	
							nx_state = s619;
						end
					else nx_state = s56;
				s57 : if( x70 && x62 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s18;
						end
					else if( x70 && x62 && ~x3 && x1 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s46;
						end
					else if( x70 && x62 && ~x3 && x1 && ~x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( x70 && x62 && ~x3 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( x70 && ~x62 && x63 && x66 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y15 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s620;
						end
					else if( x70 && ~x62 && x63 && ~x66 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y5 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s621;
						end
					else if( x70 && ~x62 && ~x63 && x64 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y5 = 1'b1;	
							y10 = 1'b1;	y16 = 1'b1;	
							nx_state = s622;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x66 && x67 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y5 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s623;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x66 && ~x67 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y5 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s624;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x66 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y5 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s621;
						end
					else if( ~x70 && x65 && x22 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && x65 && ~x22 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s625;
						end
					else if( ~x70 && ~x65 && x21 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x65 && ~x21 && x23 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x70 && ~x65 && ~x21 && ~x23 && x22 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x70 && ~x65 && ~x21 && ~x23 && ~x22 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else nx_state = s57;
				s58 : if( x70 && x62 && x6 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x70 && x62 && ~x6 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( x70 && ~x62 && x64 )
						begin
							y3 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s626;
						end
					else if( x70 && ~x62 && ~x64 && x65 && x15 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && ~x62 && ~x64 && x65 && ~x15 && x6 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x70 && ~x62 && ~x64 && x65 && ~x15 && ~x6 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( x70 && ~x62 && ~x64 && ~x65 && x10 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && ~x62 && ~x64 && ~x65 && ~x10 && x11 )
						begin
							y14 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s401;
						end
					else if( x70 && ~x62 && ~x64 && ~x65 && ~x10 && ~x11 )
						begin
							y10 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s402;
						end
					else if( ~x70 && x65 && x67 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && x67 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && x67 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x65 && x67 && x22 && ~x17 )
						nx_state = s1;
					else if( ~x70 && x65 && x67 && ~x22 && x18 && x13 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && x65 && x67 && ~x22 && x18 && x13 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x65 && x67 && ~x22 && x18 && ~x13 && x12 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && x65 && x67 && ~x22 && x18 && ~x13 && x12 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x65 && x67 && ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && x65 && x67 && ~x22 && ~x18 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x67 && x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x67 && x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x67 && x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x67 && x21 && x20 && ~x17 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x67 && x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x65 && ~x67 && x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x65 && ~x67 && x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x67 && x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x67 && ~x21 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( ~x70 && ~x65 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y21 = 1'b1;	
							nx_state = s121;
						end
					else nx_state = s58;
				s59 : if( x69 && x62 && x4 && x5 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( x69 && x62 && x4 && ~x5 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s627;
						end
					else if( x69 && x62 && ~x4 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else if( x69 && ~x62 && x16 && x15 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( x69 && ~x62 && x16 && ~x15 && x4 && x5 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( x69 && ~x62 && x16 && ~x15 && x4 && ~x5 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s627;
						end
					else if( x69 && ~x62 && x16 && ~x15 && ~x4 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else if( x69 && ~x62 && ~x16 && x15 && x6 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else if( x69 && ~x62 && ~x16 && x15 && ~x6 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y22 = 1'b1;	
							nx_state = s61;
						end
					else if( x69 && ~x62 && ~x16 && ~x15 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x69 && x10 && x6 && x7 && x2 && x64 && x3 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x69 && x10 && x6 && x7 && x2 && x64 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x69 && x10 && x6 && x7 && x2 && x64 && ~x3 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x69 && x10 && x6 && x7 && x2 && ~x64 && x41 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x69 && x10 && x6 && x7 && x2 && ~x64 && ~x41 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x69 && x10 && x6 && x7 && x2 && ~x64 && ~x41 && ~x4 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s631;
						end
					else if( ~x69 && x10 && x6 && x7 && ~x2 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x10 && x6 && ~x7 && x8 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x69 && x10 && x6 && ~x7 && ~x8 && x2 && x64 && x3 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x69 && x10 && x6 && ~x7 && ~x8 && x2 && x64 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x69 && x10 && x6 && ~x7 && ~x8 && x2 && x64 && ~x3 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x69 && x10 && x6 && ~x7 && ~x8 && x2 && ~x64 && x41 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x69 && x10 && x6 && ~x7 && ~x8 && x2 && ~x64 && ~x41 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x69 && x10 && x6 && ~x7 && ~x8 && x2 && ~x64 && ~x41 && ~x4 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s631;
						end
					else if( ~x69 && x10 && x6 && ~x7 && ~x8 && ~x2 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x10 && ~x6 && x64 && x2 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x69 && x10 && ~x6 && x64 && ~x2 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && x10 && ~x6 && ~x64 && x34 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x69 && x10 && ~x6 && ~x64 && ~x34 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x69 && ~x10 && x11 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x69 && ~x10 && x11 && ~x5 && x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && ~x10 && x11 && ~x5 && ~x6 && x64 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && ~x10 && x11 && ~x5 && ~x6 && ~x64 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else if( ~x69 && ~x10 && ~x11 && x64 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && ~x10 && ~x11 && ~x64 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else nx_state = s59;
				s60 : if( x62 && x4 && x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x62 && x4 && ~x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s633;
						end
					else if( x62 && ~x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s634;
						end
					else if( ~x62 && x15 && x6 && x16 && x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( ~x62 && x15 && x6 && x16 && ~x5 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x62 && x15 && x6 && ~x16 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x62 && x15 && ~x6 && x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( ~x62 && x15 && ~x6 && ~x16 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s636;
						end
					else if( ~x62 && ~x15 && x16 && x4 && x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x62 && ~x15 && x16 && x4 && ~x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s637;
						end
					else if( ~x62 && ~x15 && x16 && ~x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s634;
						end
					else if( ~x62 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else nx_state = s60;
				s61 : if( x62 && x4 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s627;
						end
					else if( x62 && ~x4 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else if( ~x62 && x16 && x15 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else if( ~x62 && x16 && ~x15 && x4 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s627;
						end
					else if( ~x62 && x16 && ~x15 && ~x4 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else if( ~x62 && ~x16 && x15 && x12 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x62 && ~x16 && x15 && ~x12 )
						nx_state = s61;
					else if( ~x62 && ~x16 && ~x15 && x14 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else if( ~x62 && ~x16 && ~x15 && ~x14 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else nx_state = s61;
				s62 : if( x69 && x15 && x16 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s477;
						end
					else if( x69 && x15 && ~x16 && x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( x69 && x15 && ~x16 && ~x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s477;
						end
					else if( x69 && ~x15 && x16 && x4 && x5 && x1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s477;
						end
					else if( x69 && ~x15 && x16 && x4 && x5 && ~x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s60;
						end
					else if( x69 && ~x15 && x16 && x4 && ~x5 && x1 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( x69 && ~x15 && x16 && x4 && ~x5 && ~x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x69 && ~x15 && x16 && ~x4 && x1 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( x69 && ~x15 && x16 && ~x4 && ~x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x69 && ~x15 && ~x16 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s477;
						end
					else if( ~x69 && x64 && x40 && x13 && x23 && x51 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s507;
						end
					else if( ~x69 && x64 && x40 && x13 && x23 && ~x51 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && x64 && x40 && x13 && ~x23 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s507;
						end
					else if( ~x69 && x64 && x40 && ~x13 && x28 && x35 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s507;
						end
					else if( ~x69 && x64 && x40 && ~x13 && x28 && x35 && ~x5 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x64 && x40 && ~x13 && x28 && ~x35 && x41 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && x64 && x40 && ~x13 && x28 && ~x35 && ~x41 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x64 && x40 && ~x13 && ~x28 && x6 && x35 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s638;
						end
					else if( ~x69 && x64 && x40 && ~x13 && ~x28 && x6 && ~x35 && x41 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && x64 && x40 && ~x13 && ~x28 && x6 && ~x35 && ~x41 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x64 && x40 && ~x13 && ~x28 && ~x6 && x39 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x64 && x40 && ~x13 && ~x28 && ~x6 && ~x39 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x69 && x64 && ~x40 && x11 && x10 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x69 && x64 && ~x40 && x11 && ~x10 && x1 )
						begin
							y3 = 1'b1;	y13 = 1'b1;	y18 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s639;
						end
					else if( ~x69 && x64 && ~x40 && x11 && ~x10 && ~x1 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && x64 && ~x40 && x11 && ~x10 && ~x1 && ~x3 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x69 && x64 && ~x40 && ~x11 && x10 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x64 && ~x40 && ~x11 && ~x10 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && x64 && ~x40 && ~x11 && ~x10 && ~x5 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x69 && ~x64 && x44 && x13 && x23 && x51 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s511;
						end
					else if( ~x69 && ~x64 && x44 && x13 && x23 && ~x51 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else if( ~x69 && ~x64 && x44 && x13 && ~x23 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s511;
						end
					else if( ~x69 && ~x64 && x44 && ~x13 && x28 && x35 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s511;
						end
					else if( ~x69 && ~x64 && x44 && ~x13 && x28 && x35 && ~x5 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && ~x64 && x44 && ~x13 && x28 && ~x35 && x45 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x69 && ~x64 && x44 && ~x13 && x28 && ~x35 && ~x45 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && ~x64 && x44 && ~x13 && ~x28 && x6 && x35 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s638;
						end
					else if( ~x69 && ~x64 && x44 && ~x13 && ~x28 && x6 && ~x35 && x45 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x69 && ~x64 && x44 && ~x13 && ~x28 && x6 && ~x35 && ~x45 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && ~x64 && x44 && ~x13 && ~x28 && ~x6 && x39 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && ~x64 && x44 && ~x13 && ~x28 && ~x6 && ~x39 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x69 && ~x64 && ~x44 && x10 && x11 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x69 && ~x64 && ~x44 && x10 && ~x11 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && ~x64 && ~x44 && ~x10 && x11 && x37 )
						begin
							y3 = 1'b1;	y13 = 1'b1;	y22 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s640;
						end
					else if( ~x69 && ~x64 && ~x44 && ~x10 && x11 && ~x37 && x41 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else if( ~x69 && ~x64 && ~x44 && ~x10 && x11 && ~x37 && ~x41 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x69 && ~x64 && ~x44 && ~x10 && ~x11 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && ~x64 && ~x44 && ~x10 && ~x11 && ~x5 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s631;
						end
					else nx_state = s62;
				s63 : if( x69 && x70 && x63 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s641;
						end
					else if( x69 && x70 && ~x63 && x64 && x65 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x69 && x70 && ~x63 && x64 && x65 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x69 && x70 && ~x63 && x64 && x65 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x63 && x64 && x65 && ~x14 )
						nx_state = s1;
					else if( x69 && x70 && ~x63 && x64 && ~x65 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x63 && x64 && ~x65 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x63 && x64 && ~x65 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x63 && x64 && ~x65 && ~x9 )
						nx_state = s1;
					else if( x69 && x70 && ~x63 && ~x64 && x67 && x11 && x12 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && x70 && ~x63 && ~x64 && x67 && x11 && ~x12 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && x70 && ~x63 && ~x64 && x67 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x69 && x70 && ~x63 && ~x64 && x67 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x63 && ~x64 && ~x67 && x28 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x63 && ~x64 && ~x67 && x28 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x63 && ~x64 && ~x67 && x28 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x69 && x70 && ~x63 && ~x64 && ~x67 && x28 && ~x23 )
						nx_state = s1;
					else if( x69 && x70 && ~x63 && ~x64 && ~x67 && ~x28 )
						begin
							y8 = 1'b1;	
							nx_state = s642;
						end
					else if( x69 && ~x70 && x67 && x65 && x21 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x69 && ~x70 && x67 && x65 && x21 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x69 && ~x70 && x67 && x65 && x21 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x65 && x21 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x65 && ~x21 && x23 && x22 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x67 && x65 && ~x21 && x23 && x22 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x67 && x65 && ~x21 && x23 && x22 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x65 && ~x21 && x23 && x22 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x65 && ~x21 && x23 && ~x22 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x67 && x65 && ~x21 && x23 && ~x22 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x67 && x65 && ~x21 && x23 && ~x22 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x65 && ~x21 && x23 && ~x22 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x65 && ~x21 && ~x23 && x8 && x22 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x67 && x65 && ~x21 && ~x23 && x8 && x22 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x67 && x65 && ~x21 && ~x23 && x8 && x22 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x65 && ~x21 && ~x23 && x8 && ~x22 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x67 && x65 && ~x21 && ~x23 && x8 && ~x22 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x67 && x65 && ~x21 && ~x23 && x8 && ~x22 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && x65 && ~x21 && ~x23 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x65 && x66 && x68 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x70 && x67 && ~x65 && x66 && x68 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x70 && x67 && ~x65 && x66 && x68 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x65 && x66 && x68 && x21 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x65 && x66 && x68 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( x69 && ~x70 && x67 && ~x65 && x66 && x68 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( x69 && ~x70 && x67 && ~x65 && x66 && x68 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x65 && x66 && x68 && ~x21 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x65 && x66 && ~x68 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x65 && ~x66 && x24 && x26 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s430;
						end
					else if( x69 && ~x70 && x67 && ~x65 && ~x66 && x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( x69 && ~x70 && x67 && ~x65 && ~x66 && x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( x69 && ~x70 && x67 && ~x65 && ~x66 && x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x65 && ~x66 && x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x65 && ~x66 && ~x24 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && x67 && ~x65 && ~x66 && ~x24 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && x67 && ~x65 && ~x66 && ~x24 && x25 && x19 && ~x14 && ~x13 && x26 )
						nx_state = s63;
					else if( x69 && ~x70 && x67 && ~x65 && ~x66 && ~x24 && x25 && x19 && ~x14 && ~x13 && ~x26 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x65 && ~x66 && ~x24 && x25 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x65 && ~x66 && ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && x67 && ~x65 && ~x66 && ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && x67 && ~x65 && ~x66 && ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x65 && ~x66 && ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x65 && ~x66 && ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && x67 && ~x65 && ~x66 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && x67 && ~x65 && ~x66 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x67 && ~x65 && ~x66 && ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x65 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x67 && x65 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x67 && x65 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x67 && x65 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x65 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x65 && ~x21 && x23 && x22 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( x69 && ~x70 && ~x67 && x65 && ~x21 && x23 && x22 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && ~x67 && x65 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && ~x67 && x65 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x65 && ~x21 && x23 && x22 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x65 && ~x21 && x23 && ~x22 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && ~x67 && x65 && ~x21 && x23 && ~x22 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && ~x67 && x65 && ~x21 && x23 && ~x22 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x65 && ~x21 && x23 && ~x22 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x65 && ~x21 && ~x23 && x18 && x14 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && ~x67 && x65 && ~x21 && ~x23 && x18 && x14 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && ~x67 && x65 && ~x21 && ~x23 && x18 && ~x14 && x13 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && ~x67 && x65 && ~x21 && ~x23 && x18 && ~x14 && x13 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && ~x67 && x65 && ~x21 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && x65 && ~x21 && ~x23 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x65 && x21 && x66 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && ~x67 && ~x65 && x21 && x66 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && ~x67 && ~x65 && x21 && x66 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x65 && x21 && x66 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x65 && x21 && ~x66 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x69 && ~x70 && ~x67 && ~x65 && x21 && ~x66 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x69 && ~x70 && ~x67 && ~x65 && x21 && ~x66 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x65 && x21 && ~x66 && ~x3 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x65 && ~x21 && x22 && x66 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && ~x70 && ~x67 && ~x65 && ~x21 && x22 && ~x66 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && ~x67 && ~x65 && ~x21 && ~x22 && x66 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && ~x67 && ~x65 && ~x21 && ~x22 && x66 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && ~x67 && ~x65 && ~x21 && ~x22 && x66 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x65 && ~x21 && ~x22 && x66 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x65 && ~x21 && ~x22 && ~x66 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( x69 && ~x70 && ~x67 && ~x65 && ~x21 && ~x22 && ~x66 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( x69 && ~x70 && ~x67 && ~x65 && ~x21 && ~x22 && ~x66 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x67 && ~x65 && ~x21 && ~x22 && ~x66 && ~x8 )
						nx_state = s1;
					else if( ~x69 && x70 && x1 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s644;
						end
					else if( ~x69 && x70 && ~x1 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x69 && ~x70 && x45 && x12 && x1 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x69 && ~x70 && x45 && x12 && ~x1 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x69 && ~x70 && x45 && ~x12 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x45 && x11 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x45 && ~x11 && x46 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x45 && ~x11 && ~x46 && x1 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x11 && ~x46 && ~x1 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else nx_state = s63;
				s64 : if( x62 && x64 )
						begin
							y1 = 1'b1;	y12 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s382;
						end
					else if( x62 && ~x64 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y37 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x62 && x63 && x67 && x11 && x14 && x13 && x1 )
						begin
							y5 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x62 && x63 && x67 && x11 && x14 && x13 && ~x1 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( ~x62 && x63 && x67 && x11 && x14 && ~x13 && x4 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y4 = 1'b1;	
							nx_state = s71;
						end
					else if( ~x62 && x63 && x67 && x11 && x14 && ~x13 && x4 && ~x2 )
						nx_state = s64;
					else if( ~x62 && x63 && x67 && x11 && x14 && ~x13 && ~x4 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s68;
						end
					else if( ~x62 && x63 && x67 && x11 && x14 && ~x13 && ~x4 && ~x2 )
						nx_state = s64;
					else if( ~x62 && x63 && x67 && x11 && ~x14 && x4 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y4 = 1'b1;	
							nx_state = s71;
						end
					else if( ~x62 && x63 && x67 && x11 && ~x14 && x4 && ~x2 )
						nx_state = s64;
					else if( ~x62 && x63 && x67 && x11 && ~x14 && ~x4 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s68;
						end
					else if( ~x62 && x63 && x67 && x11 && ~x14 && ~x4 && ~x2 )
						nx_state = s64;
					else if( ~x62 && x63 && x67 && ~x11 && x10 && x13 )
						nx_state = s1;
					else if( ~x62 && x63 && x67 && ~x11 && x10 && ~x13 && x4 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y4 = 1'b1;	
							nx_state = s71;
						end
					else if( ~x62 && x63 && x67 && ~x11 && x10 && ~x13 && x4 && ~x2 )
						nx_state = s64;
					else if( ~x62 && x63 && x67 && ~x11 && x10 && ~x13 && ~x4 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s68;
						end
					else if( ~x62 && x63 && x67 && ~x11 && x10 && ~x13 && ~x4 && ~x2 )
						nx_state = s64;
					else if( ~x62 && x63 && x67 && ~x11 && ~x10 && x4 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y4 = 1'b1;	
							nx_state = s71;
						end
					else if( ~x62 && x63 && x67 && ~x11 && ~x10 && x4 && ~x2 )
						nx_state = s64;
					else if( ~x62 && x63 && x67 && ~x11 && ~x10 && ~x4 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s68;
						end
					else if( ~x62 && x63 && x67 && ~x11 && ~x10 && ~x4 && ~x2 )
						nx_state = s64;
					else if( ~x62 && x63 && ~x67 && x13 && x10 )
						nx_state = s1;
					else if( ~x62 && x63 && ~x67 && x13 && ~x10 && x15 && x14 && x1 )
						begin
							y5 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x62 && x63 && ~x67 && x13 && ~x10 && x15 && x14 && ~x1 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( ~x62 && x63 && ~x67 && x13 && ~x10 && x15 && ~x14 && x4 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y4 = 1'b1;	
							nx_state = s71;
						end
					else if( ~x62 && x63 && ~x67 && x13 && ~x10 && x15 && ~x14 && x4 && ~x2 )
						nx_state = s64;
					else if( ~x62 && x63 && ~x67 && x13 && ~x10 && x15 && ~x14 && ~x4 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s68;
						end
					else if( ~x62 && x63 && ~x67 && x13 && ~x10 && x15 && ~x14 && ~x4 && ~x2 )
						nx_state = s64;
					else if( ~x62 && x63 && ~x67 && x13 && ~x10 && ~x15 && x11 )
						nx_state = s1;
					else if( ~x62 && x63 && ~x67 && x13 && ~x10 && ~x15 && ~x11 && x4 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y4 = 1'b1;	
							nx_state = s71;
						end
					else if( ~x62 && x63 && ~x67 && x13 && ~x10 && ~x15 && ~x11 && x4 && ~x2 )
						nx_state = s64;
					else if( ~x62 && x63 && ~x67 && x13 && ~x10 && ~x15 && ~x11 && ~x4 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s68;
						end
					else if( ~x62 && x63 && ~x67 && x13 && ~x10 && ~x15 && ~x11 && ~x4 && ~x2 )
						nx_state = s64;
					else if( ~x62 && x63 && ~x67 && ~x13 && x4 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y4 = 1'b1;	
							nx_state = s71;
						end
					else if( ~x62 && x63 && ~x67 && ~x13 && x4 && ~x2 )
						nx_state = s64;
					else if( ~x62 && x63 && ~x67 && ~x13 && ~x4 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s68;
						end
					else if( ~x62 && x63 && ~x67 && ~x13 && ~x4 && ~x2 )
						nx_state = s64;
					else if( ~x62 && ~x63 )
						begin
							y12 = 1'b1;	y48 = 1'b1;	
							nx_state = s646;
						end
					else nx_state = s64;
				s65 : if( x13 && x67 && x14 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x13 && x67 && ~x14 && x11 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x13 && x67 && ~x14 && ~x11 && x10 && x6 && x2 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s577;
						end
					else if( x13 && x67 && ~x14 && ~x11 && x10 && x6 && ~x2 )
						nx_state = s65;
					else if( x13 && x67 && ~x14 && ~x11 && x10 && ~x6 && x2 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x13 && x67 && ~x14 && ~x11 && x10 && ~x6 && ~x2 )
						nx_state = s65;
					else if( x13 && x67 && ~x14 && ~x11 && ~x10 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x13 && ~x67 && x15 && x14 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x13 && ~x67 && x15 && ~x14 && x10 && x6 && x2 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s577;
						end
					else if( x13 && ~x67 && x15 && ~x14 && x10 && x6 && ~x2 )
						nx_state = s65;
					else if( x13 && ~x67 && x15 && ~x14 && x10 && ~x6 && x2 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x13 && ~x67 && x15 && ~x14 && x10 && ~x6 && ~x2 )
						nx_state = s65;
					else if( x13 && ~x67 && x15 && ~x14 && ~x10 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x13 && ~x67 && ~x15 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x13 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else nx_state = s65;
				s66 : if( x70 && x62 && x64 )
						begin
							y1 = 1'b1;	y12 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s647;
						end
					else if( x70 && x62 && ~x64 )
						begin
							y27 = 1'b1;	
							nx_state = s648;
						end
					else if( x70 && ~x62 && x63 && x67 && x14 && x13 && x11 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( x70 && ~x62 && x63 && x67 && x14 && x13 && ~x11 && x10 && x4 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && ~x62 && x63 && x67 && x14 && x13 && ~x11 && x10 && ~x4 )
						nx_state = s66;
					else if( x70 && ~x62 && x63 && x67 && x14 && x13 && ~x11 && ~x10 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && ~x62 && x63 && x67 && x14 && x13 && ~x11 && ~x10 && ~x3 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s68;
						end
					else if( x70 && ~x62 && x63 && x67 && x14 && x13 && ~x11 && ~x10 && ~x3 && ~x2 )
						nx_state = s66;
					else if( x70 && ~x62 && x63 && x67 && x14 && ~x13 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && ~x62 && x63 && x67 && x14 && ~x13 && ~x3 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s68;
						end
					else if( x70 && ~x62 && x63 && x67 && x14 && ~x13 && ~x3 && ~x2 )
						nx_state = s66;
					else if( x70 && ~x62 && x63 && x67 && ~x14 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && ~x62 && x63 && x67 && ~x14 && ~x3 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s68;
						end
					else if( x70 && ~x62 && x63 && x67 && ~x14 && ~x3 && ~x2 )
						nx_state = s66;
					else if( x70 && ~x62 && x63 && ~x67 && x15 && x13 && x14 && x10 && x4 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && ~x62 && x63 && ~x67 && x15 && x13 && x14 && x10 && ~x4 )
						nx_state = s66;
					else if( x70 && ~x62 && x63 && ~x67 && x15 && x13 && x14 && ~x10 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( x70 && ~x62 && x63 && ~x67 && x15 && x13 && ~x14 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && ~x62 && x63 && ~x67 && x15 && x13 && ~x14 && ~x3 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s68;
						end
					else if( x70 && ~x62 && x63 && ~x67 && x15 && x13 && ~x14 && ~x3 && ~x2 )
						nx_state = s66;
					else if( x70 && ~x62 && x63 && ~x67 && x15 && ~x13 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && ~x62 && x63 && ~x67 && x15 && ~x13 && ~x3 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s68;
						end
					else if( x70 && ~x62 && x63 && ~x67 && x15 && ~x13 && ~x3 && ~x2 )
						nx_state = s66;
					else if( x70 && ~x62 && x63 && ~x67 && ~x15 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x15 && ~x3 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s68;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x15 && ~x3 && ~x2 )
						nx_state = s66;
					else if( x70 && ~x62 && ~x63 && x64 && x21 )
						begin
							y6 = 1'b1;	
							nx_state = s649;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x21 )
						begin
							y6 = 1'b1;	
							nx_state = s368;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 )
						begin
							y33 = 1'b1;	
							nx_state = s589;
						end
					else if( ~x70 && x66 && x21 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x70 && x66 && ~x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && ~x66 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s377;
						end
					else nx_state = s66;
				s67 : if( x70 && x13 && x67 && x11 && x14 )
						nx_state = s1;
					else if( x70 && x13 && x67 && x11 && ~x14 )
						begin
							y5 = 1'b1;	
							nx_state = s66;
						end
					else if( x70 && x13 && x67 && ~x11 && x10 && x4 && x3 && x14 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( x70 && x13 && x67 && ~x11 && x10 && x4 && x3 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s68;
						end
					else if( x70 && x13 && x67 && ~x11 && x10 && x4 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && x13 && x67 && ~x11 && x10 && ~x4 )
						nx_state = s67;
					else if( x70 && x13 && x67 && ~x11 && ~x10 )
						nx_state = s1;
					else if( x70 && x13 && ~x67 && x15 && x10 && x4 && x3 && x14 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( x70 && x13 && ~x67 && x15 && x10 && x4 && x3 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s68;
						end
					else if( x70 && x13 && ~x67 && x15 && x10 && x4 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && x13 && ~x67 && x15 && x10 && ~x4 )
						nx_state = s67;
					else if( x70 && x13 && ~x67 && x15 && ~x10 && x14 )
						nx_state = s1;
					else if( x70 && x13 && ~x67 && x15 && ~x10 && ~x14 )
						begin
							y5 = 1'b1;	
							nx_state = s66;
						end
					else if( x70 && x13 && ~x67 && ~x15 && x11 && x4 && x14 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && x13 && ~x67 && ~x15 && x11 && x4 && ~x14 && x3 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s132;
						end
					else if( x70 && x13 && ~x67 && ~x15 && x11 && x4 && ~x14 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && x13 && ~x67 && ~x15 && x11 && ~x4 )
						nx_state = s67;
					else if( x70 && x13 && ~x67 && ~x15 && ~x11 && x10 && x4 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && x13 && ~x67 && ~x15 && ~x11 && x10 && ~x4 )
						nx_state = s67;
					else if( x70 && x13 && ~x67 && ~x15 && ~x11 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x13 )
						begin
							y5 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x70 && x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x23 && x15 && x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && ~x21 && x23 && x15 && ~x10 && x12 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && ~x21 && x23 && x15 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s366;
						end
					else if( ~x70 && ~x21 && x23 && ~x15 && x16 && x10 && x12 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else if( ~x70 && ~x21 && x23 && ~x15 && x16 && x10 && ~x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x70 && ~x21 && x23 && ~x15 && x16 && ~x10 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else if( ~x70 && ~x21 && x23 && ~x15 && ~x16 )
						nx_state = s47;
					else if( ~x70 && ~x21 && ~x23 && x15 && x10 && x11 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x70 && ~x21 && ~x23 && x15 && x10 && ~x11 && x12 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x70 && ~x21 && ~x23 && x15 && x10 && ~x11 && ~x12 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && ~x21 && ~x23 && x15 && ~x10 && x12 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( ~x70 && ~x21 && ~x23 && x15 && ~x10 && x12 && ~x11 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && ~x21 && ~x23 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( ~x70 && ~x21 && ~x23 && ~x15 && x16 && x10 && x12 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x21 && ~x23 && ~x15 && x16 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s365;
						end
					else if( ~x70 && ~x21 && ~x23 && ~x15 && x16 && ~x10 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x21 && ~x23 && ~x15 && ~x16 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s151;
						end
					else nx_state = s67;
				s68 : if( x67 && x11 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( x67 && ~x11 && x13 && x14 && x10 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( x67 && ~x11 && x13 && x14 && ~x10 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y4 = 1'b1;	
							nx_state = s71;
						end
					else if( x67 && ~x11 && x13 && x14 && ~x10 && ~x1 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x67 && ~x11 && x13 && x14 && ~x10 && ~x1 && ~x2 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x67 && ~x11 && x13 && ~x14 && x10 && x6 && x2 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s577;
						end
					else if( x67 && ~x11 && x13 && ~x14 && x10 && x6 && ~x2 )
						nx_state = s68;
					else if( x67 && ~x11 && x13 && ~x14 && x10 && ~x6 && x2 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x67 && ~x11 && x13 && ~x14 && x10 && ~x6 && ~x2 )
						nx_state = s68;
					else if( x67 && ~x11 && x13 && ~x14 && ~x10 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( x67 && ~x11 && ~x13 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( ~x67 && x10 && x13 && x14 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( ~x67 && x10 && x13 && ~x14 && x15 && x6 && x2 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s577;
						end
					else if( ~x67 && x10 && x13 && ~x14 && x15 && x6 && ~x2 )
						nx_state = s68;
					else if( ~x67 && x10 && x13 && ~x14 && x15 && ~x6 && x2 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x67 && x10 && x13 && ~x14 && x15 && ~x6 && ~x2 )
						nx_state = s68;
					else if( ~x67 && x10 && x13 && ~x14 && ~x15 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( ~x67 && x10 && ~x13 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( ~x67 && ~x10 && x11 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( ~x67 && ~x10 && ~x11 && x13 && x14 && x15 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( ~x67 && ~x10 && ~x11 && x13 && x14 && ~x15 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y4 = 1'b1;	
							nx_state = s71;
						end
					else if( ~x67 && ~x10 && ~x11 && x13 && x14 && ~x15 && ~x1 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( ~x67 && ~x10 && ~x11 && x13 && x14 && ~x15 && ~x1 && ~x2 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x67 && ~x10 && ~x11 && x13 && ~x14 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( ~x67 && ~x10 && ~x11 && ~x13 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else nx_state = s68;
				s69 : if( x13 && x67 && x11 && x14 && x8 && x1 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x13 && x67 && x11 && x14 && x8 && ~x1 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x13 && x67 && x11 && x14 && ~x8 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x13 && x67 && x11 && ~x14 )
						begin
							y5 = 1'b1;	
							nx_state = s64;
						end
					else if( x13 && x67 && ~x11 && x10 && x14 && x3 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s66;
						end
					else if( x13 && x67 && ~x11 && x10 && x14 && x3 && ~x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x13 && x67 && ~x11 && x10 && x14 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x13 && x67 && ~x11 && x10 && ~x14 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s65;
						end
					else if( x13 && x67 && ~x11 && x10 && ~x14 && ~x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x13 && x67 && ~x11 && ~x10 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x13 && x67 && ~x11 && ~x10 && ~x1 && x3 )
						nx_state = s1;
					else if( x13 && x67 && ~x11 && ~x10 && ~x1 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x13 && ~x67 && x15 && x10 && x14 && x3 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s66;
						end
					else if( x13 && ~x67 && x15 && x10 && x14 && x3 && ~x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x13 && ~x67 && x15 && x10 && x14 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x13 && ~x67 && x15 && x10 && ~x14 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s65;
						end
					else if( x13 && ~x67 && x15 && x10 && ~x14 && ~x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x13 && ~x67 && x15 && ~x10 && x14 && x8 && x1 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x13 && ~x67 && x15 && ~x10 && x14 && x8 && ~x1 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x13 && ~x67 && x15 && ~x10 && x14 && ~x8 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x13 && ~x67 && x15 && ~x10 && ~x14 )
						begin
							y5 = 1'b1;	
							nx_state = s64;
						end
					else if( x13 && ~x67 && ~x15 && x11 && x5 && x14 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x13 && ~x67 && ~x15 && x11 && x5 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x13 && ~x67 && ~x15 && x11 && ~x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x13 && ~x67 && ~x15 && ~x11 && x10 && x5 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x13 && ~x67 && ~x15 && ~x11 && x10 && ~x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x13 && ~x67 && ~x15 && ~x11 && ~x10 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x13 && ~x67 && ~x15 && ~x11 && ~x10 && ~x1 && x3 )
						nx_state = s1;
					else if( x13 && ~x67 && ~x15 && ~x11 && ~x10 && ~x1 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( ~x13 )
						begin
							y5 = 1'b1;	
							nx_state = s64;
						end
					else nx_state = s69;
				s70 : if( x69 && x70 && x67 && x3 )
						nx_state = s1;
					else if( x69 && x70 && x67 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x69 && x70 && ~x67 && x11 && x14 && x3 )
						nx_state = s1;
					else if( x69 && x70 && ~x67 && x11 && x14 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x69 && x70 && ~x67 && x11 && ~x14 && x2 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( x69 && x70 && ~x67 && x11 && ~x14 && ~x2 )
						nx_state = s70;
					else if( x69 && x70 && ~x67 && ~x11 && x3 )
						nx_state = s1;
					else if( x69 && x70 && ~x67 && ~x11 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x69 && ~x70 && x65 && x66 && x61 && x60 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x66 && x61 && ~x60 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x65 && x66 && x61 && ~x60 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x65 && x66 && x61 && ~x60 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x66 && x61 && ~x60 && x62 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x66 && x61 && ~x60 && ~x62 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x61 && x60 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x61 && ~x60 && x62 && x7 && x15 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s491;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x61 && ~x60 && x62 && x7 && x15 && ~x12 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s135;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x61 && ~x60 && x62 && x7 && ~x15 && x16 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s490;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x61 && ~x60 && x62 && x7 && ~x15 && x16 && ~x12 && x2 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s269;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x61 && ~x60 && x62 && x7 && ~x15 && x16 && ~x12 && ~x2 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s565;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x61 && ~x60 && x62 && x7 && ~x15 && ~x16 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x61 && ~x60 && x62 && ~x7 && x15 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s490;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x61 && ~x60 && x62 && ~x7 && x15 && ~x12 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s566;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x61 && ~x60 && x62 && ~x7 && ~x15 && x16 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x61 && ~x60 && x62 && ~x7 && ~x15 && ~x16 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x61 && ~x60 && ~x62 && x4 && x15 && x7 )
						nx_state = s47;
					else if( x69 && ~x70 && x65 && x66 && ~x61 && ~x60 && ~x62 && x4 && x15 && ~x7 && x11 )
						nx_state = s47;
					else if( x69 && ~x70 && x65 && x66 && ~x61 && ~x60 && ~x62 && x4 && x15 && ~x7 && ~x11 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x61 && ~x60 && ~x62 && x4 && ~x15 && x16 )
						nx_state = s141;
					else if( x69 && ~x70 && x65 && x66 && ~x61 && ~x60 && ~x62 && x4 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x61 && ~x60 && ~x62 && ~x4 )
						nx_state = s141;
					else if( x69 && ~x70 && x65 && ~x66 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( x69 && ~x70 && ~x65 && x21 && x66 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && ~x65 && x21 && x66 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && ~x65 && x21 && x66 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x21 && x66 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x21 && ~x66 && x19 && x20 && x12 && x17 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	
							nx_state = s569;
						end
					else if( x69 && ~x70 && ~x65 && x21 && ~x66 && x19 && x20 && x12 && ~x17 )
						begin
							y8 = 1'b1;	y22 = 1'b1;	
							nx_state = s570;
						end
					else if( x69 && ~x70 && ~x65 && x21 && ~x66 && x19 && x20 && ~x12 && x16 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x65 && x21 && ~x66 && x19 && x20 && ~x12 && ~x16 && x17 && x5 )
						begin
							y8 = 1'b1;	
							nx_state = s373;
						end
					else if( x69 && ~x70 && ~x65 && x21 && ~x66 && x19 && x20 && ~x12 && ~x16 && x17 && ~x5 )
						begin
							y8 = 1'b1;	
							nx_state = s568;
						end
					else if( x69 && ~x70 && ~x65 && x21 && ~x66 && x19 && x20 && ~x12 && ~x16 && ~x17 && x4 )
						begin
							y8 = 1'b1;	
							nx_state = s373;
						end
					else if( x69 && ~x70 && ~x65 && x21 && ~x66 && x19 && x20 && ~x12 && ~x16 && ~x17 && ~x4 )
						begin
							y8 = 1'b1;	
							nx_state = s568;
						end
					else if( x69 && ~x70 && ~x65 && x21 && ~x66 && x19 && ~x20 && x16 && x12 )
						begin
							y8 = 1'b1;	y18 = 1'b1;	
							nx_state = s650;
						end
					else if( x69 && ~x70 && ~x65 && x21 && ~x66 && x19 && ~x20 && x16 && ~x12 && x17 )
						begin
							y8 = 1'b1;	y18 = 1'b1;	
							nx_state = s152;
						end
					else if( x69 && ~x70 && ~x65 && x21 && ~x66 && x19 && ~x20 && x16 && ~x12 && ~x17 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x65 && x21 && ~x66 && x19 && ~x20 && ~x16 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x65 && x21 && ~x66 && ~x19 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x65 && ~x21 && x66 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && ~x21 && ~x66 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && x2 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x69 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else nx_state = s70;
				s71 : if( x64 && x65 && x4 && x5 && x3 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x64 && x65 && x4 && x5 && ~x3 && x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s651;
						end
					else if( x64 && x65 && x4 && x5 && ~x3 && ~x6 && x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s651;
						end
					else if( x64 && x65 && x4 && x5 && ~x3 && ~x6 && ~x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s652;
						end
					else if( x64 && x65 && x4 && ~x5 && x3 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( x64 && x65 && x4 && ~x5 && ~x3 && x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s653;
						end
					else if( x64 && x65 && x4 && ~x5 && ~x3 && ~x6 && x7 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s653;
						end
					else if( x64 && x65 && x4 && ~x5 && ~x3 && ~x6 && ~x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s654;
						end
					else if( x64 && x65 && ~x4 && x5 && x3 )
						begin
							y51 = 1'b1;	
							nx_state = s655;
						end
					else if( x64 && x65 && ~x4 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s654;
						end
					else if( x64 && x65 && ~x4 && ~x5 && x3 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y48 = 1'b1;	
							y50 = 1'b1;	
							nx_state = s654;
						end
					else if( x64 && x65 && ~x4 && ~x5 && ~x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s654;
						end
					else if( x64 && ~x65 && x13 && x10 && x67 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x64 && ~x65 && x13 && x10 && ~x67 && x2 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x64 && ~x65 && x13 && x10 && ~x67 && ~x2 && x15 )
						nx_state = s71;
					else if( x64 && ~x65 && x13 && x10 && ~x67 && ~x2 && ~x15 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x64 && ~x65 && x13 && ~x10 && x11 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x64 && ~x65 && x13 && ~x10 && ~x11 && x67 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x64 && ~x65 && x13 && ~x10 && ~x11 && x67 && ~x2 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x64 && ~x65 && x13 && ~x10 && ~x11 && ~x67 && x15 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x64 && ~x65 && x13 && ~x10 && ~x11 && ~x67 && ~x15 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x64 && ~x65 && x13 && ~x10 && ~x11 && ~x67 && ~x15 && ~x2 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x64 && ~x65 && ~x13 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x64 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s656;
						end
					else nx_state = s71;
				s72 : if( x22 && x23 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x22 && ~x23 && x16 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x22 && ~x23 && x16 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x22 && ~x23 && x16 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x22 && ~x23 && x16 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x22 && ~x23 && x16 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x22 && ~x23 && ~x16 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s657;
						end
					else if( ~x22 && x23 && x16 )
						begin
							y50 = 1'b1;	
							nx_state = s658;
						end
					else if( ~x22 && x23 && ~x16 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s657;
						end
					else if( ~x22 && ~x23 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else nx_state = s72;
				s73 : if( x22 )
						begin
							y6 = 1'b1;	
							nx_state = s659;
						end
					else if( ~x22 )
						begin
							y6 = 1'b1;	
							nx_state = s431;
						end
					else nx_state = s73;
				s74 : if( 1'b1 )
						begin
							y37 = 1'b1;	y38 = 1'b1;	
							nx_state = s660;
						end
					else nx_state = s74;
				s75 : if( x70 && x62 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s661;
						end
					else if( x70 && ~x62 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s662;
						end
					else if( ~x70 && x65 && x21 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s663;
						end
					else if( ~x70 && x65 && ~x21 && x22 && x23 && x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( ~x70 && x65 && ~x21 && x22 && x23 && ~x15 && x19 && x18 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( ~x70 && x65 && ~x21 && x22 && x23 && ~x15 && x19 && ~x18 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s461;
						end
					else if( ~x70 && x65 && ~x21 && x22 && x23 && ~x15 && ~x19 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( ~x70 && x65 && ~x21 && x22 && ~x23 && x11 && x18 && x15 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x70 && x65 && ~x21 && x22 && ~x23 && x11 && x18 && ~x15 )
						begin
							y15 = 1'b1;	y20 = 1'b1;	
							nx_state = s665;
						end
					else if( ~x70 && x65 && ~x21 && x22 && ~x23 && x11 && ~x18 && x19 && x15 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s666;
						end
					else if( ~x70 && x65 && ~x21 && x22 && ~x23 && x11 && ~x18 && x19 && ~x15 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x70 && x65 && ~x21 && x22 && ~x23 && x11 && ~x18 && ~x19 )
						begin
							y12 = 1'b1;	
							nx_state = s245;
						end
					else if( ~x70 && x65 && ~x21 && x22 && ~x23 && ~x11 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x70 && x65 && ~x21 && ~x22 && x23 && x16 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( ~x70 && x65 && ~x21 && ~x22 && x23 && ~x16 && x20 && x19 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( ~x70 && x65 && ~x21 && ~x22 && x23 && ~x16 && x20 && ~x19 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && ~x22 && x23 && ~x16 && x20 && ~x19 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && ~x22 && x23 && ~x16 && x20 && ~x19 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && ~x22 && x23 && ~x16 && x20 && ~x19 && ~x9 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && ~x22 && x23 && ~x16 && ~x20 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( ~x70 && x65 && ~x21 && ~x22 && ~x23 && x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( ~x70 && x65 && ~x21 && ~x22 && ~x23 && ~x15 && x19 && x18 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( ~x70 && x65 && ~x21 && ~x22 && ~x23 && ~x15 && x19 && ~x18 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s461;
						end
					else if( ~x70 && x65 && ~x21 && ~x22 && ~x23 && ~x15 && ~x19 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( ~x70 && ~x65 && x24 && x16 && x26 && x11 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s309;
						end
					else if( ~x70 && ~x65 && x24 && x16 && x26 && ~x11 && x7 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x65 && x24 && x16 && x26 && ~x11 && ~x7 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s309;
						end
					else if( ~x70 && ~x65 && x24 && x16 && ~x26 && x6 && x11 && x12 )
						begin
							y11 = 1'b1;	
							nx_state = s272;
						end
					else if( ~x70 && ~x65 && x24 && x16 && ~x26 && x6 && x11 && ~x12 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x70 && ~x65 && x24 && x16 && ~x26 && x6 && x11 && ~x12 && ~x13 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s300;
						end
					else if( ~x70 && ~x65 && x24 && x16 && ~x26 && x6 && ~x11 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && ~x65 && x24 && x16 && ~x26 && ~x6 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && x26 && x7 && x17 && x13 && x11 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && x26 && x7 && x17 && x13 && ~x11 && x12 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && x26 && x7 && x17 && x13 && ~x11 && ~x12 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && x26 && x7 && x17 && ~x13 && x11 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s430;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && x26 && x7 && x17 && ~x13 && ~x11 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && x26 && x7 && ~x17 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && x26 && ~x7 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s309;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && x11 && x9 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && x11 && ~x9 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && x11 && ~x9 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && x11 && ~x9 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && x11 && ~x9 && ~x20 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && ~x11 && x7 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && ~x11 && ~x7 && x12 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && ~x11 && ~x7 && ~x12 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && ~x11 && ~x7 && ~x12 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && ~x11 && ~x7 && ~x12 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && ~x11 && ~x7 && ~x12 && ~x20 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && x11 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && ~x11 && x12 && x10 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && ~x11 && x12 && ~x10 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && ~x11 && x12 && ~x10 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && ~x11 && x12 && ~x10 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && ~x11 && x12 && ~x10 && ~x20 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && ~x11 && ~x12 && x8 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && ~x11 && ~x12 && ~x8 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && ~x11 && ~x12 && ~x8 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && ~x11 && ~x12 && ~x8 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && ~x11 && ~x12 && ~x8 && ~x20 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && ~x17 && x6 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x65 && x24 && ~x16 && ~x26 && ~x17 && ~x6 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && ~x65 && ~x24 && x25 && x26 && x1 )
						begin
							y8 = 1'b1;	y17 = 1'b1;	y23 = 1'b1;	
							nx_state = s303;
						end
					else if( ~x70 && ~x65 && ~x24 && x25 && x26 && ~x1 && x18 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x24 && x25 && x26 && ~x1 && ~x18 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && ~x65 && ~x24 && x25 && ~x26 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( ~x70 && ~x65 && ~x24 && x25 && ~x26 && ~x2 && x18 && x15 && x10 && x11 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s433;
						end
					else if( ~x70 && ~x65 && ~x24 && x25 && ~x26 && ~x2 && x18 && x15 && x10 && ~x11 && x12 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s432;
						end
					else if( ~x70 && ~x65 && ~x24 && x25 && ~x26 && ~x2 && x18 && x15 && x10 && ~x11 && ~x12 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s300;
						end
					else if( ~x70 && ~x65 && ~x24 && x25 && ~x26 && ~x2 && x18 && x15 && ~x10 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s126;
						end
					else if( ~x70 && ~x65 && ~x24 && x25 && ~x26 && ~x2 && x18 && ~x15 && x16 && x10 && x12 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x70 && ~x65 && ~x24 && x25 && ~x26 && ~x2 && x18 && ~x15 && x16 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x70 && ~x65 && ~x24 && x25 && ~x26 && ~x2 && x18 && ~x15 && x16 && ~x10 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x70 && ~x65 && ~x24 && x25 && ~x26 && ~x2 && x18 && ~x15 && ~x16 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( ~x70 && ~x65 && ~x24 && x25 && ~x26 && ~x2 && ~x18 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && ~x65 && ~x24 && ~x25 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else nx_state = s75;
				s76 : if( x70 && x21 && x20 )
						begin
							y15 = 1'b1;	y59 = 1'b1;	
							nx_state = s667;
						end
					else if( x70 && x21 && ~x20 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x70 && ~x21 && x20 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x70 && ~x21 && ~x20 )
						begin
							y5 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x70 && x20 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s668;
						end
					else if( ~x70 && ~x20 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else nx_state = s76;
				s77 : if( x69 && x70 && x62 && x64 && x9 && x32 && x33 )
						begin
							y6 = 1'b1;	y40 = 1'b1;	y41 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s346;
						end
					else if( x69 && x70 && x62 && x64 && x9 && x32 && ~x33 && x14 && x15 && x13 )
						begin
							y6 = 1'b1;	y35 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s338;
						end
					else if( x69 && x70 && x62 && x64 && x9 && x32 && ~x33 && x14 && x15 && ~x13 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s352;
						end
					else if( x69 && x70 && x62 && x64 && x9 && x32 && ~x33 && x14 && ~x15 && x13 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s349;
						end
					else if( x69 && x70 && x62 && x64 && x9 && x32 && ~x33 && x14 && ~x15 && ~x13 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s354;
						end
					else if( x69 && x70 && x62 && x64 && x9 && x32 && ~x33 && ~x14 && x15 && x13 && x16 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s347;
						end
					else if( x69 && x70 && x62 && x64 && x9 && x32 && ~x33 && ~x14 && x15 && x13 && ~x16 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s348;
						end
					else if( x69 && x70 && x62 && x64 && x9 && x32 && ~x33 && ~x14 && x15 && ~x13 && x17 )
						nx_state = s1;
					else if( x69 && x70 && x62 && x64 && x9 && x32 && ~x33 && ~x14 && x15 && ~x13 && ~x17 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s353;
						end
					else if( x69 && x70 && x62 && x64 && x9 && x32 && ~x33 && ~x14 && ~x15 && x13 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s350;
						end
					else if( x69 && x70 && x62 && x64 && x9 && x32 && ~x33 && ~x14 && ~x15 && ~x13 && x18 )
						nx_state = s1;
					else if( x69 && x70 && x62 && x64 && x9 && x32 && ~x33 && ~x14 && ~x15 && ~x13 && ~x18 )
						nx_state = s77;
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && x13 && x33 && x15 && x14 && x5 )
						begin
							y6 = 1'b1;	y35 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s338;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && x13 && x33 && x15 && x14 && ~x5 && x7 )
						begin
							y6 = 1'b1;	y35 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s338;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && x13 && x33 && x15 && x14 && ~x5 && ~x7 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y27 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s339;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && x13 && x33 && x15 && ~x14 && x31 && x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s340;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && x13 && x33 && x15 && ~x14 && x31 && ~x5 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && x13 && x33 && x15 && ~x14 && ~x31 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && x13 && x33 && x15 && ~x14 && ~x31 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && x13 && x33 && x15 && ~x14 && ~x31 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && x13 && x33 && x15 && ~x14 && ~x31 && ~x10 )
						nx_state = s1;
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && x13 && x33 && ~x15 && x14 && x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s343;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && x13 && x33 && ~x15 && x14 && ~x5 )
						begin
							y53 = 1'b1;	
							nx_state = s344;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && x13 && x33 && ~x15 && ~x14 && x16 && x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s340;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && x13 && x33 && ~x15 && ~x14 && x16 && ~x5 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && x13 && x33 && ~x15 && ~x14 && ~x16 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && x13 && x33 && ~x15 && ~x14 && ~x16 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && x13 && x33 && ~x15 && ~x14 && ~x16 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && x13 && x33 && ~x15 && ~x14 && ~x16 && ~x10 )
						nx_state = s1;
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && x13 && ~x33 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y35 = 1'b1;	y40 = 1'b1;	
							nx_state = s351;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && ~x13 && x33 && x14 && x15 && x8 && x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s340;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && ~x13 && x33 && x14 && x15 && x8 && ~x5 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && ~x13 && x33 && x14 && x15 && ~x8 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && ~x13 && x33 && x14 && x15 && ~x8 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && ~x13 && x33 && x14 && x15 && ~x8 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && ~x13 && x33 && x14 && x15 && ~x8 && ~x10 )
						nx_state = s1;
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && ~x13 && x33 && x14 && ~x15 && x30 && x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s340;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && ~x13 && x33 && x14 && ~x15 && x30 && ~x5 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && ~x13 && x33 && x14 && ~x15 && ~x30 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && ~x13 && x33 && x14 && ~x15 && ~x30 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && ~x13 && x33 && x14 && ~x15 && ~x30 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && ~x13 && x33 && x14 && ~x15 && ~x30 && ~x10 )
						nx_state = s1;
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && ~x13 && x33 && ~x14 && x15 && x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s340;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && ~x13 && x33 && ~x14 && x15 && ~x5 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && ~x13 && x33 && ~x14 && ~x15 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s345;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && ~x13 && ~x33 && x4 && x6 )
						begin
							y6 = 1'b1;	y35 = 1'b1;	y40 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s355;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && ~x13 && ~x33 && x4 && ~x6 )
						begin
							y15 = 1'b1;	
							nx_state = s22;
						end
					else if( x69 && x70 && x62 && x64 && x9 && ~x32 && ~x13 && ~x33 && ~x4 )
						begin
							y15 = 1'b1;	
							nx_state = s356;
						end
					else if( x69 && x70 && x62 && x64 && ~x9 )
						begin
							y6 = 1'b1;	y40 = 1'b1;	y41 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s346;
						end
					else if( x69 && x70 && x62 && ~x64 && x66 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x64 && ~x66 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x66 && ~x7 && x9 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x66 && ~x7 && ~x9 && x10 && x6 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x66 && ~x7 && ~x9 && x10 && ~x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x66 && ~x7 && ~x9 && ~x10 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && x62 && ~x64 && ~x66 && ~x7 && ~x9 && ~x10 && ~x11 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && x64 && x63 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x69 && x70 && ~x62 && x64 && x63 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x69 && x70 && ~x62 && x64 && x63 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && x63 && ~x14 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && x66 && x63 && x30 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && x66 && x63 && ~x30 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && x66 && ~x63 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && x3 && x11 && x2 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && x3 && x11 && ~x2 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && x3 && ~x11 && x4 && x12 && x13 && x2 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && x3 && ~x11 && x4 && x12 && x13 && ~x2 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && x3 && ~x11 && x4 && x12 && ~x13 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && x3 && ~x11 && x4 && ~x12 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && x3 && ~x11 && ~x4 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && x4 && x11 && x2 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s670;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && x4 && x11 && ~x2 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && x4 && ~x11 && x12 && x13 && x14 && x2 )
						begin
							y3 = 1'b1;	y22 = 1'b1;	y23 = 1'b1;	
							nx_state = s671;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && x4 && ~x11 && x12 && x13 && x14 && ~x2 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && x4 && ~x11 && x12 && x13 && ~x14 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s230;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && x4 && ~x11 && x12 && x13 && ~x14 && ~x2 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && x4 && ~x11 && x12 && ~x13 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && x4 && ~x11 && x12 && ~x13 && ~x2 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && x4 && ~x11 && ~x12 && x2 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && x4 && ~x11 && ~x12 && ~x2 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && x5 && x6 && x2 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && x5 && x6 && ~x2 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && x7 && x8 && x2 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && x7 && x8 && ~x2 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && x7 && ~x8 && x2 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	
							nx_state = s276;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && x7 && ~x8 && ~x2 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && x8 && x2 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	
							nx_state = s276;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && x8 && ~x2 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && ~x8 && x2 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && ~x8 && ~x2 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && x7 && x9 && x2 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && x7 && x9 && ~x2 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && x7 && ~x9 && x2 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	
							nx_state = s276;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && x7 && ~x9 && ~x2 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && x9 && x2 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	
							nx_state = s276;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && x9 && ~x2 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && ~x9 && x2 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && ~x9 && ~x2 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && x10 && x2 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && x10 && ~x2 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && ~x10 && x2 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	
							nx_state = s276;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && ~x10 && ~x2 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && x10 && x2 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	
							nx_state = s276;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && x10 && ~x2 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && ~x10 && x2 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && ~x10 && ~x2 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && ~x15 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && ~x15 && ~x7 && x9 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && ~x15 && ~x7 && ~x9 && x10 && x6 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && ~x15 && ~x7 && ~x9 && x10 && ~x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && ~x15 && ~x7 && ~x9 && ~x10 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && x63 && ~x15 && ~x7 && ~x9 && ~x10 && ~x11 )
						nx_state = s77;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && x6 && x5 && x7 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && x6 && x5 && x7 && ~x9 )
						begin
							y75 = 1'b1;	
							nx_state = s672;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && x6 && x5 && ~x7 && x8 && x9 && x12 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && x6 && x5 && ~x7 && x8 && x9 && ~x12 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && x6 && x5 && ~x7 && x8 && x9 && ~x12 && x20 && ~x13 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && x6 && x5 && ~x7 && x8 && x9 && ~x12 && ~x20 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && x6 && x5 && ~x7 && x8 && ~x9 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && x6 && x5 && ~x7 && x8 && ~x9 && ~x13 && x20 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && x6 && x5 && ~x7 && x8 && ~x9 && ~x13 && x20 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && x6 && x5 && ~x7 && x8 && ~x9 && ~x13 && ~x20 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && x6 && x5 && ~x7 && ~x8 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y24 = 1'b1;	
							y25 = 1'b1;	y26 = 1'b1;	
							nx_state = s672;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && x6 && x5 && ~x7 && ~x8 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	y29 = 1'b1;	
							nx_state = s673;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && x6 && ~x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s674;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && ~x6 && x11 && x8 && x9 && x5 && x7 )
						begin
							y47 = 1'b1;	
							nx_state = s675;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && ~x6 && x11 && x8 && x9 && x5 && ~x7 )
						begin
							y51 = 1'b1;	
							nx_state = s655;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && ~x6 && x11 && x8 && x9 && ~x5 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	y16 = 1'b1;	
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s672;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && ~x6 && x11 && x8 && ~x9 && x5 && x7 )
						begin
							y48 = 1'b1;	
							nx_state = s676;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && ~x6 && x11 && x8 && ~x9 && x5 && ~x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s677;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && ~x6 && x11 && x8 && ~x9 && ~x5 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s672;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && ~x6 && x11 && ~x8 && x5 && x7 && x9 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && ~x6 && x11 && ~x8 && x5 && x7 && ~x9 )
						begin
							y50 = 1'b1;	
							nx_state = s658;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && ~x6 && x11 && ~x8 && x5 && ~x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y55 = 1'b1;	
							nx_state = s672;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && ~x6 && x11 && ~x8 && ~x5 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	y16 = 1'b1;	
							y18 = 1'b1;	y20 = 1'b1;	
							nx_state = s672;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && x3 && ~x6 && ~x11 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s674;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && x67 && ~x3 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s678;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && ~x67 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && ~x67 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && ~x67 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && x65 && ~x66 && ~x63 && ~x67 && ~x15 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && x66 && x16 && x63 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && x66 && x16 && x63 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && x66 && x16 && x63 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && x66 && x16 && ~x63 )
						begin
							y11 = 1'b1;	
							nx_state = s271;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && x66 && ~x16 && x63 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && x66 && ~x16 && ~x63 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && x66 && ~x16 && ~x63 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && x66 && ~x16 && ~x63 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && x66 && ~x16 && ~x63 && ~x8 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && ~x66 && x63 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && ~x66 && x63 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && ~x66 && x63 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && ~x66 && x63 && ~x1 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && ~x66 && ~x63 && x67 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && ~x66 && ~x63 && x67 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && ~x66 && ~x63 && x67 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && ~x66 && ~x63 && x67 && ~x17 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && ~x66 && ~x63 && ~x67 && x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && ~x66 && ~x63 && ~x67 && x26 && ~x25 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && ~x66 && ~x63 && ~x67 && x26 && ~x25 && ~x24 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && ~x65 && ~x66 && ~x63 && ~x67 && ~x26 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && x67 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x66 && x65 && x67 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x66 && x65 && x67 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && x67 && x22 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && x67 && ~x22 && x18 && x13 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && ~x70 && x66 && x65 && x67 && ~x22 && x18 && x13 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x66 && x65 && x67 && ~x22 && x18 && ~x13 && x12 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && ~x70 && x66 && x65 && x67 && ~x22 && x18 && ~x13 && x12 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x66 && x65 && x67 && ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && x67 && ~x22 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && x20 && x12 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && x20 && x12 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && x20 && x12 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && x20 && x12 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && x20 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && ~x67 && x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && ~x67 && ~x21 && x12 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && ~x21 && x12 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x67 && ~x21 && x12 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && ~x67 && ~x21 && x12 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && ~x67 && ~x21 && ~x12 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && x62 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && x62 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && x62 && ~x15 && x16 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && x62 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y28 = 1'b1;	
							nx_state = s299;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && x63 && x6 && x15 && x8 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && x63 && x6 && x15 && ~x8 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && x63 && x6 && ~x15 && x16 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && x63 && x6 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s468;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && x63 && ~x6 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && ~x63 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && x21 && x16 && x15 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s181;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && x21 && x16 && x15 && ~x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s441;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && x21 && x16 && ~x15 && x10 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && x21 && x16 && ~x15 && ~x10 )
						begin
							y14 = 1'b1;	y16 = 1'b1;	
							nx_state = s492;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && x21 && ~x16 && x17 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s679;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && x21 && ~x16 && x17 && ~x10 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	
							nx_state = s220;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && x21 && ~x16 && ~x17 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s680;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && x21 && ~x16 && ~x17 && ~x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s443;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x10 && x22 && x4 && x17 && x15 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x10 && x22 && x4 && x17 && ~x15 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x10 && x22 && x4 && ~x17 && x18 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x10 && x22 && x4 && ~x17 && ~x18 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x10 && x22 && ~x4 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x10 && ~x22 && x7 && x16 && x15 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x10 && ~x22 && x7 && x16 && ~x15 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s579;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x10 && ~x22 && x7 && ~x16 && x17 && x15 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x10 && ~x22 && x7 && ~x16 && x17 && ~x15 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s579;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x10 && ~x22 && x7 && ~x16 && ~x17 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x10 && ~x22 && ~x7 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s579;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && x17 && x4 && x15 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && x17 && x4 && ~x15 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	
							nx_state = s268;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && x17 && ~x4 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && x15 && x12 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && x15 && ~x12 && x14 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && x15 && ~x12 && ~x14 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && x15 && ~x12 && ~x14 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && x15 && ~x12 && ~x14 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && x15 && ~x12 && ~x14 && ~x7 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && ~x15 && x14 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && ~x15 && x14 && ~x13 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && ~x15 && x14 && ~x13 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && ~x15 && x14 && ~x13 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && ~x15 && x14 && ~x13 && ~x7 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && ~x15 && ~x14 && x11 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && ~x15 && ~x14 && ~x11 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && ~x15 && ~x14 && ~x11 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && ~x15 && ~x14 && ~x11 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && ~x15 && ~x14 && ~x11 && ~x7 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && ~x18 && x4 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s579;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && ~x18 && ~x4 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && x16 && x7 && x15 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s681;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && x16 && x7 && ~x15 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && x16 && ~x7 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s579;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && x14 && x13 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s579;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && x14 && ~x13 && x15 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s579;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && x14 && ~x13 && ~x15 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && x14 && ~x13 && ~x15 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && x14 && ~x13 && ~x15 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && x14 && ~x13 && ~x15 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && ~x14 && x15 && x12 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s579;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && ~x14 && x15 && ~x12 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && ~x14 && x15 && ~x12 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && ~x14 && x15 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && ~x14 && x15 && ~x12 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && ~x14 && ~x15 && x11 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s579;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && ~x14 && ~x15 && ~x11 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && ~x14 && ~x15 && ~x11 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && ~x14 && ~x15 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && ~x14 && ~x15 && ~x11 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && ~x17 && x7 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && ~x17 && ~x7 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s579;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x21 && x67 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && x21 && ~x67 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x21 && ~x67 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x21 && ~x67 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && x21 && ~x67 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x22 && x67 && x23 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x22 && x67 && x23 && ~x18 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x22 && x67 && x23 && ~x18 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x22 && x67 && x23 && ~x18 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x22 && x67 && x23 && ~x18 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x22 && x67 && ~x23 )
						begin
							y6 = 1'b1;	y19 = 1'b1;	
							nx_state = s682;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x22 && ~x67 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x22 && ~x67 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x22 && ~x67 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x22 && ~x67 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && x22 && ~x67 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && x67 && x23 )
						begin
							y6 = 1'b1;	y19 = 1'b1;	
							nx_state = s682;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && x67 && ~x23 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && x67 && ~x23 && ~x19 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && x67 && ~x23 && ~x19 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && x67 && ~x23 && ~x19 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && x67 && ~x23 && ~x19 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && x7 && x23 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && x7 && x23 && ~x9 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && x7 && ~x23 && x9 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && x7 && ~x23 && ~x9 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s296;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && x8 && x23 && x9 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s296;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && x8 && x23 && ~x9 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s297;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && x8 && ~x23 && x9 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s297;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && x8 && ~x23 && ~x9 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s333;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && x23 && x13 && x9 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && x23 && x13 && ~x9 && x14 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && x23 && x13 && ~x9 && ~x14 && x20 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && x23 && x13 && ~x9 && ~x14 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && x23 && ~x13 && x14 && x9 && x20 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && x23 && ~x13 && x14 && x9 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && x23 && ~x13 && x14 && ~x9 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && x23 && ~x13 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && ~x23 && x13 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s683;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && ~x23 && x13 && ~x9 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s683;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && ~x23 && x13 && ~x9 && ~x14 && x18 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && ~x23 && x13 && ~x9 && ~x14 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && ~x23 && ~x13 && x14 && x9 && x18 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && ~x23 && ~x13 && x14 && x9 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && ~x23 && ~x13 && x14 && ~x9 )
						begin
							y22 = 1'b1;	
							nx_state = s683;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && ~x23 && ~x13 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && ~x16 && x7 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && ~x16 && ~x7 && x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && ~x16 && ~x7 && ~x8 && x5 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && ~x16 && ~x7 && ~x8 && ~x5 && x2 && x23 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && ~x16 && ~x7 && ~x8 && ~x5 && x2 && ~x23 && x9 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && ~x16 && ~x7 && ~x8 && ~x5 && x2 && ~x23 && ~x9 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && ~x16 && ~x7 && ~x8 && ~x5 && ~x2 && x9 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && ~x16 && ~x7 && ~x8 && ~x5 && ~x2 && ~x9 && x23 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && ~x16 && ~x7 && ~x8 && ~x5 && ~x2 && ~x9 && ~x23 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && x5 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && x9 && x10 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && x9 && ~x10 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && x9 && ~x10 && ~x8 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && x9 && ~x10 && ~x8 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && x9 && ~x10 && ~x8 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && x9 && ~x10 && ~x8 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && ~x9 && x8 && x12 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && ~x9 && x8 && ~x12 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && ~x9 && x8 && ~x12 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && ~x9 && x8 && ~x12 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && ~x9 && x8 && ~x12 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && ~x9 && ~x8 && x11 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && ~x9 && ~x8 && ~x11 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && ~x9 && ~x8 && ~x11 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && ~x9 && ~x8 && ~x11 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && ~x9 && ~x8 && ~x11 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && ~x16 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && ~x16 && ~x2 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s333;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && x9 && ~x10 && x8 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && x9 && ~x10 && ~x8 && x18 && x14 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && x9 && ~x10 && ~x8 && x18 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && x9 && ~x10 && ~x8 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && x9 && ~x10 && ~x8 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && ~x9 && x8 && x12 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && ~x9 && x8 && ~x12 && x18 && x14 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && ~x9 && x8 && ~x12 && x18 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && ~x9 && x8 && ~x12 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && ~x9 && x8 && ~x12 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && ~x9 && ~x8 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && ~x9 && ~x8 && ~x11 && x18 && x14 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && ~x9 && ~x8 && ~x11 && x18 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && ~x9 && ~x8 && ~x11 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && ~x9 && ~x8 && ~x11 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && ~x16 && x2 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && ~x16 && ~x2 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s495;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x20 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && x21 && x9 && x3 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && x21 && x9 && ~x3 && x4 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && x21 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && x21 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && x12 && x19 && x15 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && x12 && x19 && ~x15 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s315;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && x12 && ~x19 && x20 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && x12 && ~x19 && ~x20 )
						begin
							y6 = 1'b1;	y21 = 1'b1;	
							nx_state = s684;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else if( ~x69 )
						nx_state = s1;
					else nx_state = s77;
				s78 : if( x70 && x69 && x62 && x5 && x4 && x2 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x70 && x69 && x62 && x5 && x4 && ~x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s479;
						end
					else if( x70 && x69 && x62 && x5 && ~x4 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s633;
						end
					else if( x70 && x69 && x62 && ~x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s633;
						end
					else if( x70 && x69 && ~x62 && x63 && x15 && x16 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s637;
						end
					else if( x70 && x69 && ~x62 && x63 && x15 && x16 && ~x1 && x5 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y22 = 1'b1;	
							nx_state = s61;
						end
					else if( x70 && x69 && ~x62 && x63 && x15 && x16 && ~x1 && ~x5 && x6 && x2 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( x70 && x69 && ~x62 && x63 && x15 && x16 && ~x1 && ~x5 && x6 && x2 && ~x3 )
						nx_state = s1;
					else if( x70 && x69 && ~x62 && x63 && x15 && x16 && ~x1 && ~x5 && x6 && ~x2 )
						nx_state = s1;
					else if( x70 && x69 && ~x62 && x63 && x15 && x16 && ~x1 && ~x5 && ~x6 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s638;
						end
					else if( x70 && x69 && ~x62 && x63 && x15 && ~x16 && x7 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s638;
						end
					else if( x70 && x69 && ~x62 && x63 && x15 && ~x16 && ~x7 && x9 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s638;
						end
					else if( x70 && x69 && ~x62 && x63 && x15 && ~x16 && ~x7 && ~x9 && x10 && x6 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x70 && x69 && ~x62 && x63 && x15 && ~x16 && ~x7 && ~x9 && x10 && ~x6 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s636;
						end
					else if( x70 && x69 && ~x62 && x63 && x15 && ~x16 && ~x7 && ~x9 && ~x10 && x11 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s637;
						end
					else if( x70 && x69 && ~x62 && x63 && x15 && ~x16 && ~x7 && ~x9 && ~x10 && ~x11 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && x16 && x5 && x4 && x2 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && x16 && x5 && x4 && ~x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && x16 && x5 && ~x4 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s637;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && x16 && ~x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s637;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && x3 && x11 && x2 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && x3 && x11 && ~x2 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && x3 && ~x11 && x4 && x12 && x13 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && x3 && ~x11 && x4 && x12 && x13 && ~x2 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && x3 && ~x11 && x4 && x12 && ~x13 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && x3 && ~x11 && x4 && ~x12 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && x3 && ~x11 && ~x4 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && x4 && x11 && x2 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s670;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && x4 && x11 && ~x2 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && x4 && ~x11 && x12 && x13 && x14 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s686;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && x4 && ~x11 && x12 && x13 && x14 && ~x2 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && x4 && ~x11 && x12 && x13 && ~x14 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && x4 && ~x11 && x12 && x13 && ~x14 && ~x2 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && x4 && ~x11 && x12 && ~x13 && x2 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y22 = 1'b1;	
							nx_state = s61;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && x4 && ~x11 && x12 && ~x13 && ~x2 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && x4 && ~x11 && ~x12 && x2 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && x4 && ~x11 && ~x12 && ~x2 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && x5 && x6 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s637;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && x5 && x6 && ~x2 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && x7 && x8 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s637;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && x7 && x8 && ~x2 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && x7 && ~x8 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && x7 && ~x8 && ~x2 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && x8 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && x8 && ~x2 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && ~x8 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s637;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && ~x8 && ~x2 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && x7 && x9 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s637;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && x7 && x9 && ~x2 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && x7 && ~x9 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && x7 && ~x9 && ~x2 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && x9 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && x9 && ~x2 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && ~x9 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s637;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && ~x9 && ~x2 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && x10 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s637;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && x10 && ~x2 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && ~x10 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && ~x10 && ~x2 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && x10 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && x10 && ~x2 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && ~x10 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s637;
						end
					else if( x70 && x69 && ~x62 && x63 && ~x15 && ~x16 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && ~x10 && ~x2 )
						nx_state = s78;
					else if( x70 && x69 && ~x62 && ~x63 && x18 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x70 && x69 && ~x62 && ~x63 && ~x18 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( x70 && ~x69 && x63 && x46 && x34 && x42 && x2 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y12 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s687;
						end
					else if( x70 && ~x69 && x63 && x46 && x34 && x42 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && x63 && x46 && x34 && ~x42 && x3 && x35 && x43 && x44 && x2 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s688;
						end
					else if( x70 && ~x69 && x63 && x46 && x34 && ~x42 && x3 && x35 && x43 && x44 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && x63 && x46 && x34 && ~x42 && x3 && x35 && x43 && ~x44 )
						nx_state = s78;
					else if( x70 && ~x69 && x63 && x46 && x34 && ~x42 && x3 && x35 && ~x43 )
						nx_state = s78;
					else if( x70 && ~x69 && x63 && x46 && x34 && ~x42 && x3 && ~x35 )
						nx_state = s78;
					else if( x70 && ~x69 && x63 && x46 && x34 && ~x42 && ~x3 && x35 && x43 && x44 && x2 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s689;
						end
					else if( x70 && ~x69 && x63 && x46 && x34 && ~x42 && ~x3 && x35 && x43 && x44 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && x63 && x46 && x34 && ~x42 && ~x3 && x35 && x43 && ~x44 )
						nx_state = s78;
					else if( x70 && ~x69 && x63 && x46 && x34 && ~x42 && ~x3 && x35 && ~x43 )
						nx_state = s78;
					else if( x70 && ~x69 && x63 && x46 && x34 && ~x42 && ~x3 && ~x35 )
						nx_state = s78;
					else if( x70 && ~x69 && x63 && x46 && ~x34 && x33 && x4 && x11 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y29 = 1'b1;	
							nx_state = s690;
						end
					else if( x70 && ~x69 && x63 && x46 && ~x34 && x33 && x4 && ~x11 && x12 && x13 && x14 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s689;
						end
					else if( x70 && ~x69 && x63 && x46 && ~x34 && x33 && x4 && ~x11 && x12 && x13 && ~x14 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s691;
						end
					else if( x70 && ~x69 && x63 && x46 && ~x34 && x33 && x4 && ~x11 && x12 && ~x13 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s692;
						end
					else if( x70 && ~x69 && x63 && x46 && ~x34 && x33 && x4 && ~x11 && ~x12 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s693;
						end
					else if( x70 && ~x69 && x63 && x46 && ~x34 && x33 && ~x4 && x5 && x37 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( x70 && ~x69 && x63 && x46 && ~x34 && x33 && ~x4 && x5 && ~x37 && x7 && x39 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( x70 && ~x69 && x63 && x46 && ~x34 && x33 && ~x4 && x5 && ~x37 && x7 && ~x39 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( x70 && ~x69 && x63 && x46 && ~x34 && x33 && ~x4 && x5 && ~x37 && ~x7 && x8 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( x70 && ~x69 && x63 && x46 && ~x34 && x33 && ~x4 && x5 && ~x37 && ~x7 && ~x8 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( x70 && ~x69 && x63 && x46 && ~x34 && x33 && ~x4 && ~x5 && x6 && x38 && x40 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( x70 && ~x69 && x63 && x46 && ~x34 && x33 && ~x4 && ~x5 && x6 && x38 && ~x40 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( x70 && ~x69 && x63 && x46 && ~x34 && x33 && ~x4 && ~x5 && x6 && ~x38 && x9 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( x70 && ~x69 && x63 && x46 && ~x34 && x33 && ~x4 && ~x5 && x6 && ~x38 && ~x9 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( x70 && ~x69 && x63 && x46 && ~x34 && x33 && ~x4 && ~x5 && ~x6 && x7 && x10 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( x70 && ~x69 && x63 && x46 && ~x34 && x33 && ~x4 && ~x5 && ~x6 && x7 && ~x10 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( x70 && ~x69 && x63 && x46 && ~x34 && x33 && ~x4 && ~x5 && ~x6 && ~x7 && x41 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( x70 && ~x69 && x63 && x46 && ~x34 && x33 && ~x4 && ~x5 && ~x6 && ~x7 && ~x41 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( x70 && ~x69 && x63 && x46 && ~x34 && ~x33 )
						nx_state = s78;
					else if( x70 && ~x69 && x63 && ~x46 && x38 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y27 = 1'b1;	
							nx_state = s696;
						end
					else if( x70 && ~x69 && x63 && ~x46 && ~x38 && x40 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y27 = 1'b1;	
							nx_state = s696;
						end
					else if( x70 && ~x69 && x63 && ~x46 && ~x38 && ~x40 && x10 && x37 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x70 && ~x69 && x63 && ~x46 && ~x38 && ~x40 && x10 && ~x37 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s697;
						end
					else if( x70 && ~x69 && x63 && ~x46 && ~x38 && ~x40 && ~x10 && x42 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( x70 && ~x69 && x63 && ~x46 && ~x38 && ~x40 && ~x10 && ~x42 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && x3 && x11 && x64 && x2 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s698;
						end
					else if( x70 && ~x69 && ~x63 && x15 && x3 && x11 && x64 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && x3 && x11 && ~x64 && x2 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s447;
						end
					else if( x70 && ~x69 && ~x63 && x15 && x3 && x11 && ~x64 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && x3 && ~x11 && x4 && x12 && x13 && x2 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s688;
						end
					else if( x70 && ~x69 && ~x63 && x15 && x3 && ~x11 && x4 && x12 && x13 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && x3 && ~x11 && x4 && x12 && ~x13 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && x3 && ~x11 && x4 && ~x12 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && x3 && ~x11 && ~x4 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && x4 && x11 && x64 && x2 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s670;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && x4 && x11 && x64 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && x4 && x11 && ~x64 && x33 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s670;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && x4 && x11 && ~x64 && ~x33 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && x4 && ~x11 && x12 && x13 && x14 && x64 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s699;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && x4 && ~x11 && x12 && x13 && x14 && x64 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && x4 && ~x11 && x12 && x13 && x14 && ~x64 && x33 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s699;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && x4 && ~x11 && x12 && x13 && x14 && ~x64 && ~x33 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && x4 && ~x11 && x12 && x13 && ~x14 && x64 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && x4 && ~x11 && x12 && x13 && ~x14 && x64 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && x4 && ~x11 && x12 && x13 && ~x14 && ~x64 && x33 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s700;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && x4 && ~x11 && x12 && x13 && ~x14 && ~x64 && ~x33 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && x4 && ~x11 && x12 && ~x13 && x64 && x2 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s692;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && x4 && ~x11 && x12 && ~x13 && x64 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && x4 && ~x11 && x12 && ~x13 && ~x64 && x33 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s701;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && x4 && ~x11 && x12 && ~x13 && ~x64 && ~x33 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && x4 && ~x11 && ~x12 && x64 && x2 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s693;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && x4 && ~x11 && ~x12 && x64 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && x4 && ~x11 && ~x12 && ~x64 && x33 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s702;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && x4 && ~x11 && ~x12 && ~x64 && ~x33 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && x5 && x6 && x64 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && x5 && x6 && x64 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && x5 && x6 && ~x64 && x33 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s703;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && x5 && x6 && ~x64 && ~x33 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && x7 && x8 && x64 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && x7 && x8 && x64 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && x7 && x8 && ~x64 && x33 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s703;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && x7 && x8 && ~x64 && ~x33 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && x7 && ~x8 && x64 && x2 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && x7 && ~x8 && x64 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && x7 && ~x8 && ~x64 && x33 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && x7 && ~x8 && ~x64 && ~x33 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && x8 && x64 && x2 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && x8 && x64 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && x8 && ~x64 && x33 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && x8 && ~x64 && ~x33 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && ~x8 && x64 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && ~x8 && x64 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && ~x8 && ~x64 && x33 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s703;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && ~x8 && ~x64 && ~x33 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && x7 && x9 && x64 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && x7 && x9 && x64 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && x7 && x9 && ~x64 && x33 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s703;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && x7 && x9 && ~x64 && ~x33 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && x7 && ~x9 && x64 && x2 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && x7 && ~x9 && x64 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && x7 && ~x9 && ~x64 && x33 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && x7 && ~x9 && ~x64 && ~x33 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && x9 && x64 && x2 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && x9 && x64 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && x9 && ~x64 && x33 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && x9 && ~x64 && ~x33 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && ~x9 && x64 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && ~x9 && x64 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && ~x9 && ~x64 && x33 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s703;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && ~x9 && ~x64 && ~x33 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && x10 && x64 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && x10 && x64 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && x10 && ~x64 && x33 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s703;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && x10 && ~x64 && ~x33 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && ~x10 && x64 && x2 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && ~x10 && x64 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && ~x10 && ~x64 && x33 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && ~x10 && ~x64 && ~x33 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && x10 && x64 && x2 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && x10 && x64 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && x10 && ~x64 && x33 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && x10 && ~x64 && ~x33 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && ~x10 && x64 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && ~x10 && x64 && ~x2 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && ~x10 && ~x64 && x33 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s703;
						end
					else if( x70 && ~x69 && ~x63 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && ~x10 && ~x64 && ~x33 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && ~x15 && x7 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s704;
						end
					else if( x70 && ~x69 && ~x63 && ~x15 && ~x7 && x9 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s704;
						end
					else if( x70 && ~x69 && ~x63 && ~x15 && ~x7 && ~x9 && x10 && x6 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x70 && ~x69 && ~x63 && ~x15 && ~x7 && ~x9 && x10 && ~x6 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s705;
						end
					else if( x70 && ~x69 && ~x63 && ~x15 && ~x7 && ~x9 && ~x10 && x64 && x11 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( x70 && ~x69 && ~x63 && ~x15 && ~x7 && ~x9 && ~x10 && x64 && ~x11 )
						nx_state = s78;
					else if( x70 && ~x69 && ~x63 && ~x15 && ~x7 && ~x9 && ~x10 && ~x64 && x11 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s703;
						end
					else if( x70 && ~x69 && ~x63 && ~x15 && ~x7 && ~x9 && ~x10 && ~x64 && ~x11 )
						nx_state = s78;
					else if( ~x70 && x69 && x61 && x60 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s139;
						end
					else if( ~x70 && x69 && x61 && ~x60 && x62 )
						nx_state = s1;
					else if( ~x70 && x69 && x61 && ~x60 && ~x62 )
						nx_state = s118;
					else if( ~x70 && x69 && ~x61 && x60 )
						nx_state = s118;
					else if( ~x70 && x69 && ~x61 && ~x60 && x62 && x4 && x15 && x12 && x7 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s592;
						end
					else if( ~x70 && x69 && ~x61 && ~x60 && x62 && x4 && x15 && x12 && ~x7 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s706;
						end
					else if( ~x70 && x69 && ~x61 && ~x60 && x62 && x4 && x15 && ~x12 && x7 )
						nx_state = s331;
					else if( ~x70 && x69 && ~x61 && ~x60 && x62 && x4 && x15 && ~x12 && ~x7 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x69 && ~x61 && ~x60 && x62 && x4 && ~x15 && x16 && x7 && x12 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s706;
						end
					else if( ~x70 && x69 && ~x61 && ~x60 && x62 && x4 && ~x15 && x16 && x7 && ~x12 )
						nx_state = s331;
					else if( ~x70 && x69 && ~x61 && ~x60 && x62 && x4 && ~x15 && x16 && ~x7 )
						nx_state = s331;
					else if( ~x70 && x69 && ~x61 && ~x60 && x62 && x4 && ~x15 && ~x16 && x7 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s707;
						end
					else if( ~x70 && x69 && ~x61 && ~x60 && x62 && x4 && ~x15 && ~x16 && ~x7 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && x69 && ~x61 && ~x60 && x62 && ~x4 )
						nx_state = s331;
					else if( ~x70 && x69 && ~x61 && ~x60 && ~x62 && x15 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( ~x70 && x69 && ~x61 && ~x60 && ~x62 && x15 && ~x7 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x69 && ~x61 && ~x60 && ~x62 && x15 && ~x7 && ~x11 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x70 && x69 && ~x61 && ~x60 && ~x62 && ~x15 && x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( ~x70 && x69 && ~x61 && ~x60 && ~x62 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && ~x69 && x5 && x6 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x69 && x5 && ~x6 && x7 )
						nx_state = s1;
					else if( ~x70 && ~x69 && x5 && ~x6 && ~x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							nx_state = s38;
						end
					else if( ~x70 && ~x69 && ~x5 && x4 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && ~x69 && ~x5 && ~x4 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else nx_state = s78;
				s79 : if( 1'b1 )
						begin
							y2 = 1'b1;	
							nx_state = s708;
						end
					else nx_state = s79;
				s80 : if( 1'b1 )
						begin
							y19 = 1'b1;	
							nx_state = s13;
						end
					else nx_state = s80;
				s81 : if( x62 && x32 && x33 )
						begin
							y9 = 1'b1;	
							nx_state = s709;
						end
					else if( x62 && x32 && ~x33 && x8 )
						begin
							y9 = 1'b1;	
							nx_state = s709;
						end
					else if( x62 && x32 && ~x33 && ~x8 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s470;
						end
					else if( x62 && ~x32 && x8 )
						begin
							y9 = 1'b1;	
							nx_state = s709;
						end
					else if( x62 && ~x32 && ~x8 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s470;
						end
					else if( ~x62 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else nx_state = s81;
				s82 : if( x69 && x64 && x65 )
						begin
							y8 = 1'b1;	
							nx_state = s568;
						end
					else if( x69 && x64 && ~x65 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x69 && ~x64 && x65 && x31 && x30 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( x69 && ~x64 && x65 && x31 && ~x30 )
						begin
							y3 = 1'b1;	
							nx_state = s710;
						end
					else if( x69 && ~x64 && x65 && ~x31 && x30 )
						begin
							y3 = 1'b1;	
							nx_state = s462;
						end
					else if( x69 && ~x64 && x65 && ~x31 && ~x30 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( x69 && ~x64 && ~x65 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s57;
						end
					else if( ~x69 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else nx_state = s82;
				s83 : if( 1'b1 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s712;
						end
					else nx_state = s83;
				s84 : if( 1'b1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y26 = 1'b1;	
							nx_state = s713;
						end
					else nx_state = s84;
				s85 : if( 1'b1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else nx_state = s85;
				s86 : if( x22 )
						nx_state = s1;
					else if( ~x22 && x15 && x8 )
						begin
							y11 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x22 && x15 && ~x8 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s591;
						end
					else if( ~x22 && ~x15 && x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s126;
						end
					else if( ~x22 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else nx_state = s86;
				s87 : if( x70 && x63 && x64 && x19 && x20 && x2 && x1 && x4 && x3 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x70 && x63 && x64 && x19 && x20 && x2 && x1 && x4 && x3 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x70 && x63 && x64 && x19 && x20 && x2 && x1 && x4 && x3 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( x70 && x63 && x64 && x19 && x20 && x2 && x1 && x4 && x3 && ~x22 )
						nx_state = s1;
					else if( x70 && x63 && x64 && x19 && x20 && x2 && x1 && x4 && ~x3 && x5 && x18 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && x63 && x64 && x19 && x20 && x2 && x1 && x4 && ~x3 && x5 && ~x18 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x70 && x63 && x64 && x19 && x20 && x2 && x1 && x4 && ~x3 && x5 && ~x18 && x22 && ~x21 )
						nx_state = s1;
					else if( x70 && x63 && x64 && x19 && x20 && x2 && x1 && x4 && ~x3 && x5 && ~x18 && ~x22 )
						nx_state = s1;
					else if( x70 && x63 && x64 && x19 && x20 && x2 && x1 && x4 && ~x3 && ~x5 && x21 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && x63 && x64 && x19 && x20 && x2 && x1 && x4 && ~x3 && ~x5 && ~x21 && x22 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x70 && x63 && x64 && x19 && x20 && x2 && x1 && x4 && ~x3 && ~x5 && ~x21 && x22 && ~x18 )
						nx_state = s1;
					else if( x70 && x63 && x64 && x19 && x20 && x2 && x1 && x4 && ~x3 && ~x5 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x70 && x63 && x64 && x19 && x20 && x2 && x1 && ~x4 && x5 && x3 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x70 && x63 && x64 && x19 && x20 && x2 && x1 && ~x4 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	y36 = 1'b1;	
							nx_state = s654;
						end
					else if( x70 && x63 && x64 && x19 && x20 && x2 && x1 && ~x4 && ~x5 && x3 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x70 && x63 && x64 && x19 && x20 && x2 && x1 && ~x4 && ~x5 && ~x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y34 = 1'b1;	y37 = 1'b1;	
							nx_state = s654;
						end
					else if( x70 && x63 && x64 && x19 && x20 && x2 && ~x1 )
						begin
							y26 = 1'b1;	
							nx_state = s413;
						end
					else if( x70 && x63 && x64 && x19 && x20 && ~x2 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s715;
						end
					else if( x70 && x63 && x64 && x19 && x20 && ~x2 && ~x8 )
						begin
							y26 = 1'b1;	
							nx_state = s413;
						end
					else if( x70 && x63 && x64 && x19 && ~x20 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s716;
						end
					else if( x70 && x63 && x64 && ~x19 )
						begin
							y28 = 1'b1;	
							nx_state = s717;
						end
					else if( x70 && x63 && ~x64 && x66 && x31 && x15 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x70 && x63 && ~x64 && x66 && x31 && ~x15 && x16 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && x63 && ~x64 && x66 && x31 && ~x15 && ~x16 )
						begin
							y35 = 1'b1;	
							nx_state = s718;
						end
					else if( x70 && x63 && ~x64 && x66 && ~x31 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x70 && x63 && ~x64 && ~x66 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x70 && x63 && ~x64 && ~x66 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x70 && x63 && ~x64 && ~x66 && x19 && ~x14 && ~x13 && x11 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( x70 && x63 && ~x64 && ~x66 && x19 && ~x14 && ~x13 && x11 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( x70 && x63 && ~x64 && ~x66 && x19 && ~x14 && ~x13 && ~x11 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( x70 && x63 && ~x64 && ~x66 && ~x19 )
						nx_state = s1;
					else if( x70 && ~x63 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x63 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x63 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x17 )
						nx_state = s1;
					else if( ~x70 && x65 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x21 && x16 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s233;
						end
					else if( ~x70 && ~x65 && x21 && x16 && ~x10 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && ~x65 && x21 && ~x16 )
						begin
							y5 = 1'b1;	y17 = 1'b1;	
							nx_state = s721;
						end
					else if( ~x70 && ~x65 && ~x21 )
						nx_state = s1;
					else nx_state = s87;
				s88 : if( x69 && x70 && x62 && x20 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x69 && x70 && x62 && x20 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x69 && x70 && x62 && x20 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( x69 && x70 && x62 && x20 && ~x21 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x20 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && x70 && ~x62 && x63 && x65 && x64 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x69 && x70 && ~x62 && x63 && x65 && x64 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x69 && x70 && ~x62 && x63 && x65 && x64 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x65 && x64 && ~x22 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x65 && ~x64 && x66 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && x70 && ~x62 && x63 && x65 && ~x64 && ~x66 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x69 && x70 && ~x62 && x63 && x65 && ~x64 && ~x66 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x69 && x70 && ~x62 && x63 && x65 && ~x64 && ~x66 && x19 && ~x14 && ~x13 && x11 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( x69 && x70 && ~x62 && x63 && x65 && ~x64 && ~x66 && x19 && ~x14 && ~x13 && x11 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( x69 && x70 && ~x62 && x63 && x65 && ~x64 && ~x66 && x19 && ~x14 && ~x13 && ~x11 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( x69 && x70 && ~x62 && x63 && x65 && ~x64 && ~x66 && ~x19 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x64 && x17 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y22 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s722;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x64 && ~x17 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x64 && ~x17 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x64 && ~x17 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x64 && ~x17 && ~x10 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x65 && ~x64 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && ~x64 && ~x2 && x5 && x3 && x1 )
						nx_state = s88;
					else if( x69 && x70 && ~x62 && x63 && ~x65 && ~x64 && ~x2 && x5 && x3 && ~x1 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && ~x64 && ~x2 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && ~x64 && ~x2 && ~x5 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	
							nx_state = s7;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x66 && x65 && x23 && x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x66 && x65 && x23 && x11 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x66 && x65 && x23 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x66 && x65 && x23 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x66 && x65 && ~x23 && x24 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x66 && x65 && ~x23 && x24 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x66 && x65 && ~x23 && x24 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x66 && x65 && ~x23 && x24 && ~x20 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x66 && x65 && ~x23 && ~x24 && x11 && x12 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x66 && x65 && ~x23 && ~x24 && x11 && ~x12 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x66 && x65 && ~x23 && ~x24 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x66 && x65 && ~x23 && ~x24 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x66 && ~x65 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x66 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && x66 && x22 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y10 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s92;
						end
					else if( x69 && ~x70 && x65 && x67 && x66 && ~x22 && x23 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y10 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s92;
						end
					else if( x69 && ~x70 && x65 && x67 && x66 && ~x22 && ~x23 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x66 && x21 && x18 )
						begin
							y14 = 1'b1;	y19 = 1'b1;	
							nx_state = s723;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x66 && x21 && ~x18 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s724;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x66 && ~x21 && x22 && x8 && x23 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x66 && ~x21 && x22 && x8 && x23 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x66 && ~x21 && x22 && x8 && x23 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x66 && ~x21 && x22 && x8 && ~x23 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x66 && ~x21 && x22 && x8 && ~x23 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x66 && ~x21 && x22 && x8 && ~x23 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x66 && ~x21 && x22 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x66 && ~x21 && ~x22 && x23 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x66 && ~x21 && ~x22 && x23 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x66 && ~x21 && ~x22 && x23 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x66 && ~x21 && ~x22 && x23 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x66 && ~x21 && ~x22 && ~x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x66 && ~x21 && ~x22 && ~x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x66 && ~x21 && ~x22 && ~x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x66 && ~x21 && ~x22 && ~x23 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && x68 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && x61 && x60 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && x61 && x60 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && x61 && x60 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && x61 && x60 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && x61 && ~x60 && x62 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && x61 && ~x60 && ~x62 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s559;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && ~x61 && x60 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s559;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && ~x61 && ~x60 )
						nx_state = s47;
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && x23 && x22 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && x23 && x22 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && x23 && x22 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && x23 && ~x22 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && x23 && ~x22 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && x23 && ~x22 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && x23 && ~x22 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && ~x23 && x18 && x14 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && ~x23 && x18 && x14 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && ~x23 && x18 && ~x14 && x13 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && ~x23 && x18 && ~x14 && x13 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && ~x23 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x68 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x70 && ~x65 && x68 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x70 && ~x65 && x68 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x68 && x21 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x68 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( x69 && ~x70 && ~x65 && x68 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( x69 && ~x70 && ~x65 && x68 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x68 && ~x21 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x68 && x62 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else if( ~x69 && x9 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && ~x9 && x7 )
						nx_state = s1;
					else if( ~x69 && ~x9 && ~x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else nx_state = s88;
				s89 : if( x22 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	
							nx_state = s486;
						end
					else if( ~x22 )
						nx_state = s1;
					else nx_state = s89;
				s90 : if( x69 && x70 && x63 && x64 )
						begin
							y2 = 1'b1;	y17 = 1'b1;	y19 = 1'b1;	
							nx_state = s725;
						end
					else if( x69 && x70 && x63 && ~x64 )
						begin
							y66 = 1'b1;	
							nx_state = s726;
						end
					else if( x69 && x70 && ~x63 && x23 && x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x69 && x70 && ~x63 && x23 && x11 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x69 && x70 && ~x63 && x23 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x69 && x70 && ~x63 && x23 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x63 && ~x23 && x24 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && x70 && ~x63 && ~x23 && x24 && ~x12 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x63 && ~x23 && x24 && ~x12 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x63 && ~x23 && x24 && ~x12 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x69 && x70 && ~x63 && ~x23 && x24 && ~x12 && ~x20 )
						nx_state = s1;
					else if( x69 && x70 && ~x63 && ~x23 && ~x24 && x11 && x12 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && x70 && ~x63 && ~x23 && ~x24 && x11 && ~x12 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && x70 && ~x63 && ~x23 && ~x24 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x69 && x70 && ~x63 && ~x23 && ~x24 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && x66 && x22 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && x66 && ~x22 && x23 && x19 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x69 && ~x70 && x65 && x67 && x66 && ~x22 && x23 && x19 && x15 && ~x8 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && x65 && x67 && x66 && ~x22 && x23 && x19 && ~x15 && x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s126;
						end
					else if( x69 && ~x70 && x65 && x67 && x66 && ~x22 && x23 && x19 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( x69 && ~x70 && x65 && x67 && x66 && ~x22 && x23 && ~x19 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x65 && x67 && x66 && ~x22 && ~x23 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x66 && x21 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x66 && ~x21 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && x68 && x20 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && x68 && ~x20 && x21 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && x68 && ~x20 && x21 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && x68 && ~x20 && x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && x68 && ~x20 && x21 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && x68 && ~x20 && ~x21 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && x60 && x61 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && x60 && x61 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && x60 && x61 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && x60 && x61 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && x60 && ~x61 )
						nx_state = s118;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && x62 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && ~x62 )
						nx_state = s118;
					else if( x69 && ~x70 && x65 && ~x67 && x66 && ~x68 && ~x60 && ~x61 )
						nx_state = s47;
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && x23 && x22 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && x23 && x22 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && x23 && x22 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && x23 && ~x22 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && x23 && ~x22 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && x23 && ~x22 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && x23 && ~x22 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && ~x23 && x18 && x14 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && ~x23 && x18 && x14 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && ~x23 && x18 && ~x14 && x13 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && ~x23 && x18 && ~x14 && x13 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x66 && ~x21 && ~x23 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x68 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x68 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x68 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x68 && x21 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x68 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x68 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x68 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x68 && ~x21 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x21 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x21 && x22 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s170;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x21 && ~x22 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s315;
						end
					else if( ~x69 && x5 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x69 && ~x5 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x5 && ~x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else nx_state = s90;
				s91 : if( x65 && x70 && x64 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( x65 && x70 && ~x64 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && x70 && ~x64 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && x70 && ~x64 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x65 && x70 && ~x64 && ~x23 )
						nx_state = s1;
					else if( x65 && ~x70 && x23 )
						begin
							y2 = 1'b1;	y16 = 1'b1;	y24 = 1'b1;	
							nx_state = s270;
						end
					else if( x65 && ~x70 && ~x23 && x18 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x65 && ~x70 && ~x23 && x18 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x65 && ~x70 && ~x23 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && ~x70 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x70 && x64 )
						begin
							y5 = 1'b1;	y13 = 1'b1;	y30 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s727;
						end
					else if( ~x65 && x70 && ~x64 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x65 && x70 && ~x64 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x65 && x70 && ~x64 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x64 && ~x8 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x65 && ~x70 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x65 && ~x70 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x9 )
						nx_state = s1;
					else nx_state = s91;
				s92 : if( x22 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s426;
						end
					else if( ~x22 && x23 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x22 && x23 && x15 && ~x8 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x22 && x23 && ~x15 && x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s126;
						end
					else if( ~x22 && x23 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( ~x22 && ~x23 )
						begin
							y2 = 1'b1;	y16 = 1'b1;	y24 = 1'b1;	
							nx_state = s270;
						end
					else nx_state = s92;
				s93 : if( x69 && x65 && x66 && x67 && x22 && x16 && x15 && x8 && x14 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && x15 && x8 && ~x14 && x7 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s358;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && x15 && x8 && ~x14 && ~x7 && x12 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && x15 && x8 && ~x14 && ~x7 && ~x12 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && x15 && x8 && ~x14 && ~x7 && ~x12 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && x15 && x8 && ~x14 && ~x7 && ~x12 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && x65 && x66 && x67 && x22 && x16 && x15 && x8 && ~x14 && ~x7 && ~x12 && ~x17 )
						nx_state = s1;
					else if( x69 && x65 && x66 && x67 && x22 && x16 && x15 && ~x8 && x14 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && x15 && ~x8 && ~x14 && x7 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s728;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && x15 && ~x8 && ~x14 && ~x7 && x13 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && x15 && ~x8 && ~x14 && ~x7 && ~x13 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && x15 && ~x8 && ~x14 && ~x7 && ~x13 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && x15 && ~x8 && ~x14 && ~x7 && ~x13 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && x65 && x66 && x67 && x22 && x16 && x15 && ~x8 && ~x14 && ~x7 && ~x13 && ~x17 )
						nx_state = s1;
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && x8 && x9 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && x8 && x9 && ~x2 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && x8 && x9 && ~x2 && ~x4 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s486;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && x8 && ~x9 && x7 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && x8 && ~x9 && x7 && ~x2 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && x8 && ~x9 && x7 && ~x2 && ~x4 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s486;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && x8 && ~x9 && ~x7 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && x8 && ~x9 && ~x7 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && x8 && ~x9 && ~x7 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && x8 && ~x9 && ~x7 && ~x17 )
						nx_state = s1;
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && x7 && x11 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && x7 && x11 && ~x2 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && x7 && x11 && ~x2 && ~x4 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s486;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && x7 && ~x11 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && x7 && ~x11 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && x7 && ~x11 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && x7 && ~x11 && ~x17 )
						nx_state = s1;
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && ~x7 && x10 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && ~x7 && x10 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && ~x7 && x10 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && ~x7 && x10 && ~x17 )
						nx_state = s1;
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x2 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x69 && x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x2 && ~x4 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s486;
						end
					else if( x69 && x65 && x66 && x67 && x22 && ~x16 && x15 && x7 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && x65 && x66 && x67 && x22 && ~x16 && x15 && ~x7 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( x69 && x65 && x66 && x67 && x22 && ~x16 && x15 && ~x7 && ~x2 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x69 && x65 && x66 && x67 && x22 && ~x16 && x15 && ~x7 && ~x2 && ~x4 && x8 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y28 = 1'b1;	
							nx_state = s729;
						end
					else if( x69 && x65 && x66 && x67 && x22 && ~x16 && x15 && ~x7 && ~x2 && ~x4 && ~x8 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s591;
						end
					else if( x69 && x65 && x66 && x67 && x22 && ~x16 && ~x15 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( x69 && x65 && x66 && x67 && x22 && ~x16 && ~x15 && ~x2 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x69 && x65 && x66 && x67 && x22 && ~x16 && ~x15 && ~x2 && ~x4 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && x65 && x66 && x67 && ~x22 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( x69 && x65 && x66 && ~x67 && x21 && x20 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s553;
						end
					else if( x69 && x65 && x66 && ~x67 && x21 && ~x20 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s731;
						end
					else if( x69 && x65 && x66 && ~x67 && ~x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s731;
						end
					else if( x69 && x65 && ~x66 && x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s111;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x23 && x22 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && x23 && ~x22 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s110;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x23 && x22 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s111;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x23 && ~x22 )
						nx_state = s1;
					else if( x69 && ~x65 && x20 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && ~x65 && ~x20 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x69 && x70 && x19 && x62 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s320;
						end
					else if( ~x69 && x70 && x19 && ~x62 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( ~x69 && x70 && ~x19 && x26 && x62 && x5 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x69 && x70 && ~x19 && x26 && x62 && ~x5 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s733;
						end
					else if( ~x69 && x70 && ~x19 && x26 && ~x62 && x63 && x64 && x5 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s734;
						end
					else if( ~x69 && x70 && ~x19 && x26 && ~x62 && x63 && x64 && ~x5 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s735;
						end
					else if( ~x69 && x70 && ~x19 && x26 && ~x62 && x63 && ~x64 && x5 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x70 && ~x19 && x26 && ~x62 && x63 && ~x64 && ~x5 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x69 && x70 && ~x19 && x26 && ~x62 && ~x63 && x5 && x64 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s736;
						end
					else if( ~x69 && x70 && ~x19 && x26 && ~x62 && ~x63 && x5 && ~x64 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s737;
						end
					else if( ~x69 && x70 && ~x19 && x26 && ~x62 && ~x63 && ~x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( ~x69 && x70 && ~x19 && ~x26 && x62 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s738;
						end
					else if( ~x69 && x70 && ~x19 && ~x26 && ~x62 && x64 && x63 )
						begin
							y11 = 1'b1;	y36 = 1'b1;	
							nx_state = s739;
						end
					else if( ~x69 && x70 && ~x19 && ~x26 && ~x62 && x64 && ~x63 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s738;
						end
					else if( ~x69 && x70 && ~x19 && ~x26 && ~x62 && ~x64 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s738;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x4 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s320;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x4 && x1 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x4 && x1 && ~x3 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s733;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x4 && ~x1 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x19 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x19 && x26 && x5 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x19 && x26 && ~x5 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x19 && ~x26 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s738;
						end
					else if( ~x69 && ~x70 && ~x44 && x4 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s320;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x4 && x1 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x4 && x1 && ~x3 )
						begin
							y5 = 1'b1;	y13 = 1'b1;	
							nx_state = s740;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x4 && ~x1 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s738;
						end
					else nx_state = s93;
				s94 : if( x69 && x70 && x62 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x69 && x70 && x62 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x69 && x70 && x62 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x19 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x65 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && x22 && x19 && x8 && x9 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && x22 && x19 && x8 && x9 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && x22 && x19 && x8 && x9 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && x22 && x19 && x8 && x9 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && x22 && x19 && x8 && x9 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && x22 && x19 && x8 && ~x9 && x10 )
						begin
							y33 = 1'b1;	y54 = 1'b1;	
							nx_state = s1;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && x22 && x19 && x8 && ~x9 && ~x10 )
						begin
							y37 = 1'b1;	y55 = 1'b1;	
							nx_state = s1;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && x22 && x19 && ~x8 && x9 && x5 && x10 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && x22 && x19 && ~x8 && x9 && x5 && ~x10 && x4 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && x22 && x19 && ~x8 && x9 && x5 && ~x10 && ~x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && x22 && x19 && ~x8 && x9 && ~x5 && x4 && x10 && x6 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && x22 && x19 && ~x8 && x9 && ~x5 && x4 && x10 && ~x6 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && x22 && x19 && ~x8 && x9 && ~x5 && x4 && ~x10 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && x22 && x19 && ~x8 && x9 && ~x5 && ~x4 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && x22 && x19 && ~x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y26 = 1'b1;	
							y51 = 1'b1;	y56 = 1'b1;	
							nx_state = s741;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && x22 && x19 && ~x8 && ~x9 && ~x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y23 = 1'b1;	
							y52 = 1'b1;	y53 = 1'b1;	
							nx_state = s741;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && x22 && ~x19 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s742;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && ~x22 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && ~x22 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && ~x22 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && ~x22 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && x23 && ~x22 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x65 && ~x23 && x19 && x20 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s523;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && ~x23 && x19 && ~x20 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s743;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x65 && ~x23 && ~x19 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s742;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x65 && x12 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x65 && x12 && ~x8 && x7 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x65 && x12 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x65 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x18 )
						begin
							y59 = 1'b1;	y60 = 1'b1;	
							nx_state = s284;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x18 && x19 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x18 && ~x19 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && x24 && x23 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && x24 && ~x23 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x24 && x11 && x12 && x23 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x24 && x11 && x12 && ~x23 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x24 && x11 && ~x12 && x13 && x23 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x24 && x11 && ~x12 && x13 && ~x23 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x24 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x67 && ~x24 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && ~x67 && x29 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && ~x67 && x29 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && ~x67 && x29 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && ~x67 && x29 && ~x23 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && ~x67 && ~x29 )
						begin
							y8 = 1'b1;	
							nx_state = s744;
						end
					else if( x69 && ~x70 && x65 && x66 && x60 && x61 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && x66 && x60 && x61 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && x66 && x60 && x61 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x65 && x66 && x60 && x61 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x65 && x66 && x60 && ~x61 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x66 && x60 && ~x61 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x66 && x60 && ~x61 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( x69 && ~x70 && x65 && x66 && x60 && ~x61 && ~x18 )
						nx_state = s118;
					else if( x69 && ~x70 && x65 && x66 && ~x60 && x61 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x60 && x61 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x60 && x61 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x66 && ~x60 && x61 && x62 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x66 && ~x60 && x61 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x60 && x61 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x66 && ~x60 && x61 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( x69 && ~x70 && x65 && x66 && ~x60 && x61 && ~x62 && ~x18 )
						nx_state = s118;
					else if( x69 && ~x70 && x65 && x66 && ~x60 && ~x61 )
						nx_state = s47;
					else if( x69 && ~x70 && x65 && ~x66 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && x65 && ~x66 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && ~x66 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && ~x66 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x23 && x22 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x23 && x22 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x23 && x22 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x23 && ~x22 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x23 && ~x22 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x23 && ~x22 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && x23 && ~x22 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && ~x23 && x18 && x14 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && ~x23 && x18 && x14 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && ~x23 && x18 && ~x14 && x13 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && ~x23 && x18 && ~x14 && x13 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x66 && ~x21 && ~x23 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x68 && x5 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x65 && x68 && x5 && ~x18 && x21 && x6 )
						nx_state = s94;
					else if( x69 && ~x70 && ~x65 && x68 && x5 && ~x18 && x21 && ~x6 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && ~x65 && x68 && x5 && ~x18 && ~x21 && x4 )
						nx_state = s94;
					else if( x69 && ~x70 && ~x65 && x68 && x5 && ~x18 && ~x21 && ~x4 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && ~x65 && x68 && ~x5 && x21 && x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( x69 && ~x70 && ~x65 && x68 && ~x5 && x21 && ~x4 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s97;
						end
					else if( x69 && ~x70 && ~x65 && x68 && ~x5 && ~x21 && x6 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && ~x70 && ~x65 && x68 && ~x5 && ~x21 && ~x6 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s97;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x68 && x62 && ~x61 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x68 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else if( ~x69 && x70 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y26 = 1'b1;	
							nx_state = s745;
						end
					else if( ~x69 && ~x70 && x45 && x12 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x69 && ~x70 && x45 && x12 && ~x5 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x45 && x12 && ~x5 && ~x1 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x69 && ~x70 && x45 && ~x12 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( ~x69 && ~x70 && ~x45 && x11 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x11 && x46 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x11 && ~x46 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x11 && ~x46 && ~x5 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x11 && ~x46 && ~x5 && ~x1 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else nx_state = s94;
				s95 : if( x69 && x70 && x64 && x63 )
						begin
							y13 = 1'b1;	y16 = 1'b1;	
							nx_state = s335;
						end
					else if( x69 && x70 && x64 && ~x63 && x65 && x66 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x69 && x70 && x64 && ~x63 && x65 && x66 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x69 && x70 && x64 && ~x63 && x65 && x66 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x63 && x65 && x66 && ~x14 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x63 && x65 && ~x66 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x63 && ~x65 && x66 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && x8 && x6 && x11 && x10 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && x8 && x6 && x11 && x10 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && x8 && x6 && x11 && x10 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && x8 && x6 && x11 && x10 && ~x18 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && x8 && x6 && x11 && ~x10 && x12 && x13 )
						begin
							y7 = 1'b1;	
							nx_state = s747;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && x8 && x6 && x11 && ~x10 && x12 && ~x13 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && x8 && x6 && x11 && ~x10 && x12 && ~x13 && x18 && ~x14 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && x8 && x6 && x11 && ~x10 && x12 && ~x13 && ~x18 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && x8 && x6 && x11 && ~x10 && ~x12 && x14 )
						begin
							y7 = 1'b1;	
							nx_state = s748;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && x8 && x6 && x11 && ~x10 && ~x12 && ~x14 && x18 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && x8 && x6 && x11 && ~x10 && ~x12 && ~x14 && x18 && ~x13 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && x8 && x6 && x11 && ~x10 && ~x12 && ~x14 && ~x18 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && x8 && x6 && ~x11 && x12 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && x8 && x6 && ~x11 && x12 && ~x10 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y27 = 1'b1;	y45 = 1'b1;	
							nx_state = s749;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && x8 && x6 && ~x11 && ~x12 && x10 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && x8 && x6 && ~x11 && ~x12 && ~x10 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y38 = 1'b1;	y46 = 1'b1;	
							nx_state = s749;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && x8 && ~x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s750;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && ~x8 && x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s750;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && ~x8 && ~x7 && x6 && x11 && x12 && x10 )
						begin
							y40 = 1'b1;	
							nx_state = s751;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && ~x8 && ~x7 && x6 && x11 && x12 && ~x10 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s752;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && ~x8 && ~x7 && x6 && x11 && ~x12 && x10 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && ~x8 && ~x7 && x6 && x11 && ~x12 && ~x10 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y35 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s749;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && ~x8 && ~x7 && x6 && ~x11 && x12 && x10 )
						begin
							y42 = 1'b1;	
							nx_state = s754;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && ~x8 && ~x7 && x6 && ~x11 && x12 && ~x10 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y33 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s749;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && ~x8 && ~x7 && x6 && ~x11 && ~x12 && x10 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && ~x8 && ~x7 && x6 && ~x11 && ~x12 && ~x10 )
						begin
							y44 = 1'b1;	
							nx_state = s755;
						end
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 && ~x8 && ~x7 && ~x6 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s756;
						end
					else if( x69 && x70 && ~x64 && x63 && x11 && x4 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x70 && ~x64 && x63 && x11 && ~x4 )
						begin
							y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s757;
						end
					else if( x69 && x70 && ~x64 && x63 && ~x11 && x4 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( x69 && x70 && ~x64 && x63 && ~x11 && ~x4 && x7 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x69 && x70 && ~x64 && x63 && ~x11 && ~x4 && ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x67 && x23 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x67 && ~x23 && x24 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x67 && ~x23 && x24 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x67 && ~x23 && x24 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x69 && x70 && ~x64 && ~x63 && x67 && ~x23 && x24 && ~x20 )
						nx_state = s1;
					else if( x69 && x70 && ~x64 && ~x63 && x67 && ~x23 && ~x24 && x11 && x12 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x67 && ~x23 && ~x24 && x11 && ~x12 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x67 && ~x23 && ~x24 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x69 && x70 && ~x64 && ~x63 && x67 && ~x23 && ~x24 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x64 && ~x63 && ~x67 && x29 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x64 && ~x63 && ~x67 && x29 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x64 && ~x63 && ~x67 && x29 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x69 && x70 && ~x64 && ~x63 && ~x67 && x29 && ~x23 )
						nx_state = s1;
					else if( x69 && x70 && ~x64 && ~x63 && ~x67 && ~x29 )
						begin
							y8 = 1'b1;	
							nx_state = s373;
						end
					else if( x69 && ~x70 && x65 && x67 && x21 && x68 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x69 && ~x70 && x65 && x67 && x21 && x68 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x69 && ~x70 && x65 && x67 && x21 && x68 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && x21 && x68 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && x21 && ~x68 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && x67 && x21 && ~x68 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && x67 && x21 && ~x68 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && x21 && ~x68 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x68 && x23 && x22 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x68 && x23 && x22 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x68 && x23 && x22 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x68 && x23 && x22 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x68 && x23 && ~x22 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x68 && x23 && ~x22 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x68 && x23 && ~x22 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x68 && x23 && ~x22 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x68 && ~x23 && x8 && x22 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x68 && ~x23 && x8 && x22 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x68 && ~x23 && x8 && x22 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x68 && ~x23 && x8 && ~x22 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x68 && ~x23 && x8 && ~x22 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x68 && ~x23 && x8 && ~x22 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x68 && ~x23 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x68 && x22 && x19 && x18 && x11 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x68 && x22 && x19 && x18 && ~x11 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x68 && x22 && x19 && x18 && ~x11 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x68 && x22 && x19 && x18 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x68 && x22 && x19 && x18 && ~x11 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x68 && x22 && x19 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x68 && x22 && ~x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x68 && x22 && ~x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x68 && x22 && ~x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x68 && x22 && ~x19 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x68 && ~x22 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x68 && ~x22 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x68 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x68 && ~x22 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x21 && x23 && x22 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x21 && x23 && x22 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x21 && x23 && x22 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x21 && x23 && ~x22 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x21 && x23 && ~x22 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x21 && x23 && ~x22 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x21 && x23 && ~x22 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x21 && ~x23 && x18 && x14 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x21 && ~x23 && x18 && x14 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x21 && ~x23 && x18 && ~x14 && x13 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x21 && ~x23 && x18 && ~x14 && x13 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x21 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x21 && ~x23 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && x68 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x68 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x68 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x68 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x68 && x62 && ~x61 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && x21 && x17 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && x21 && x17 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && x21 && x17 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && x21 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && x22 && ~x8 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && ~x22 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x67 && ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x22 && x21 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x22 && ~x21 && x16 && x12 && x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x22 && ~x21 && x16 && x12 && ~x19 && x18 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x22 && ~x21 && x16 && x12 && ~x19 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x22 && ~x21 && x16 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x22 && ~x21 && ~x16 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x22 )
						nx_state = s1;
					else if( ~x69 && x70 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && x70 && ~x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x69 && ~x70 && x45 && x12 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && x45 && x12 && ~x1 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x69 && ~x70 && x45 && ~x12 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && ~x70 && ~x45 && x10 && x46 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && ~x70 && ~x45 && x10 && ~x46 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x70 && ~x45 && x10 && ~x46 && ~x1 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x10 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else nx_state = s95;
				s96 : if( x69 && x21 )
						begin
							y10 = 1'b1;	
							nx_state = s405;
						end
					else if( x69 && ~x21 && x19 && x16 && x10 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( x69 && ~x21 && x19 && x16 && ~x10 )
						begin
							y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s233;
						end
					else if( x69 && ~x21 && x19 && ~x16 && x17 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x21 && x19 && ~x16 && ~x17 )
						begin
							y5 = 1'b1;	y17 = 1'b1;	
							nx_state = s721;
						end
					else if( x69 && ~x21 && ~x19 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	
							nx_state = s758;
						end
					else if( ~x69 && x10 && x12 && x70 && x64 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( ~x69 && x10 && x12 && x70 && ~x64 )
						nx_state = s1;
					else if( ~x69 && x10 && x12 && ~x70 )
						nx_state = s1;
					else if( ~x69 && x10 && ~x12 && x1 && x2 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && x10 && ~x12 && x1 && ~x2 && x70 && x64 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( ~x69 && x10 && ~x12 && x1 && ~x2 && x70 && ~x64 )
						nx_state = s1;
					else if( ~x69 && x10 && ~x12 && x1 && ~x2 && ~x70 )
						nx_state = s1;
					else if( ~x69 && x10 && ~x12 && ~x1 && x70 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( ~x69 && x10 && ~x12 && ~x1 && ~x70 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s733;
						end
					else if( ~x69 && ~x10 && x11 && x1 && x70 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s759;
						end
					else if( ~x69 && ~x10 && x11 && x1 && ~x70 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && ~x10 && x11 && ~x1 && x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && ~x10 && x11 && ~x1 && ~x3 && x70 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && ~x10 && x11 && ~x1 && ~x3 && ~x70 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x10 && ~x11 && x12 && x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && ~x10 && ~x11 && x12 && ~x3 && x70 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s201;
						end
					else if( ~x69 && ~x10 && ~x11 && x12 && ~x3 && ~x70 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( ~x69 && ~x10 && ~x11 && ~x12 && x6 && x70 && x64 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( ~x69 && ~x10 && ~x11 && ~x12 && x6 && x70 && ~x64 )
						nx_state = s1;
					else if( ~x69 && ~x10 && ~x11 && ~x12 && x6 && ~x70 )
						nx_state = s1;
					else if( ~x69 && ~x10 && ~x11 && ~x12 && ~x6 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else nx_state = s96;
				s97 : if( x65 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x65 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	
							nx_state = s594;
						end
					else nx_state = s97;
				s98 : if( x70 && x63 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x70 && x63 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x70 && x63 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x70 && x63 && ~x1 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x63 && x64 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x63 && x64 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x66 && x67 && x11 && x12 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x70 && ~x63 && ~x64 && x66 && x67 && x11 && ~x12 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x70 && ~x63 && ~x64 && x66 && x67 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x66 && x67 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x66 && ~x67 && x28 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x63 && ~x64 && x66 && ~x67 && x28 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x63 && ~x64 && x66 && ~x67 && x28 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x66 && ~x67 && x28 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x66 && ~x67 && ~x28 )
						begin
							y8 = 1'b1;	
							nx_state = s642;
						end
					else if( x70 && ~x63 && ~x64 && ~x66 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && ~x63 && ~x64 && ~x66 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && ~x63 && ~x64 && ~x66 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && ~x66 && ~x15 )
						nx_state = s1;
					else if( ~x70 && x66 && x67 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x67 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x70 && x66 && ~x67 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x70 && x66 && ~x67 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x67 && ~x4 )
						nx_state = s1;
					else if( ~x70 && ~x66 && x24 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x66 && ~x24 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s761;
						end
					else nx_state = s98;
				s99 : if( x69 )
						nx_state = s1;
					else if( ~x69 && x42 && x43 && x13 && x10 && x4 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x69 && x42 && x43 && x13 && x10 && ~x4 )
						nx_state = s99;
					else if( ~x69 && x42 && x43 && x13 && ~x10 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x42 && x43 && x13 && ~x10 && ~x3 && x33 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && x42 && x43 && x13 && ~x10 && ~x3 && ~x33 )
						nx_state = s99;
					else if( ~x69 && x42 && x43 && ~x13 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x42 && x43 && ~x13 && ~x3 && x33 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && x42 && x43 && ~x13 && ~x3 && ~x33 )
						nx_state = s99;
					else if( ~x69 && x42 && ~x43 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x42 && ~x43 && ~x3 && x33 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && x42 && ~x43 && ~x3 && ~x33 )
						nx_state = s99;
					else if( ~x69 && ~x42 && x12 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && ~x42 && x12 && ~x3 && x33 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && ~x42 && x12 && ~x3 && ~x33 )
						nx_state = s99;
					else if( ~x69 && ~x42 && ~x12 && x44 && x45 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && ~x42 && ~x12 && x44 && x45 && ~x3 && x33 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && ~x42 && ~x12 && x44 && x45 && ~x3 && ~x33 )
						nx_state = s99;
					else if( ~x69 && ~x42 && ~x12 && x44 && ~x45 && x41 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( ~x69 && ~x42 && ~x12 && x44 && ~x45 && ~x41 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && ~x42 && ~x12 && x44 && ~x45 && ~x41 && ~x3 && x33 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && ~x42 && ~x12 && x44 && ~x45 && ~x41 && ~x3 && ~x33 )
						nx_state = s99;
					else if( ~x69 && ~x42 && ~x12 && ~x44 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && ~x42 && ~x12 && ~x44 && ~x3 && x33 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && ~x42 && ~x12 && ~x44 && ~x3 && ~x33 )
						nx_state = s99;
					else nx_state = s99;
				s100 : if( x63 && x62 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x63 && ~x62 && x15 && x8 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x63 && ~x62 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x63 && ~x62 && ~x15 && x16 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x63 && ~x62 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s299;
						end
					else if( ~x63 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else nx_state = s100;
				s101 : if( x66 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( ~x66 && x26 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x66 && ~x26 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else nx_state = s101;
				s102 : if( x64 )
						nx_state = s1;
					else if( ~x64 && x63 && x18 && x15 && x8 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x64 && x63 && x18 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x64 && x63 && x18 && ~x15 && x16 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x64 && x63 && x18 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s299;
						end
					else if( ~x64 && x63 && ~x18 )
						begin
							y31 = 1'b1;	
							nx_state = s164;
						end
					else if( ~x64 && ~x63 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else nx_state = s102;
				s103 : if( x70 && x62 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x70 && x62 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x70 && x62 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( x70 && x62 && ~x27 )
						nx_state = s1;
					else if( x70 && ~x62 && x64 && x63 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x70 && ~x62 && x64 && x63 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x70 && ~x62 && x64 && x63 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && x64 && x63 && ~x14 )
						nx_state = s1;
					else if( x70 && ~x62 && x64 && ~x63 && x65 && x67 )
						nx_state = s1;
					else if( x70 && ~x62 && x64 && ~x63 && x65 && ~x67 && x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x70 && ~x62 && x64 && ~x63 && x65 && ~x67 && x10 && ~x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x70 && ~x62 && x64 && ~x63 && x65 && ~x67 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x62 && x64 && ~x63 && x65 && ~x67 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x62 && x64 && ~x63 && ~x65 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && x64 && ~x63 && ~x65 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && x64 && ~x63 && ~x65 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && x64 && ~x63 && ~x65 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x64 && x63 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x70 && ~x62 && ~x64 && x63 && ~x15 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && ~x64 && ~x63 && x21 && x22 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( x70 && ~x62 && ~x64 && ~x63 && x21 && ~x22 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( x70 && ~x62 && ~x64 && ~x63 && x21 && ~x22 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x64 && ~x63 && ~x21 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( x70 && ~x62 && ~x64 && ~x63 && ~x21 && ~x23 )
						nx_state = s1;
					else if( ~x70 && x63 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x70 && ~x63 && x62 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x70 && ~x63 && ~x62 && x64 && x16 && x8 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x63 && ~x62 && x64 && x16 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && ~x63 && ~x62 && x64 && ~x16 && x4 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x70 && ~x63 && ~x62 && x64 && ~x16 && ~x4 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s299;
						end
					else if( ~x70 && ~x63 && ~x62 && ~x64 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x70 && ~x63 && ~x62 && ~x64 && x15 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && ~x63 && ~x62 && ~x64 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( ~x70 && ~x63 && ~x62 && ~x64 && ~x15 && ~x16 && x14 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s299;
						end
					else if( ~x70 && ~x63 && ~x62 && ~x64 && ~x15 && ~x16 && ~x14 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s295;
						end
					else nx_state = s103;
				s104 : if( x69 && x70 && x62 && x24 && x2 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && x70 && x62 && x24 && x2 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x69 && x70 && x62 && x24 && ~x2 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x69 && x70 && x62 && ~x24 && x2 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( x69 && x70 && x62 && ~x24 && ~x2 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( x69 && x70 && x62 && ~x24 && ~x2 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x69 && x70 && ~x62 && x63 && x64 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && x64 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x63 && ~x64 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s328;
						end
					else if( x69 && x70 && ~x62 && ~x63 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && x65 && x21 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && x65 && ~x21 && x22 && x23 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && x65 && ~x21 && x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && x65 && ~x21 && ~x22 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x65 && x67 && x64 && x63 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x65 && x67 && x64 && ~x63 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x67 && ~x64 && x63 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && ~x65 && x67 && ~x64 && ~x63 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && x21 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x23 && x22 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x23 && x22 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x23 && x22 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x23 && x22 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && x23 && ~x22 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x67 && ~x21 && ~x23 )
						nx_state = s1;
					else if( ~x69 && x70 && x15 && x3 && x11 && x2 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s698;
						end
					else if( ~x69 && x70 && x15 && x3 && x11 && ~x2 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && x3 && ~x11 && x4 && x12 && x13 && x2 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( ~x69 && x70 && x15 && x3 && ~x11 && x4 && x12 && x13 && ~x2 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && x3 && ~x11 && x4 && x12 && ~x13 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && x3 && ~x11 && x4 && ~x12 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && x3 && ~x11 && ~x4 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && ~x3 && x4 && x11 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s762;
						end
					else if( ~x69 && x70 && x15 && ~x3 && x4 && x11 && ~x2 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && ~x3 && x4 && ~x11 && x12 && x13 && x14 && x2 )
						begin
							y13 = 1'b1;	
							nx_state = s763;
						end
					else if( ~x69 && x70 && x15 && ~x3 && x4 && ~x11 && x12 && x13 && x14 && ~x2 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && ~x3 && x4 && ~x11 && x12 && x13 && ~x14 && x2 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s764;
						end
					else if( ~x69 && x70 && x15 && ~x3 && x4 && ~x11 && x12 && x13 && ~x14 && ~x2 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && ~x3 && x4 && ~x11 && x12 && ~x13 && x2 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s765;
						end
					else if( ~x69 && x70 && x15 && ~x3 && x4 && ~x11 && x12 && ~x13 && ~x2 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && ~x3 && x4 && ~x11 && ~x12 && x2 )
						begin
							y10 = 1'b1;	
							nx_state = s766;
						end
					else if( ~x69 && x70 && x15 && ~x3 && x4 && ~x11 && ~x12 && ~x2 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && x5 && x6 && x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s767;
						end
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && x5 && x6 && ~x2 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && x5 && ~x6 && x7 && x8 && x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s767;
						end
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && x5 && ~x6 && x7 && x8 && ~x2 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && x5 && ~x6 && x7 && ~x8 && x2 )
						begin
							y2 = 1'b1;	
							nx_state = s768;
						end
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && x5 && ~x6 && x7 && ~x8 && ~x2 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && x8 && x2 )
						begin
							y2 = 1'b1;	
							nx_state = s768;
						end
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && x8 && ~x2 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && ~x8 && x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s767;
						end
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && x5 && ~x6 && ~x7 && ~x8 && ~x2 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && ~x5 && x6 && x7 && x9 && x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s767;
						end
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && ~x5 && x6 && x7 && x9 && ~x2 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && ~x5 && x6 && x7 && ~x9 && x2 )
						begin
							y2 = 1'b1;	
							nx_state = s768;
						end
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && ~x5 && x6 && x7 && ~x9 && ~x2 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && x9 && x2 )
						begin
							y2 = 1'b1;	
							nx_state = s768;
						end
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && x9 && ~x2 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && ~x9 && x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s767;
						end
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && ~x5 && x6 && ~x7 && ~x9 && ~x2 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && x10 && x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s767;
						end
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && x10 && ~x2 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && ~x10 && x2 )
						begin
							y2 = 1'b1;	
							nx_state = s768;
						end
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && x7 && ~x10 && ~x2 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && x10 && x2 )
						begin
							y2 = 1'b1;	
							nx_state = s768;
						end
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && x10 && ~x2 )
						nx_state = s104;
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && ~x10 && x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s767;
						end
					else if( ~x69 && x70 && x15 && ~x3 && ~x4 && ~x5 && ~x6 && ~x7 && ~x10 && ~x2 )
						nx_state = s104;
					else if( ~x69 && x70 && ~x15 && x7 )
						begin
							y13 = 1'b1;	
							nx_state = s769;
						end
					else if( ~x69 && x70 && ~x15 && ~x7 && x9 )
						begin
							y13 = 1'b1;	
							nx_state = s769;
						end
					else if( ~x69 && x70 && ~x15 && ~x7 && ~x9 && x10 && x6 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x69 && x70 && ~x15 && ~x7 && ~x9 && x10 && ~x6 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s770;
						end
					else if( ~x69 && x70 && ~x15 && ~x7 && ~x9 && ~x10 && x11 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s767;
						end
					else if( ~x69 && x70 && ~x15 && ~x7 && ~x9 && ~x10 && ~x11 )
						nx_state = s104;
					else if( ~x69 && ~x70 && x44 && x45 && x26 && x42 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x26 && ~x42 && x15 && x40 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x26 && ~x42 && x15 && ~x40 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x26 && ~x42 && ~x15 && x34 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x26 && ~x42 && ~x15 && ~x34 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x26 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x2 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x70 && ~x44 && x10 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 && x2 && x11 && x13 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 && x2 && x11 && ~x13 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 && x2 && ~x11 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 && x2 && ~x11 && ~x12 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 && ~x2 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else nx_state = s104;
				s105 : if( x70 && x62 && x66 && x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x70 && x62 && x66 && ~x6 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x70 && x62 && ~x66 && x17 && x18 && x5 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x70 && x62 && ~x66 && x17 && x18 && ~x5 && x6 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x70 && x62 && ~x66 && x17 && x18 && ~x5 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x70 && x62 && ~x66 && x17 && ~x18 && x9 && x10 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x70 && x62 && ~x66 && x17 && ~x18 && x9 && ~x10 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x70 && x62 && ~x66 && x17 && ~x18 && ~x9 && x6 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x70 && x62 && ~x66 && x17 && ~x18 && ~x9 && ~x6 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x70 && x62 && ~x66 && ~x17 && x18 )
						nx_state = s1;
					else if( x70 && x62 && ~x66 && ~x17 && ~x18 && x6 && x7 && x2 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x70 && x62 && ~x66 && ~x17 && ~x18 && x6 && x7 && x2 && ~x3 && x4 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x70 && x62 && ~x66 && ~x17 && ~x18 && x6 && x7 && x2 && ~x3 && ~x4 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x70 && x62 && ~x66 && ~x17 && ~x18 && x6 && x7 && ~x2 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	
							nx_state = s20;
						end
					else if( x70 && x62 && ~x66 && ~x17 && ~x18 && x6 && ~x7 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x70 && x62 && ~x66 && ~x17 && ~x18 && x6 && ~x7 && ~x8 && x2 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x70 && x62 && ~x66 && ~x17 && ~x18 && x6 && ~x7 && ~x8 && x2 && ~x3 && x4 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x70 && x62 && ~x66 && ~x17 && ~x18 && x6 && ~x7 && ~x8 && x2 && ~x3 && ~x4 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x70 && x62 && ~x66 && ~x17 && ~x18 && x6 && ~x7 && ~x8 && ~x2 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	
							nx_state = s20;
						end
					else if( x70 && x62 && ~x66 && ~x17 && ~x18 && ~x6 && x2 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x70 && x62 && ~x66 && ~x17 && ~x18 && ~x6 && ~x2 )
						nx_state = s1;
					else if( x70 && ~x62 && x63 && x67 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s18;
						end
					else if( x70 && ~x62 && x63 && ~x67 && x29 && x5 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x70 && ~x62 && x63 && ~x67 && x29 && x5 && ~x4 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x70 && ~x62 && x63 && ~x67 && x29 && ~x5 && x4 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x70 && ~x62 && x63 && ~x67 && x29 && ~x5 && ~x4 )
						begin
							y8 = 1'b1;	
							nx_state = s568;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && x30 && x4 && x31 && x15 && x5 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && x30 && x4 && x31 && x15 && ~x5 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && x30 && x4 && x31 && ~x15 && x16 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && x30 && x4 && x31 && ~x15 && ~x16 && x5 )
						begin
							y47 = 1'b1;	
							nx_state = s675;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && x30 && x4 && x31 && ~x15 && ~x16 && ~x5 )
						begin
							y48 = 1'b1;	
							nx_state = s676;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && x30 && x4 && ~x31 && x5 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && x30 && x4 && ~x31 && ~x5 )
						begin
							y19 = 1'b1;	
							nx_state = s13;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && x30 && ~x4 && x5 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && x30 && ~x4 && ~x5 && x31 && x15 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && x30 && ~x4 && ~x5 && x31 && ~x15 && x16 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && x30 && ~x4 && ~x5 && x31 && ~x15 && ~x16 )
						begin
							y35 = 1'b1;	
							nx_state = s718;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && x30 && ~x4 && ~x5 && ~x31 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && ~x30 && x5 && x31 && x4 && x13 )
						begin
							y29 = 1'b1;	
							nx_state = s771;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && ~x30 && x5 && x31 && x4 && ~x13 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && ~x30 && x5 && x31 && ~x4 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && ~x30 && x5 && ~x31 && x4 && x8 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && ~x30 && x5 && ~x31 && x4 && ~x8 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && ~x30 && x5 && ~x31 && ~x4 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && ~x30 && ~x5 && x31 && x4 && x8 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && ~x30 && ~x5 && x31 && x4 && ~x8 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && ~x30 && ~x5 && x31 && ~x4 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && ~x30 && ~x5 && ~x31 && x4 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && ~x30 && ~x5 && ~x31 && ~x4 && x9 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && ~x30 && ~x5 && ~x31 && ~x4 && ~x9 && x7 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x29 && ~x30 && ~x5 && ~x31 && ~x4 && ~x9 && ~x7 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x65 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && x5 && x18 && x19 && x12 )
						begin
							y54 = 1'b1;	
							nx_state = s772;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && x5 && x18 && x19 && ~x12 )
						begin
							y55 = 1'b1;	
							nx_state = s773;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && x5 && x18 && ~x19 && x12 && x6 )
						begin
							y50 = 1'b1;	y52 = 1'b1;	
							nx_state = s774;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && x5 && x18 && ~x19 && x12 && ~x6 && x16 )
						begin
							y51 = 1'b1;	
							nx_state = s655;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && x5 && x18 && ~x19 && x12 && ~x6 && ~x16 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && x5 && x18 && ~x19 && x12 && ~x6 && ~x16 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && x5 && x18 && ~x19 && x12 && ~x6 && ~x16 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && x5 && x18 && ~x19 && x12 && ~x6 && ~x16 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && x5 && x18 && ~x19 && ~x12 && x6 )
						begin
							y6 = 1'b1;	
							nx_state = s368;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && x5 && x18 && ~x19 && ~x12 && ~x6 && x15 )
						begin
							y51 = 1'b1;	
							nx_state = s655;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && x5 && x18 && ~x19 && ~x12 && ~x6 && ~x15 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && x5 && x18 && ~x19 && ~x12 && ~x6 && ~x15 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && x5 && x18 && ~x19 && ~x12 && ~x6 && ~x15 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && x5 && x18 && ~x19 && ~x12 && ~x6 && ~x15 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && x5 && ~x18 && x19 )
						begin
							y27 = 1'b1;	y39 = 1'b1;	y40 = 1'b1;	
							nx_state = s284;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && x5 && ~x18 && ~x19 && x6 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && x5 && ~x18 && ~x19 && ~x6 )
						begin
							y22 = 1'b1;	
							nx_state = s130;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && x19 && x6 && x12 && x11 )
						begin
							y46 = 1'b1;	
							nx_state = s775;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && x19 && x6 && x12 && ~x11 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && x19 && x6 && x12 && ~x11 && x9 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && x19 && x6 && x12 && ~x11 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && x19 && x6 && ~x12 && x10 )
						begin
							y46 = 1'b1;	
							nx_state = s775;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && x19 && x6 && ~x12 && ~x10 && x9 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && x19 && x6 && ~x12 && ~x10 && x9 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && x19 && x6 && ~x12 && ~x10 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && x19 && ~x6 && x12 )
						begin
							y59 = 1'b1;	y61 = 1'b1;	
							nx_state = s284;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && x19 && ~x6 && ~x12 )
						begin
							y56 = 1'b1;	y57 = 1'b1;	
							nx_state = s284;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && ~x19 && x6 && x12 && x14 )
						begin
							y51 = 1'b1;	
							nx_state = s655;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && ~x19 && x6 && x12 && ~x14 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && ~x19 && x6 && x12 && ~x14 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && ~x19 && x6 && x12 && ~x14 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && ~x19 && x6 && x12 && ~x14 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && ~x19 && x6 && ~x12 && x13 )
						begin
							y51 = 1'b1;	
							nx_state = s655;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && ~x19 && x6 && ~x12 && ~x13 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && ~x19 && x6 && ~x12 && ~x13 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && ~x19 && x6 && ~x12 && ~x13 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && ~x19 && x6 && ~x12 && ~x13 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && x18 && ~x19 && ~x6 )
						begin
							y51 = 1'b1;	
							nx_state = s655;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && ~x18 && x19 && x12 && x6 )
						begin
							y44 = 1'b1;	
							nx_state = s755;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && ~x18 && x19 && x12 && ~x6 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && ~x18 && x19 && ~x12 && x6 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && ~x18 && x19 && ~x12 && ~x6 )
						begin
							y42 = 1'b1;	
							nx_state = s754;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x7 && ~x5 && ~x18 && ~x19 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && ~x7 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x3 && x24 && x23 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x3 && x24 && x23 && ~x7 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x3 && x24 && ~x23 && x5 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x3 && x24 && ~x23 && x5 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x3 && x24 && ~x23 && x5 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && x3 && x24 && ~x23 && x5 && ~x20 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && x3 && x24 && ~x23 && ~x5 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x3 && ~x24 && x5 && x11 && x12 && x23 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x3 && ~x24 && x5 && x11 && x12 && ~x23 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x3 && ~x24 && x5 && x11 && ~x12 && x13 && x23 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x3 && ~x24 && x5 && x11 && ~x12 && x13 && ~x23 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x3 && ~x24 && x5 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && x3 && ~x24 && x5 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && x3 && ~x24 && ~x5 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x66 && x65 && x15 && x16 && x12 && x10 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && x66 && x65 && x15 && x16 && x12 && ~x10 && x20 && x13 && x11 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s358;
						end
					else if( ~x70 && x66 && x65 && x15 && x16 && x12 && ~x10 && x20 && x13 && ~x11 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( ~x70 && x66 && x65 && x15 && x16 && x12 && ~x10 && x20 && ~x13 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x66 && x65 && x15 && x16 && x12 && ~x10 && x20 && ~x13 && x19 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && x15 && x16 && x12 && ~x10 && x20 && ~x13 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && x15 && x16 && x12 && ~x10 && ~x20 && x21 && x11 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s358;
						end
					else if( ~x70 && x66 && x65 && x15 && x16 && x12 && ~x10 && ~x20 && x21 && ~x11 && x13 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s426;
						end
					else if( ~x70 && x66 && x65 && x15 && x16 && x12 && ~x10 && ~x20 && x21 && ~x11 && ~x13 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x66 && x65 && x15 && x16 && x12 && ~x10 && ~x20 && x21 && ~x11 && ~x13 && x19 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && x15 && x16 && x12 && ~x10 && ~x20 && x21 && ~x11 && ~x13 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && x15 && x16 && x12 && ~x10 && ~x20 && ~x21 && x13 && x11 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s358;
						end
					else if( ~x70 && x66 && x65 && x15 && x16 && x12 && ~x10 && ~x20 && ~x21 && x13 && ~x11 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( ~x70 && x66 && x65 && x15 && x16 && x12 && ~x10 && ~x20 && ~x21 && ~x13 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x66 && x65 && x15 && x16 && x12 && ~x10 && ~x20 && ~x21 && ~x13 && x19 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && x15 && x16 && x12 && ~x10 && ~x20 && ~x21 && ~x13 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && x15 && x16 && ~x12 && x10 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && x66 && x65 && x15 && x16 && ~x12 && ~x10 && x11 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s600;
						end
					else if( ~x70 && x66 && x65 && x15 && x16 && ~x12 && ~x10 && ~x11 && x14 && x20 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( ~x70 && x66 && x65 && x15 && x16 && ~x12 && ~x10 && ~x11 && x14 && ~x20 && x21 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s426;
						end
					else if( ~x70 && x66 && x65 && x15 && x16 && ~x12 && ~x10 && ~x11 && x14 && ~x20 && ~x21 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( ~x70 && x66 && x65 && x15 && x16 && ~x12 && ~x10 && ~x11 && ~x14 && x19 && x13 && x20 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x66 && x65 && x15 && x16 && ~x12 && ~x10 && ~x11 && ~x14 && x19 && x13 && ~x20 && x21 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x66 && x65 && x15 && x16 && ~x12 && ~x10 && ~x11 && ~x14 && x19 && x13 && ~x20 && ~x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x66 && x65 && x15 && x16 && ~x12 && ~x10 && ~x11 && ~x14 && x19 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && x15 && x16 && ~x12 && ~x10 && ~x11 && ~x14 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && x15 && ~x16 && x10 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && x10 && ~x2 && x20 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && x10 && ~x2 && x20 && ~x4 && x11 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && x10 && ~x2 && x20 && ~x4 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s601;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && x10 && ~x2 && x20 && ~x4 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s776;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && x10 && ~x2 && ~x20 && x21 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && x10 && ~x2 && ~x20 && x21 && ~x3 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && x10 && ~x2 && ~x20 && x21 && ~x3 && ~x11 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s601;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && x10 && ~x2 && ~x20 && x21 && ~x3 && ~x11 && ~x12 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s606;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && x10 && ~x2 && ~x20 && ~x21 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && x10 && ~x2 && ~x20 && ~x21 && ~x4 && x11 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && x10 && ~x2 && ~x20 && ~x21 && ~x4 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s601;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && x10 && ~x2 && ~x20 && ~x21 && ~x4 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s776;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && ~x10 && x11 && x20 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && ~x10 && x11 && ~x20 && x21 && x12 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && ~x10 && x11 && ~x20 && x21 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s776;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && ~x10 && x11 && ~x20 && ~x21 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && ~x10 && ~x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && ~x10 && ~x11 && ~x2 && x20 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && ~x10 && ~x11 && ~x2 && x20 && ~x4 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s777;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && ~x10 && ~x11 && ~x2 && x20 && ~x4 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s602;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && ~x10 && ~x11 && ~x2 && ~x20 && x21 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && ~x10 && ~x11 && ~x2 && ~x20 && x21 && ~x3 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && ~x10 && ~x11 && ~x2 && ~x20 && x21 && ~x3 && ~x12 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s556;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && ~x10 && ~x11 && ~x2 && ~x20 && ~x21 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && ~x10 && ~x11 && ~x2 && ~x20 && ~x21 && ~x4 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s777;
						end
					else if( ~x70 && x66 && x65 && x15 && ~x16 && ~x10 && ~x11 && ~x2 && ~x20 && ~x21 && ~x4 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s602;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && x10 && x12 && x8 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && x10 && x12 && ~x8 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && x10 && x12 && ~x8 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && x10 && x12 && ~x8 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s603;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && x10 && ~x12 && x9 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && x10 && ~x12 && x9 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s778;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && x10 && ~x12 && x9 && ~x2 && ~x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && x10 && ~x12 && ~x9 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && ~x10 && x12 && x7 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && ~x10 && x12 && x7 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && ~x10 && x12 && x7 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s603;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && ~x10 && x12 && ~x7 && x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && ~x10 && x12 && ~x7 && x11 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && ~x10 && x12 && ~x7 && x11 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s603;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && ~x10 && x12 && ~x7 && ~x11 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && ~x10 && ~x12 && x11 && x9 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && ~x10 && ~x12 && x11 && x9 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && ~x10 && ~x12 && x11 && x9 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s603;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && ~x10 && ~x12 && x11 && ~x9 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && ~x10 && ~x12 && ~x11 && x8 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && ~x10 && ~x12 && ~x11 && x8 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && ~x10 && ~x12 && ~x11 && x8 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s603;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && x16 && ~x10 && ~x12 && ~x11 && ~x8 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x15 && x20 && ~x16 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && ~x16 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && x66 && x65 && ~x15 && x20 && ~x16 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s604;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && x10 && x8 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s779;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && x10 && x8 && ~x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && x10 && ~x8 && x12 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && x10 && ~x8 && x12 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && x10 && ~x8 && x12 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && x10 && ~x8 && x12 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && x10 && ~x8 && ~x12 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s779;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && x10 && ~x8 && ~x12 && ~x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && x12 && x11 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && x12 && x11 && ~x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y11 = 1'b1;	
							nx_state = s600;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && x12 && ~x11 && x7 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s779;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && x12 && ~x11 && x7 && ~x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && x12 && ~x11 && ~x7 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && x12 && ~x11 && ~x7 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && x12 && ~x11 && ~x7 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && x12 && ~x11 && ~x7 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && x11 && x9 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s779;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && x11 && x9 && ~x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && x11 && ~x9 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && x11 && ~x9 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && x11 && ~x9 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && x11 && ~x9 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && ~x11 && x8 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && ~x11 && x8 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && ~x11 && x8 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && ~x11 && x8 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && ~x11 && ~x8 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s779;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && ~x11 && ~x8 && ~x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && ~x16 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && ~x16 && ~x3 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && x10 && x12 && x8 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && x10 && x12 && ~x8 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && x10 && x12 && ~x8 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && x10 && x12 && ~x8 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s603;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && x10 && ~x12 && x9 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && x10 && ~x12 && x9 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s778;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && x10 && ~x12 && x9 && ~x2 && ~x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && x10 && ~x12 && ~x9 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && x12 && x7 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && x12 && x7 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && x12 && x7 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s603;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && x12 && ~x7 && x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && x12 && ~x7 && x11 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && x12 && ~x7 && x11 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s603;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && x12 && ~x7 && ~x11 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && ~x12 && x11 && x9 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && ~x12 && x11 && x9 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && ~x12 && x11 && x9 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s603;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && ~x12 && x11 && ~x9 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && ~x12 && ~x11 && x8 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && ~x12 && ~x11 && x8 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && ~x12 && ~x11 && x8 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s603;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && ~x12 && ~x11 && ~x8 )
						nx_state = s1;
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && ~x16 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && ~x16 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && x66 && x65 && ~x15 && ~x20 && ~x21 && ~x16 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s604;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && x15 && x14 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && x15 && x14 && ~x9 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && x15 && ~x14 && x7 && x9 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s296;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && x15 && ~x14 && x7 && ~x9 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s297;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && x15 && ~x14 && ~x7 && x9 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && x15 && ~x14 && ~x7 && x9 && ~x12 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && x15 && ~x14 && ~x7 && x9 && ~x12 && x61 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x65 && x62 && x16 && x15 && ~x14 && ~x7 && x9 && ~x12 && ~x61 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x65 && x62 && x16 && x15 && ~x14 && ~x7 && ~x9 && x13 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && x15 && ~x14 && ~x7 && ~x9 && ~x13 && x61 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && x15 && ~x14 && ~x7 && ~x9 && ~x13 && x61 && ~x12 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x65 && x62 && x16 && x15 && ~x14 && ~x7 && ~x9 && ~x13 && ~x61 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x65 && x62 && x16 && ~x15 && x9 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && ~x15 && x9 && ~x3 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && ~x15 && x9 && ~x3 && ~x4 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && x7 && x11 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && x7 && x11 && ~x3 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && x7 && x11 && ~x3 && ~x4 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && x7 && ~x11 && x3 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && x7 && ~x11 && ~x3 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && x7 && ~x11 && ~x3 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && x7 && ~x11 && ~x3 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && x7 && ~x11 && ~x3 && ~x61 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && ~x7 && x10 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && ~x7 && x10 && ~x3 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && ~x7 && x10 && ~x3 && ~x4 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && ~x7 && ~x10 && x3 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && ~x7 && ~x10 && ~x3 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && ~x7 && ~x10 && ~x3 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && ~x7 && ~x10 && ~x3 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && ~x7 && ~x10 && ~x3 && ~x61 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x65 && x62 && ~x16 && x15 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && x66 && ~x65 && x62 && ~x16 && x15 && ~x7 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( ~x70 && x66 && ~x65 && x62 && ~x16 && x15 && ~x7 && ~x3 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && x66 && ~x65 && x62 && ~x16 && x15 && ~x7 && ~x3 && ~x4 && x8 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x66 && ~x65 && x62 && ~x16 && x15 && ~x7 && ~x3 && ~x4 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && x66 && ~x65 && x62 && ~x16 && ~x15 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( ~x70 && x66 && ~x65 && x62 && ~x16 && ~x15 && ~x3 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && x66 && ~x65 && x62 && ~x16 && ~x15 && ~x3 && ~x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && x66 && ~x65 && ~x62 && x63 && x64 && x17 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x66 && ~x65 && ~x62 && x63 && x64 && x17 && ~x13 && x12 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x66 && ~x65 && ~x62 && x63 && x64 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x65 && ~x62 && x63 && x64 && ~x17 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x65 && ~x62 && x63 && ~x64 && x15 && x8 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x66 && ~x65 && ~x62 && x63 && ~x64 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && x66 && ~x65 && ~x62 && x63 && ~x64 && ~x15 && x16 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x70 && x66 && ~x65 && ~x62 && x63 && ~x64 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s299;
						end
					else if( ~x70 && x66 && ~x65 && ~x62 && ~x63 && x64 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x66 && ~x65 && ~x62 && ~x63 && ~x64 && x6 && x15 && x8 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x66 && ~x65 && ~x62 && ~x63 && ~x64 && x6 && x15 && ~x8 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( ~x70 && x66 && ~x65 && ~x62 && ~x63 && ~x64 && x6 && ~x15 && x16 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x66 && ~x65 && ~x62 && ~x63 && ~x64 && x6 && ~x15 && ~x16 && x14 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s468;
						end
					else if( ~x70 && x66 && ~x65 && ~x62 && ~x63 && ~x64 && x6 && ~x15 && ~x16 && ~x14 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s102;
						end
					else if( ~x70 && x66 && ~x65 && ~x62 && ~x63 && ~x64 && ~x6 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x66 && x65 && x21 && x15 && x9 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x66 && x65 && x21 && x15 && ~x9 && x6 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && ~x66 && x65 && x21 && x15 && ~x9 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && x16 && x9 && x8 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && x16 && x9 && ~x8 && x10 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && x16 && x9 && ~x8 && ~x10 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && x16 && x9 && ~x8 && ~x10 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && x16 && x9 && ~x8 && ~x10 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && x16 && x9 && ~x8 && ~x10 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && x16 && x9 && ~x8 && ~x10 && ~x18 && ~x19 )
						nx_state = s1;
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && x8 && x12 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && x8 && ~x12 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && x8 && ~x12 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && x8 && ~x12 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && x8 && ~x12 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && x8 && ~x12 && ~x18 && ~x19 )
						nx_state = s1;
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && ~x8 && x11 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && ~x8 && ~x11 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && ~x8 && ~x11 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && ~x8 && ~x11 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && ~x8 && ~x11 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && ~x8 && ~x11 && ~x18 && ~x19 )
						nx_state = s1;
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && ~x16 && x6 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s495;
						end
					else if( ~x70 && ~x66 && x65 && x21 && ~x15 && ~x16 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x66 && x65 && ~x21 && x22 && x18 && x14 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x70 && ~x66 && x65 && ~x21 && x22 && x18 && ~x14 && x13 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x70 && ~x66 && x65 && ~x21 && x22 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x66 && x65 && ~x21 && x22 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x66 && x65 && ~x21 && ~x22 && x23 && x15 && x9 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && ~x66 && x65 && ~x21 && ~x22 && x23 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && ~x66 && x65 && ~x21 && ~x22 && x23 && ~x15 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s495;
						end
					else if( ~x70 && ~x66 && x65 && ~x21 && ~x22 && ~x23 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && x20 && x15 && x8 )
						begin
							y2 = 1'b1;	y13 = 1'b1;	
							nx_state = s780;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && x20 && x15 && ~x8 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s781;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && x20 && x15 && ~x8 && ~x6 )
						begin
							y2 = 1'b1;	y13 = 1'b1;	
							nx_state = s782;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && x20 && ~x15 && x16 && x7 && x8 )
						begin
							y2 = 1'b1;	y13 = 1'b1;	
							nx_state = s782;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && x20 && ~x15 && x16 && x7 && ~x8 )
						begin
							y2 = 1'b1;	y13 = 1'b1;	
							nx_state = s780;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && x20 && ~x15 && x16 && ~x7 )
						begin
							y2 = 1'b1;	y13 = 1'b1;	
							nx_state = s780;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && x20 && ~x15 && ~x16 && x6 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && x20 && ~x15 && ~x16 && ~x6 )
						begin
							y2 = 1'b1;	y13 = 1'b1;	
							nx_state = s782;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && x21 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && x14 && x8 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && x14 && ~x8 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s358;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && ~x14 && x7 && x8 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	y20 = 1'b1;	
							nx_state = s781;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && ~x14 && x7 && ~x8 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && ~x14 && ~x7 && x8 && x12 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && x17 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && ~x14 && ~x7 && ~x8 && x13 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && x17 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && x17 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && x7 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && x7 && ~x2 && x3 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && x7 && ~x2 && ~x3 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && ~x7 && x9 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && ~x7 && x9 && ~x2 && x3 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && ~x7 && x9 && ~x2 && ~x3 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && ~x7 && ~x9 && x2 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && ~x7 && ~x9 && ~x2 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && ~x7 && ~x9 && ~x2 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && ~x7 && ~x9 && ~x2 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && ~x7 && ~x9 && ~x2 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && x7 && x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && x7 && x11 && ~x2 && x3 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && x7 && x11 && ~x2 && ~x3 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && x7 && ~x11 && x2 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && x7 && ~x11 && ~x2 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && x7 && ~x11 && ~x2 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && x7 && ~x11 && ~x2 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && x7 && ~x11 && ~x2 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && ~x7 && x10 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && ~x7 && x10 && ~x2 && x3 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && ~x7 && x10 && ~x2 && ~x3 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && x2 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x2 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x2 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x2 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x2 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x16 && x15 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x16 && x15 && ~x7 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x16 && x15 && ~x7 && ~x2 && x3 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x16 && x15 && ~x7 && ~x2 && ~x3 && x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x16 && x15 && ~x7 && ~x2 && ~x3 && ~x8 )
						begin
							y2 = 1'b1;	y13 = 1'b1;	
							nx_state = s780;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x16 && ~x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x16 && ~x15 && ~x2 && x3 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x16 && ~x15 && ~x2 && ~x3 )
						begin
							y7 = 1'b1;	y12 = 1'b1;	
							nx_state = s610;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && x24 && x26 && x11 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s300;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && x24 && x26 && ~x11 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && x24 && x26 && ~x11 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && x24 && x26 && ~x11 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && ~x68 && x24 && x26 && ~x11 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && ~x68 && x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && ~x68 && x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && x26 && x15 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && x26 && ~x15 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && x26 && ~x15 && ~x3 && x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && x26 && ~x15 && ~x3 && ~x1 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x18 && x15 && x10 && x11 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s433;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x18 && x15 && x10 && ~x11 && x12 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s432;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x18 && x15 && x10 && ~x11 && ~x12 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s300;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x18 && x15 && ~x10 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s126;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x18 && ~x15 && x16 && x10 && x12 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x18 && ~x15 && x16 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x18 && ~x15 && x16 && ~x10 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x18 && ~x15 && ~x16 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && ~x18 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && x10 && x12 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && x10 && x12 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && x10 && x12 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && x10 && x12 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && x10 && ~x12 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s304;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && ~x10 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && ~x10 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && ~x10 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && ~x10 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && ~x26 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else nx_state = s105;
				s106 : if( x70 && x63 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x70 && ~x63 && x64 && x10 && ~x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x70 && ~x63 && x64 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && x31 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && x31 && ~x11 && x9 && x8 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && x31 && ~x11 && x9 && x8 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && x31 && ~x11 && x9 && x8 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && x31 && ~x11 && x9 && x8 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && x31 && ~x11 && x9 && ~x8 && x10 && x25 )
						begin
							y29 = 1'b1;	
							nx_state = s771;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && x31 && ~x11 && x9 && ~x8 && x10 && ~x25 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && x31 && ~x11 && x9 && ~x8 && x10 && ~x25 && x23 && ~x24 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && x31 && ~x11 && x9 && ~x8 && x10 && ~x25 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && x31 && ~x11 && x9 && ~x8 && ~x10 && x24 )
						begin
							y29 = 1'b1;	
							nx_state = s771;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && x31 && ~x11 && x9 && ~x8 && ~x10 && ~x24 && x23 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && x31 && ~x11 && x9 && ~x8 && ~x10 && ~x24 && x23 && ~x25 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && x31 && ~x11 && x9 && ~x8 && ~x10 && ~x24 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && x31 && ~x11 && ~x9 && x10 && x8 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s253;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && x31 && ~x11 && ~x9 && x10 && ~x8 )
						begin
							y8 = 1'b1;	
							nx_state = s783;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && x31 && ~x11 && ~x9 && ~x10 && x8 )
						begin
							y10 = 1'b1;	y23 = 1'b1;	
							nx_state = s1;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && x31 && ~x11 && ~x9 && ~x10 && ~x8 )
						begin
							y8 = 1'b1;	
							nx_state = s568;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && ~x31 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && ~x31 && ~x12 && x22 && x9 && x10 && x8 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && ~x31 && ~x12 && x22 && x9 && x10 && ~x8 )
						begin
							y8 = 1'b1;	
							nx_state = s784;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && ~x31 && ~x12 && x22 && x9 && ~x10 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && ~x31 && ~x12 && x22 && x9 && ~x10 && ~x8 )
						begin
							y8 = 1'b1;	
							nx_state = s785;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && ~x31 && ~x12 && x22 && ~x9 && x10 && x8 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && ~x31 && ~x12 && x22 && ~x9 && x10 && ~x8 && x27 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && ~x31 && ~x12 && x22 && ~x9 && x10 && ~x8 && ~x27 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && ~x31 && ~x12 && x22 && ~x9 && ~x10 && x8 )
						begin
							y8 = 1'b1;	
							nx_state = s786;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && ~x31 && ~x12 && x22 && ~x9 && ~x10 && ~x8 && x26 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && ~x31 && ~x12 && x22 && ~x9 && ~x10 && ~x8 && ~x26 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && x30 && ~x31 && ~x12 && ~x22 )
						begin
							y45 = 1'b1;	y47 = 1'b1;	y50 = 1'b1;	
							y60 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							nx_state = s787;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s788;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && x9 && x10 && x8 )
						begin
							y9 = 1'b1;	
							nx_state = s790;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && x9 && x10 && ~x8 && x21 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && x9 && x10 && ~x8 && ~x21 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && x9 && x10 && ~x8 && ~x21 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && x9 && x10 && ~x8 && ~x21 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && x9 && x10 && ~x8 && ~x21 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && x9 && ~x10 && x8 )
						begin
							y3 = 1'b1;	
							nx_state = s789;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && x9 && ~x10 && ~x8 && x18 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && x9 && ~x10 && ~x8 && ~x18 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && x9 && ~x10 && ~x8 && ~x18 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && x9 && ~x10 && ~x8 && ~x18 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && x9 && ~x10 && ~x8 && ~x18 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && ~x9 && x8 && x10 && x19 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && ~x9 && x8 && x10 && ~x19 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && ~x9 && x8 && x10 && ~x19 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && ~x9 && x8 && x10 && ~x19 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && ~x9 && x8 && x10 && ~x19 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && ~x9 && x8 && ~x10 && x20 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && ~x9 && x8 && ~x10 && ~x20 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && ~x9 && x8 && ~x10 && ~x20 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && ~x9 && x8 && ~x10 && ~x20 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && ~x9 && x8 && ~x10 && ~x20 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && x31 && ~x9 && ~x8 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && x22 && ~x31 )
						begin
							y9 = 1'b1;	
							nx_state = s790;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x4 && ~x30 && ~x12 && ~x22 )
						begin
							y45 = 1'b1;	y47 = 1'b1;	y50 = 1'b1;	
							y60 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							nx_state = s787;
						end
					else if( x70 && ~x63 && ~x64 && x65 && ~x4 && x30 )
						begin
							y5 = 1'b1;	
							nx_state = s791;
						end
					else if( x70 && ~x63 && ~x64 && x65 && ~x4 && ~x30 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x70 && ~x63 && ~x64 && ~x65 && x66 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x70 && ~x63 && ~x64 && ~x65 && x66 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x70 && ~x63 && ~x64 && ~x65 && x66 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && ~x65 && x66 && ~x8 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && ~x65 && ~x66 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x63 && ~x64 && ~x65 && ~x66 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x63 && ~x64 && ~x65 && ~x66 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && ~x65 && ~x66 && ~x17 )
						nx_state = s1;
					else if( ~x70 && x65 && x21 && x15 && x9 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x70 && x65 && x21 && x15 && ~x9 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && x65 && x21 && ~x15 && x16 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x70 && x65 && x21 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s333;
						end
					else if( ~x70 && x65 && ~x21 && x23 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && ~x23 && x22 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && ~x22 && x17 && x15 && x9 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && ~x22 && x17 && x15 && ~x9 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && ~x22 && x17 && ~x15 && x16 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && ~x22 && x17 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s495;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && ~x22 && ~x17 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x70 && ~x65 && x62 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x70 && ~x65 && ~x62 && x63 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( ~x70 && ~x65 && ~x62 && ~x63 )
						nx_state = s1;
					else nx_state = s106;
				s107 : if( x21 && x65 )
						nx_state = s1;
					else if( x21 && ~x65 && x16 && x6 && x15 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s181;
						end
					else if( x21 && ~x65 && x16 && x6 && x15 && ~x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s441;
						end
					else if( x21 && ~x65 && x16 && x6 && ~x15 && x10 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x21 && ~x65 && x16 && x6 && ~x15 && ~x10 )
						begin
							y14 = 1'b1;	y16 = 1'b1;	
							nx_state = s492;
						end
					else if( x21 && ~x65 && x16 && ~x6 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s579;
						end
					else if( x21 && ~x65 && ~x16 && x17 && x10 && x6 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s679;
						end
					else if( x21 && ~x65 && ~x16 && x17 && x10 && ~x6 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s579;
						end
					else if( x21 && ~x65 && ~x16 && x17 && ~x10 && x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x21 && ~x65 && ~x16 && x17 && ~x10 && ~x6 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s792;
						end
					else if( x21 && ~x65 && ~x16 && ~x17 && x6 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s680;
						end
					else if( x21 && ~x65 && ~x16 && ~x17 && x6 && ~x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s443;
						end
					else if( x21 && ~x65 && ~x16 && ~x17 && ~x6 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s579;
						end
					else if( ~x21 && x22 && x65 && x23 && x5 && x18 && x15 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( ~x21 && x22 && x65 && x23 && x5 && x18 && ~x15 )
						begin
							y15 = 1'b1;	y20 = 1'b1;	
							nx_state = s665;
						end
					else if( ~x21 && x22 && x65 && x23 && x5 && ~x18 && x19 && x15 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s793;
						end
					else if( ~x21 && x22 && x65 && x23 && x5 && ~x18 && x19 && ~x15 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( ~x21 && x22 && x65 && x23 && x5 && ~x18 && ~x19 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s115;
						end
					else if( ~x21 && x22 && x65 && x23 && ~x5 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( ~x21 && x22 && x65 && ~x23 )
						begin
							y12 = 1'b1;	y19 = 1'b1;	
							nx_state = s794;
						end
					else if( ~x21 && x22 && ~x65 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x21 && ~x22 && x65 && x23 && x19 && x6 && x16 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && ~x22 && x65 && x23 && x19 && x6 && ~x16 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && ~x22 && x65 && x23 && x19 && ~x6 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && x20 && x16 && x6 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s793;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && x20 && x16 && ~x6 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && x20 && ~x16 && x17 && x18 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && x20 && ~x16 && x17 && x18 && ~x6 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && x20 && ~x16 && x17 && ~x18 && x14 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && x20 && ~x16 && x17 && ~x18 && ~x14 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && x20 && ~x16 && ~x17 && x18 && x14 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && x20 && ~x16 && ~x17 && x18 && ~x14 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && x20 && ~x16 && ~x17 && ~x18 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && x20 && ~x16 && ~x17 && ~x18 && ~x6 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && ~x20 && x6 )
						begin
							y12 = 1'b1;	
							nx_state = s245;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && ~x20 && ~x6 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( ~x21 && ~x22 && x65 && ~x23 && x5 && x18 && x15 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( ~x21 && ~x22 && x65 && ~x23 && x5 && x18 && ~x15 )
						begin
							y15 = 1'b1;	y20 = 1'b1;	
							nx_state = s665;
						end
					else if( ~x21 && ~x22 && x65 && ~x23 && x5 && ~x18 && x19 && x15 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s793;
						end
					else if( ~x21 && ~x22 && x65 && ~x23 && x5 && ~x18 && x19 && ~x15 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( ~x21 && ~x22 && x65 && ~x23 && x5 && ~x18 && ~x19 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s115;
						end
					else if( ~x21 && ~x22 && x65 && ~x23 && ~x5 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( ~x21 && ~x22 && ~x65 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s18;
						end
					else nx_state = s107;
				s108 : if( x69 && x65 && x21 )
						nx_state = s1;
					else if( x69 && x65 && ~x21 && x22 && x23 && x18 && x19 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && x18 && x19 && x15 && ~x17 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && x18 && x19 && ~x15 && x16 && x17 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s296;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && x18 && x19 && ~x15 && x16 && ~x17 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y20 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s795;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && x18 && x19 && ~x15 && ~x16 && x8 && x10 && x17 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && x18 && x19 && ~x15 && ~x16 && x8 && x10 && ~x17 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && x18 && x19 && ~x15 && ~x16 && x8 && ~x10 && x11 && x17 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && x18 && x19 && ~x15 && ~x16 && x8 && ~x10 && x11 && ~x17 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && x18 && x19 && ~x15 && ~x16 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x65 && ~x21 && x22 && x23 && x18 && x19 && ~x15 && ~x16 && ~x8 )
						nx_state = s1;
					else if( x69 && x65 && ~x21 && x22 && x23 && x18 && ~x19 && x16 && x15 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && x18 && ~x19 && x16 && ~x15 && x17 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && x18 && ~x19 && x16 && ~x15 && ~x17 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s796;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && x18 && ~x19 && ~x16 && x17 && x15 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && x18 && ~x19 && ~x16 && x17 && ~x15 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s797;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && x18 && ~x19 && ~x16 && ~x17 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s798;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && x18 && ~x19 && ~x16 && ~x17 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && x18 && ~x19 && ~x16 && ~x17 && ~x4 && ~x6 && x15 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s795;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && x18 && ~x19 && ~x16 && ~x17 && ~x4 && ~x6 && ~x15 )
						begin
							y16 = 1'b1;	y20 = 1'b1;	
							nx_state = s795;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && x19 && x15 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s798;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && x19 && x15 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && x19 && x15 && ~x4 && ~x6 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s724;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && x17 && x13 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s798;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && x17 && x13 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && x17 && x13 && ~x4 && ~x6 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s795;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && x17 && ~x13 && x16 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s798;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && x17 && ~x13 && x16 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && x17 && ~x13 && x16 && ~x4 && ~x6 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s795;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && x17 && ~x13 && ~x16 )
						nx_state = s1;
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && ~x17 && x16 && x14 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s798;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && ~x17 && x16 && x14 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && ~x17 && x16 && x14 && ~x4 && ~x6 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s795;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && ~x17 && x16 && ~x14 )
						nx_state = s1;
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && x12 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s798;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && x12 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && x12 && ~x4 && ~x6 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s795;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && ~x12 )
						nx_state = s1;
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && ~x19 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s798;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && ~x19 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x69 && x65 && ~x21 && x22 && x23 && ~x18 && ~x19 && ~x4 && ~x6 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x69 && x65 && ~x21 && x22 && ~x23 && x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( x69 && x65 && ~x21 && x22 && ~x23 && ~x15 && x19 && x18 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( x69 && x65 && ~x21 && x22 && ~x23 && ~x15 && x19 && ~x18 && x8 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && ~x21 && x22 && ~x23 && ~x15 && x19 && ~x18 && x8 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && ~x21 && x22 && ~x23 && ~x15 && x19 && ~x18 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x69 && x65 && ~x21 && x22 && ~x23 && ~x15 && x19 && ~x18 && ~x8 )
						nx_state = s1;
					else if( x69 && x65 && ~x21 && x22 && ~x23 && ~x15 && ~x19 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( x69 && x65 && ~x21 && ~x22 && x23 && x5 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s107;
						end
					else if( x69 && x65 && ~x21 && ~x22 && x23 && ~x5 && x19 && x6 && x16 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( x69 && x65 && ~x21 && ~x22 && x23 && ~x5 && x19 && x6 && ~x16 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x65 && ~x21 && ~x22 && x23 && ~x5 && x19 && ~x6 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( x69 && x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && x20 && x16 && x6 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s793;
						end
					else if( x69 && x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && x20 && x16 && ~x6 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( x69 && x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && x20 && ~x16 && x17 && x18 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( x69 && x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && x20 && ~x16 && x17 && x18 && ~x6 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( x69 && x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && x20 && ~x16 && x17 && ~x18 && x14 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( x69 && x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && x20 && ~x16 && x17 && ~x18 && ~x14 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( x69 && x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && x20 && ~x16 && ~x17 && x18 && x14 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( x69 && x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && x20 && ~x16 && ~x17 && x18 && ~x14 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( x69 && x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && x20 && ~x16 && ~x17 && ~x18 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( x69 && x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && x20 && ~x16 && ~x17 && ~x18 && ~x6 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( x69 && x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && ~x20 && x6 )
						begin
							y12 = 1'b1;	
							nx_state = s245;
						end
					else if( x69 && x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && ~x20 && ~x6 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && x18 && x19 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && x18 && x19 && x15 && ~x17 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && x18 && x19 && ~x15 && x16 && x17 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s296;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && x18 && x19 && ~x15 && x16 && ~x17 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y20 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s795;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && x8 && x10 && x17 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && x8 && x10 && ~x17 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && x8 && ~x10 && x11 && x17 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && x8 && ~x10 && x11 && ~x17 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && ~x8 )
						nx_state = s1;
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && x18 && ~x19 && x16 && x15 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && x18 && ~x19 && x16 && ~x15 && x17 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && x18 && ~x19 && x16 && ~x15 && ~x17 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s796;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && x18 && ~x19 && ~x16 && x17 && x15 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && x18 && ~x19 && ~x16 && x17 && ~x15 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s797;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && x18 && ~x19 && ~x16 && ~x17 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s798;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && x18 && ~x19 && ~x16 && ~x17 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && x18 && ~x19 && ~x16 && ~x17 && ~x4 && ~x6 && x15 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s795;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && x18 && ~x19 && ~x16 && ~x17 && ~x4 && ~x6 && ~x15 )
						begin
							y16 = 1'b1;	y20 = 1'b1;	
							nx_state = s795;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && x15 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s798;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && x15 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && x15 && ~x4 && ~x6 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s724;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && x17 && x13 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s798;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && x17 && x13 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && x17 && x13 && ~x4 && ~x6 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s795;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && x17 && ~x13 && x16 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s798;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && x17 && ~x13 && x16 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && x17 && ~x13 && x16 && ~x4 && ~x6 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s795;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && x17 && ~x13 && ~x16 )
						nx_state = s1;
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && ~x17 && x16 && x14 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s798;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && ~x17 && x16 && x14 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && ~x17 && x16 && x14 && ~x4 && ~x6 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s795;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && ~x17 && x16 && ~x14 )
						nx_state = s1;
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && x12 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s798;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && x12 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && x12 && ~x4 && ~x6 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s795;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && ~x12 )
						nx_state = s1;
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && ~x19 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s798;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && ~x19 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x69 && x65 && ~x21 && ~x22 && ~x23 && ~x18 && ~x19 && ~x4 && ~x6 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x69 && ~x65 && x66 && x21 && x4 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s107;
						end
					else if( x69 && ~x65 && x66 && x21 && ~x4 && x16 && x6 && x15 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s181;
						end
					else if( x69 && ~x65 && x66 && x21 && ~x4 && x16 && x6 && x15 && ~x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s441;
						end
					else if( x69 && ~x65 && x66 && x21 && ~x4 && x16 && x6 && ~x15 && x10 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x65 && x66 && x21 && ~x4 && x16 && x6 && ~x15 && ~x10 )
						begin
							y14 = 1'b1;	y16 = 1'b1;	
							nx_state = s492;
						end
					else if( x69 && ~x65 && x66 && x21 && ~x4 && x16 && ~x6 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s579;
						end
					else if( x69 && ~x65 && x66 && x21 && ~x4 && ~x16 && x17 && x10 && x6 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s679;
						end
					else if( x69 && ~x65 && x66 && x21 && ~x4 && ~x16 && x17 && x10 && ~x6 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s579;
						end
					else if( x69 && ~x65 && x66 && x21 && ~x4 && ~x16 && x17 && ~x10 && x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x69 && ~x65 && x66 && x21 && ~x4 && ~x16 && x17 && ~x10 && ~x6 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s792;
						end
					else if( x69 && ~x65 && x66 && x21 && ~x4 && ~x16 && ~x17 && x6 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s680;
						end
					else if( x69 && ~x65 && x66 && x21 && ~x4 && ~x16 && ~x17 && x6 && ~x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s443;
						end
					else if( x69 && ~x65 && x66 && x21 && ~x4 && ~x16 && ~x17 && ~x6 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s579;
						end
					else if( x69 && ~x65 && x66 && ~x21 && x22 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s443;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x66 && x24 && x26 && x16 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x69 && ~x65 && ~x66 && x24 && x26 && x16 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x69 && ~x65 && ~x66 && x24 && x26 && x16 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x66 && x24 && x26 && x16 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x66 && x24 && x26 && ~x16 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s304;
						end
					else if( x69 && ~x65 && ~x66 && x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( x69 && ~x65 && ~x66 && x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( x69 && ~x65 && ~x66 && x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x66 && x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x66 && ~x24 && x25 && x26 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x65 && ~x66 && ~x24 && x25 && x26 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x65 && ~x66 && ~x24 && x25 && x26 && x19 && ~x14 && ~x13 )
						nx_state = s108;
					else if( x69 && ~x65 && ~x66 && ~x24 && x25 && x26 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x66 && ~x24 && x25 && ~x26 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( x69 && ~x65 && ~x66 && ~x24 && ~x25 && x26 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( x69 && ~x65 && ~x66 && ~x24 && ~x25 && ~x26 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s370;
						end
					else if( ~x69 && x70 && x62 && x64 && x61 && x13 && x23 && x51 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x69 && x70 && x62 && x64 && x61 && x13 && x23 && ~x51 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && x70 && x62 && x64 && x61 && x13 && ~x23 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x69 && x70 && x62 && x64 && x61 && ~x13 && x28 && x35 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x69 && x70 && x62 && x64 && x61 && ~x13 && x28 && x35 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && x62 && x64 && x61 && ~x13 && x28 && ~x35 && x60 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( ~x69 && x70 && x62 && x64 && x61 && ~x13 && x28 && ~x35 && ~x60 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && x62 && x64 && x61 && ~x13 && ~x28 && x6 && x35 )
						begin
							y13 = 1'b1;	
							nx_state = s800;
						end
					else if( ~x69 && x70 && x62 && x64 && x61 && ~x13 && ~x28 && x6 && ~x35 && x60 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( ~x69 && x70 && x62 && x64 && x61 && ~x13 && ~x28 && x6 && ~x35 && ~x60 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && x62 && x64 && x61 && ~x13 && ~x28 && ~x6 && x39 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && x62 && x64 && x61 && ~x13 && ~x28 && ~x6 && ~x39 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x61 && x11 && x10 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x61 && x11 && ~x10 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s759;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x61 && x11 && ~x10 && ~x1 && x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x61 && x11 && ~x10 && ~x1 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x61 && ~x11 && x10 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x61 && ~x11 && ~x10 && x5 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x70 && x62 && x64 && ~x61 && ~x11 && ~x10 && ~x5 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x69 && x70 && x62 && ~x64 && x14 && x13 && x23 && x41 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x69 && x70 && x62 && ~x64 && x14 && x13 && x23 && ~x41 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && x70 && x62 && ~x64 && x14 && x13 && ~x23 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x69 && x70 && x62 && ~x64 && x14 && ~x13 && x28 && x35 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x69 && x70 && x62 && ~x64 && x14 && ~x13 && x28 && x35 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && x62 && ~x64 && x14 && ~x13 && x28 && ~x35 && x15 )
						nx_state = s1;
					else if( ~x69 && x70 && x62 && ~x64 && x14 && ~x13 && x28 && ~x35 && ~x15 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && x62 && ~x64 && x14 && ~x13 && ~x28 && x6 && x35 )
						begin
							y13 = 1'b1;	
							nx_state = s800;
						end
					else if( ~x69 && x70 && x62 && ~x64 && x14 && ~x13 && ~x28 && x6 && ~x35 && x15 )
						nx_state = s1;
					else if( ~x69 && x70 && x62 && ~x64 && x14 && ~x13 && ~x28 && x6 && ~x35 && ~x15 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && x62 && ~x64 && x14 && ~x13 && ~x28 && ~x6 && x39 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && x62 && ~x64 && x14 && ~x13 && ~x28 && ~x6 && ~x39 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( ~x69 && x70 && x62 && ~x64 && ~x14 && x11 && x10 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && x70 && x62 && ~x64 && ~x14 && x11 && ~x10 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s759;
						end
					else if( ~x69 && x70 && x62 && ~x64 && ~x14 && x11 && ~x10 && ~x1 && x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && x70 && x62 && ~x64 && ~x14 && x11 && ~x10 && ~x1 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && x70 && x62 && ~x64 && ~x14 && ~x11 && x10 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x70 && x62 && ~x64 && ~x14 && ~x11 && ~x10 && x5 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x70 && x62 && ~x64 && ~x14 && ~x11 && ~x10 && ~x5 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && x43 && x34 && x44 && x10 && x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s99;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && x43 && x34 && x44 && x10 && ~x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && x43 && x34 && x44 && ~x10 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && x43 && x34 && ~x44 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && x43 && ~x34 && x13 && x41 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && x43 && ~x34 && x13 && ~x41 && x1 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && x43 && ~x34 && x13 && ~x41 && ~x1 && x38 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s801;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && x43 && ~x34 && x13 && ~x41 && ~x1 && ~x38 )
						nx_state = s108;
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && x43 && ~x34 && ~x13 && x1 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && x43 && ~x34 && ~x13 && ~x1 && x38 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s801;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && x43 && ~x34 && ~x13 && ~x1 && ~x38 )
						nx_state = s108;
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && ~x43 && x10 && x44 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && ~x43 && x10 && ~x44 && x45 && x5 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s183;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && ~x43 && x10 && ~x44 && x45 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && ~x43 && x10 && ~x44 && ~x45 && x32 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s181;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && ~x43 && x10 && ~x44 && ~x45 && ~x32 && x3 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && ~x43 && x10 && ~x44 && ~x45 && ~x32 && x3 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && ~x43 && x10 && ~x44 && ~x45 && ~x32 && x3 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && ~x43 && x10 && ~x44 && ~x45 && ~x32 && x3 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && ~x43 && x10 && ~x44 && ~x45 && ~x32 && x3 && x15 && ~x47 && ~x1 )
						nx_state = s108;
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && ~x43 && x10 && ~x44 && ~x45 && ~x32 && x3 && ~x15 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && ~x43 && x10 && ~x44 && ~x45 && ~x32 && ~x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && ~x43 && ~x10 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && ~x43 && ~x10 && ~x34 && x1 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && ~x43 && ~x10 && ~x34 && ~x1 && x38 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s801;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && x42 && ~x43 && ~x10 && ~x34 && ~x1 && ~x38 )
						nx_state = s108;
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && x12 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && x12 && ~x34 && x1 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && x12 && ~x34 && ~x1 && x38 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s801;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && x12 && ~x34 && ~x1 && ~x38 )
						nx_state = s108;
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && ~x12 && x41 && x13 && x14 && x36 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && ~x12 && x41 && x13 && x14 && ~x36 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && ~x12 && x41 && x13 && ~x14 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s183;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && ~x12 && x41 && ~x13 && x45 && x5 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s183;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && ~x12 && x41 && ~x13 && x45 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && ~x12 && x41 && ~x13 && ~x45 && x32 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s181;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && ~x12 && x41 && ~x13 && ~x45 && ~x32 && x3 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && ~x12 && x41 && ~x13 && ~x45 && ~x32 && x3 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && ~x12 && x41 && ~x13 && ~x45 && ~x32 && x3 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && ~x12 && x41 && ~x13 && ~x45 && ~x32 && x3 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && ~x12 && x41 && ~x13 && ~x45 && ~x32 && x3 && x15 && ~x47 && ~x1 )
						nx_state = s108;
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && ~x12 && x41 && ~x13 && ~x45 && ~x32 && x3 && ~x15 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && ~x12 && x41 && ~x13 && ~x45 && ~x32 && ~x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && ~x12 && ~x41 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && ~x12 && ~x41 && ~x34 && x1 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && ~x12 && ~x41 && ~x34 && ~x1 && x38 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s801;
						end
					else if( ~x69 && x70 && ~x62 && x63 && x64 && ~x42 && ~x12 && ~x41 && ~x34 && ~x1 && ~x38 )
						nx_state = s108;
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && x15 && x19 && x28 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && x15 && x19 && x28 && ~x1 && x35 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && x15 && x19 && x28 && ~x1 && ~x35 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && x15 && x19 && ~x28 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && x15 && ~x19 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && ~x15 && x13 && x23 && x48 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && ~x15 && x13 && x23 && ~x48 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && ~x15 && x13 && ~x23 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && ~x15 && ~x13 && x28 && x35 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && ~x15 && ~x13 && x28 && x35 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && ~x15 && ~x13 && x28 && ~x35 && x21 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && ~x15 && ~x13 && x28 && ~x35 && ~x21 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && ~x15 && ~x13 && ~x28 && x6 && x35 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s443;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && ~x15 && ~x13 && ~x28 && x6 && ~x35 && x21 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && ~x15 && ~x13 && ~x28 && x6 && ~x35 && ~x21 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && ~x15 && ~x13 && ~x28 && ~x6 && x39 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && x70 && ~x62 && x63 && ~x64 && ~x15 && ~x13 && ~x28 && ~x6 && ~x39 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && x40 && x19 && x28 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && x40 && x19 && x28 && ~x1 && x35 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && x40 && x19 && x28 && ~x1 && ~x35 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && x40 && x19 && ~x28 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && x40 && ~x19 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && ~x40 && x13 && x23 && x51 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && ~x40 && x13 && x23 && ~x51 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && ~x40 && x13 && ~x23 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && ~x40 && ~x13 && x28 && x35 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && ~x40 && ~x13 && x28 && x35 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && ~x40 && ~x13 && x28 && ~x35 && x41 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && ~x40 && ~x13 && x28 && ~x35 && ~x41 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && ~x40 && ~x13 && ~x28 && x6 && x35 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s443;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && ~x40 && ~x13 && ~x28 && x6 && ~x35 && x41 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && ~x40 && ~x13 && ~x28 && x6 && ~x35 && ~x41 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && ~x40 && ~x13 && ~x28 && ~x6 && x39 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( ~x69 && x70 && ~x62 && ~x63 && ~x40 && ~x13 && ~x28 && ~x6 && ~x39 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s736;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x11 && x10 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x11 && ~x10 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x11 && ~x10 && ~x1 && x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x11 && ~x10 && ~x1 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x11 && x10 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x11 && ~x10 && x5 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x11 && ~x10 && ~x5 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x19 && x28 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x19 && x28 && ~x1 && x15 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x19 && x28 && ~x1 && ~x15 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x19 && ~x28 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x19 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && ~x44 && x10 && x5 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x69 && ~x70 && ~x44 && x10 && ~x5 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s738;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 && ~x1 && x3 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 && ~x1 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else nx_state = s108;
				s109 : if( x70 && x62 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x70 && x62 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x70 && x62 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( x70 && x62 && ~x27 )
						nx_state = s1;
					else if( x70 && ~x62 && x63 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x70 && ~x62 && x63 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x70 && ~x62 && x63 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && x63 && ~x14 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x70 && ~x62 && ~x63 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x70 && ~x62 && ~x63 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x18 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && x67 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && x66 && x67 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && x66 && x67 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && x67 && x22 && ~x17 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && x67 && ~x22 && x18 && x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && x65 && x66 && x67 && ~x22 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && x65 && x66 && x67 && ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && x67 && ~x22 && ~x18 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && ~x67 && x60 && x61 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x65 && x66 && ~x67 && x60 && x61 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x65 && x66 && ~x67 && x60 && x61 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( ~x70 && x65 && x66 && ~x67 && x60 && x61 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( ~x70 && x65 && x66 && ~x67 && x60 && ~x61 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && x66 && ~x67 && x60 && ~x61 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && x66 && ~x67 && x60 && ~x61 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( ~x70 && x65 && x66 && ~x67 && x60 && ~x61 && ~x18 )
						nx_state = s118;
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && x61 && x62 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && x61 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && x61 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && x61 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && x61 && ~x62 && ~x18 )
						nx_state = s118;
					else if( ~x70 && x65 && x66 && ~x67 && ~x60 && ~x61 )
						nx_state = s47;
					else if( ~x70 && x65 && ~x66 && x67 && x21 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( ~x70 && x65 && ~x66 && x67 && x21 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( ~x70 && x65 && ~x66 && x67 && x21 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x67 && x21 && ~x8 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && x23 && x22 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && x23 && ~x22 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s805;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && ~x23 && x22 && x3 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s805;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && ~x23 && x22 && ~x3 && x6 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && ~x23 && x22 && ~x3 && x6 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && ~x23 && x22 && ~x3 && x6 && ~x18 && x19 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && ~x23 && x22 && ~x3 && x6 && ~x18 && x19 && ~x15 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && ~x23 && x22 && ~x3 && x6 && ~x18 && ~x19 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && ~x23 && x22 && ~x3 && ~x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s107;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && ~x23 && ~x22 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	y25 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x70 && ~x65 )
						begin
							y6 = 1'b1;	y21 = 1'b1;	y26 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s109;
				s110 : if( x21 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s806;
						end
					else if( ~x21 && x23 && x22 )
						nx_state = s1;
					else if( ~x21 && x23 && ~x22 && x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x21 && x23 && ~x22 && ~x16 && x20 && x19 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x21 && x23 && ~x22 && ~x16 && x20 && ~x19 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else if( ~x21 && x23 && ~x22 && ~x16 && ~x20 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x21 && ~x23 && x22 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x21 && ~x23 && ~x22 )
						nx_state = s1;
					else nx_state = s110;
				s111 : if( x21 && x18 && x19 && x15 && x17 )
						begin
							y15 = 1'b1;	y20 = 1'b1;	
							nx_state = s665;
						end
					else if( x21 && x18 && x19 && x15 && ~x17 )
						begin
							y16 = 1'b1;	y20 = 1'b1;	
							nx_state = s795;
						end
					else if( x21 && x18 && x19 && ~x15 && x16 && x17 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( x21 && x18 && x19 && ~x15 && x16 && ~x17 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s796;
						end
					else if( x21 && x18 && x19 && ~x15 && ~x16 && x17 && x10 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x21 && x18 && x19 && ~x15 && ~x16 && x17 && ~x10 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && x18 && x19 && ~x15 && ~x16 && x17 && ~x10 && x8 && ~x9 )
						nx_state = s1;
					else if( x21 && x18 && x19 && ~x15 && ~x16 && x17 && ~x10 && ~x8 )
						nx_state = s1;
					else if( x21 && x18 && x19 && ~x15 && ~x16 && ~x17 && x9 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x21 && x18 && x19 && ~x15 && ~x16 && ~x17 && ~x9 && x8 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && x18 && x19 && ~x15 && ~x16 && ~x17 && ~x9 && x8 && ~x10 )
						nx_state = s1;
					else if( x21 && x18 && x19 && ~x15 && ~x16 && ~x17 && ~x9 && ~x8 )
						nx_state = s1;
					else if( x21 && x18 && ~x19 && x16 && x15 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s476;
						end
					else if( x21 && x18 && ~x19 && x16 && ~x15 && x17 && x14 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s795;
						end
					else if( x21 && x18 && ~x19 && x16 && ~x15 && x17 && ~x14 )
						begin
							y12 = 1'b1;	y19 = 1'b1;	
							nx_state = s794;
						end
					else if( x21 && x18 && ~x19 && x16 && ~x15 && ~x17 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( x21 && x18 && ~x19 && ~x16 && x17 && x15 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( x21 && x18 && ~x19 && ~x16 && x17 && x15 && ~x3 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x21 && x18 && ~x19 && ~x16 && x17 && x15 && ~x3 && ~x5 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s793;
						end
					else if( x21 && x18 && ~x19 && ~x16 && x17 && ~x15 )
						begin
							y6 = 1'b1;	y19 = 1'b1;	
							nx_state = s682;
						end
					else if( x21 && x18 && ~x19 && ~x16 && ~x17 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( x21 && x18 && ~x19 && ~x16 && ~x17 && ~x3 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x21 && x18 && ~x19 && ~x16 && ~x17 && ~x3 && ~x5 && x15 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y28 = 1'b1;	
							nx_state = s807;
						end
					else if( x21 && x18 && ~x19 && ~x16 && ~x17 && ~x3 && ~x5 && ~x15 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( x21 && ~x18 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( x21 && ~x18 && ~x3 && x19 && x15 && x17 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x21 && ~x18 && ~x3 && x19 && x15 && x17 && ~x5 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s793;
						end
					else if( x21 && ~x18 && ~x3 && x19 && x15 && ~x17 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s808;
						end
					else if( x21 && ~x18 && ~x3 && x19 && x15 && ~x17 && ~x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && x16 && x17 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && x16 && x17 && ~x5 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y20 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s795;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && x16 && ~x17 && x14 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && x16 && ~x17 && x14 && ~x5 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y20 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s795;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && x16 && ~x17 && ~x14 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && x16 && ~x17 && ~x14 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && x16 && ~x17 && ~x14 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && x16 && ~x17 && ~x14 && ~x8 )
						nx_state = s1;
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && x17 && x12 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && x17 && x12 && ~x5 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y20 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s795;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && x17 && ~x12 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && x17 && ~x12 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && x17 && ~x12 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && x17 && ~x12 && ~x8 )
						nx_state = s1;
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && ~x17 && x13 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && ~x17 && x13 && ~x5 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y20 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s795;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && ~x17 && ~x13 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && ~x17 && ~x13 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && ~x17 && ~x13 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && ~x17 && ~x13 && ~x8 )
						nx_state = s1;
					else if( x21 && ~x18 && ~x3 && ~x19 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( x21 && ~x18 && ~x3 && ~x19 && ~x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x21 && x22 && x23 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x21 && x22 && ~x23 && x15 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x21 && x22 && ~x23 && ~x15 && x19 && x18 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x21 && x22 && ~x23 && ~x15 && x19 && ~x18 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x21 && x22 && ~x23 && ~x15 && ~x19 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x21 && ~x22 && x23 && x4 && x19 && x16 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x21 && ~x22 && x23 && x4 && x19 && ~x16 )
						begin
							y15 = 1'b1;	y20 = 1'b1;	
							nx_state = s665;
						end
					else if( ~x21 && ~x22 && x23 && x4 && ~x19 && x20 && x16 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s724;
						end
					else if( ~x21 && ~x22 && x23 && x4 && ~x19 && x20 && ~x16 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x21 && ~x22 && x23 && x4 && ~x19 && ~x20 )
						begin
							y3 = 1'b1;	y12 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s113;
						end
					else if( ~x21 && ~x22 && x23 && ~x4 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x21 && ~x22 && ~x23 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else nx_state = s111;
				s112 : if( x21 && x18 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && x18 && x15 && ~x17 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	
							nx_state = s807;
						end
					else if( x21 && x18 && ~x15 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x21 && ~x18 && x19 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && ~x18 && x19 && x15 && ~x17 )
						begin
							y8 = 1'b1;	
							nx_state = s568;
						end
					else if( x21 && ~x18 && x19 && ~x15 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s795;
						end
					else if( x21 && ~x18 && ~x19 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x21 && x22 && x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s301;
						end
					else nx_state = s112;
				s113 : if( x21 && x6 && x18 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && x6 && x18 && x15 && ~x17 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	
							nx_state = s807;
						end
					else if( x21 && x6 && x18 && ~x15 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x21 && x6 && ~x18 && x19 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && x6 && ~x18 && x19 && x15 && ~x17 )
						begin
							y8 = 1'b1;	
							nx_state = s568;
						end
					else if( x21 && x6 && ~x18 && x19 && ~x15 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s795;
						end
					else if( x21 && x6 && ~x18 && ~x19 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s110;
						end
					else if( x21 && ~x6 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s666;
						end
					else if( ~x21 && x23 && x22 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && x23 && x22 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && x23 && x22 && ~x18 && x19 && x15 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s666;
						end
					else if( ~x21 && x23 && x22 && ~x18 && x19 && ~x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( ~x21 && x23 && x22 && ~x18 && ~x19 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x21 && x23 && ~x22 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s301;
						end
					else if( ~x21 && ~x23 && x22 )
						nx_state = s1;
					else if( ~x21 && ~x23 && ~x22 )
						begin
							y12 = 1'b1;	y19 = 1'b1;	
							nx_state = s794;
						end
					else nx_state = s113;
				s114 : if( 1'b1 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else nx_state = s114;
				s115 : if( x21 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s805;
						end
					else if( ~x21 && x22 && x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && x22 && ~x23 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s795;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && ~x19 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( ~x21 && ~x22 && x23 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s301;
						end
					else nx_state = s115;
				s116 : if( x13 && x17 && x21 && x16 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s810;
						end
					else if( x13 && x17 && x21 && ~x16 && x18 && x15 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s810;
						end
					else if( x13 && x17 && x21 && ~x16 && x18 && ~x15 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else if( x13 && x17 && x21 && ~x16 && ~x18 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s810;
						end
					else if( x13 && x17 && ~x21 && x22 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s810;
						end
					else if( x13 && x17 && ~x21 && ~x22 && x15 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s810;
						end
					else if( x13 && x17 && ~x21 && ~x22 && ~x15 && x19 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s810;
						end
					else if( x13 && x17 && ~x21 && ~x22 && ~x15 && ~x19 && x20 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s810;
						end
					else if( x13 && x17 && ~x21 && ~x22 && ~x15 && ~x19 && ~x20 && x16 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s810;
						end
					else if( x13 && x17 && ~x21 && ~x22 && ~x15 && ~x19 && ~x20 && ~x16 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else if( x13 && ~x17 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s810;
						end
					else if( ~x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s810;
						end
					else nx_state = s116;
				s117 : if( x66 && x15 && x12 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x66 && x15 && x12 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s609;
						end
					else if( x66 && x15 && ~x12 && x7 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x66 && x15 && ~x12 && ~x7 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x66 && ~x15 && x16 && x7 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s811;
						end
					else if( x66 && ~x15 && x16 && x7 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x66 && ~x15 && x16 && ~x7 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s707;
						end
					else if( x66 && ~x15 && ~x16 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s812;
						end
					else if( x66 && ~x15 && ~x16 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x66 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else nx_state = s117;
				s118 : if( x65 )
						nx_state = s1;
					else if( ~x65 && x20 )
						nx_state = s1;
					else if( ~x65 && ~x20 && x21 && x15 && x8 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x65 && ~x20 && x21 && x15 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s556;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x16 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x65 && ~x20 && ~x21 )
						begin
							y3 = 1'b1;	y20 = 1'b1;	
							nx_state = s120;
						end
					else nx_state = s118;
				s119 : if( x20 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x20 && x21 && x15 && x8 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x20 && x21 && x15 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s556;
						end
					else if( ~x20 && x21 && ~x15 && x16 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s131;
						end
					else if( ~x20 && x21 && ~x15 && ~x16 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else nx_state = s119;
				s120 : if( x21 )
						nx_state = s1;
					else if( ~x21 && x15 && x8 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && x15 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s556;
						end
					else if( ~x21 && ~x15 && x16 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x21 && ~x15 && ~x16 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s76;
						end
					else nx_state = s120;
				s121 : if( x20 )
						nx_state = s1;
					else if( ~x20 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	
							nx_state = s813;
						end
					else nx_state = s121;
				s122 : if( x24 && x26 && x19 )
						nx_state = s122;
					else if( x24 && x26 && ~x19 )
						nx_state = s1;
					else if( x24 && ~x26 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( ~x24 && x25 && x26 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x26 && x15 && x6 && x10 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s368;
						end
					else if( ~x24 && x25 && ~x26 && x15 && x6 && x10 && ~x11 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( ~x24 && x25 && ~x26 && x15 && x6 && x10 && ~x11 && ~x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x24 && x25 && ~x26 && x15 && x6 && ~x10 )
						begin
							y8 = 1'b1;	y17 = 1'b1;	y23 = 1'b1;	
							nx_state = s303;
						end
					else if( ~x24 && x25 && ~x26 && x15 && ~x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && x10 && x8 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && x10 && ~x8 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && x10 && ~x8 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && x10 && ~x8 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && x10 && ~x8 && ~x19 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && ~x10 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && ~x10 && ~x7 && x11 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && ~x10 && ~x7 && ~x11 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && ~x10 && ~x7 && ~x11 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && ~x10 && ~x7 && ~x11 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && ~x10 && ~x7 && ~x11 && ~x19 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && ~x10 && x11 && x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && ~x10 && x11 && ~x9 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && ~x10 && x11 && ~x9 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && ~x10 && x11 && ~x9 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && ~x10 && x11 && ~x9 && ~x19 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && ~x10 && ~x11 && x8 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && ~x10 && ~x11 && x8 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && ~x10 && ~x11 && x8 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && ~x10 && ~x11 && x8 && ~x19 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && ~x10 && ~x11 && ~x8 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && ~x16 && x6 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && ~x16 && ~x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x24 && ~x25 && x26 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else nx_state = s122;
				s123 : if( x68 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x68 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x68 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x68 && x20 && ~x18 )
						nx_state = s1;
					else if( x68 && ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x68 && ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x68 && ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x68 && ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( x68 && ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( x68 && ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( x68 && ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x68 && ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else if( ~x68 && x24 && x26 )
						begin
							y17 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x68 && x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x68 && x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x68 && x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x68 && x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x68 && ~x24 && x25 && x26 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x68 && ~x24 && x25 && ~x26 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 )
						nx_state = s1;
					else if( ~x68 && ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x68 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x68 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x68 && ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else nx_state = s123;
				s124 : if( x70 && x62 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x62 && x63 )
						begin
							y3 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s814;
						end
					else if( x70 && ~x62 && ~x63 && x64 )
						begin
							y16 = 1'b1;	
							nx_state = s293;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s815;
						end
					else if( ~x70 && x66 && x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && x66 && x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && x66 && x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x66 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x21 && x22 && x23 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && x66 && ~x21 && x22 && ~x23 && x18 && x14 )
						nx_state = s47;
					else if( ~x70 && x66 && ~x21 && x22 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s47;
					else if( ~x70 && x66 && ~x21 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x21 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x21 && ~x22 && x23 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( ~x70 && x66 && ~x21 && ~x22 && ~x23 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s362;
						end
					else if( ~x70 && ~x66 && x24 && x26 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x70 && ~x66 && x24 && x26 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x70 && ~x66 && x24 && x26 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && ~x66 && x24 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x66 && x24 && ~x26 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x24 && x25 && x26 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x70 && ~x66 && ~x24 && x25 && x26 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x70 && ~x66 && ~x24 && x25 && x26 && x19 && ~x14 && ~x13 )
						nx_state = s124;
					else if( ~x70 && ~x66 && ~x24 && x25 && x26 && ~x19 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x24 && x25 && ~x26 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x70 && ~x66 && ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x70 && ~x66 && ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && ~x66 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && ~x66 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else nx_state = s124;
				s125 : if( x69 && x24 && x26 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x69 && x24 && x26 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x69 && x24 && x26 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && x24 && x26 && ~x18 )
						nx_state = s1;
					else if( x69 && x24 && ~x26 )
						nx_state = s1;
					else if( x69 && ~x24 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x24 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x24 && x25 && x19 && ~x14 && ~x13 && x26 )
						nx_state = s125;
					else if( x69 && ~x24 && x25 && x19 && ~x14 && ~x13 && ~x26 )
						nx_state = s1;
					else if( x69 && ~x24 && x25 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else if( ~x69 && x62 && x14 && x13 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s816;
						end
					else if( ~x69 && x62 && x14 && ~x13 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s817;
						end
					else if( ~x69 && x62 && ~x14 )
						begin
							y13 = 1'b1;	
							nx_state = s769;
						end
					else if( ~x69 && ~x62 && x28 && x57 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && ~x62 && x28 && ~x57 )
						nx_state = s125;
					else if( ~x69 && ~x62 && ~x28 && x27 && x8 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && ~x62 && ~x28 && x27 && ~x8 && x37 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && ~x62 && ~x28 && x27 && ~x8 && ~x37 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s818;
						end
					else if( ~x69 && ~x62 && ~x28 && ~x27 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s503;
						end
					else nx_state = s125;
				s126 : if( x65 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x65 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x65 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && x22 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x22 && x18 && x13 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x65 && ~x22 && x18 && x13 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x65 && ~x22 && x18 && ~x13 && x12 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x65 && ~x22 && x18 && ~x13 && x12 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x65 && ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && ~x22 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x26 && x24 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( ~x65 && x26 && ~x24 && x25 )
						nx_state = s1;
					else if( ~x65 && x26 && ~x24 && ~x25 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && x26 && ~x24 && ~x25 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && x26 && ~x24 && ~x25 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x26 && ~x24 && ~x25 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x26 && x24 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s819;
						end
					else if( ~x65 && ~x26 && ~x24 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x65 && ~x26 && ~x24 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x65 && ~x26 && ~x24 && x25 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x26 && ~x24 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x26 && ~x24 && ~x25 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x65 && ~x26 && ~x24 && ~x25 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x65 && ~x26 && ~x24 && ~x25 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x26 && ~x24 && ~x25 && ~x17 )
						nx_state = s1;
					else nx_state = s126;
				s127 : if( x70 && x62 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x70 && ~x62 && x12 && x15 && x13 && x3 )
						begin
							y3 = 1'b1;	y22 = 1'b1;	y23 = 1'b1;	
							nx_state = s671;
						end
					else if( x70 && ~x62 && x12 && x15 && x13 && ~x3 && x14 )
						begin
							y3 = 1'b1;	y22 = 1'b1;	y23 = 1'b1;	
							nx_state = s671;
						end
					else if( x70 && ~x62 && x12 && x15 && x13 && ~x3 && ~x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s230;
						end
					else if( x70 && ~x62 && x12 && x15 && ~x13 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( x70 && ~x62 && x12 && ~x15 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x70 && ~x62 && ~x12 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( ~x70 && x66 && x21 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x70 && x66 && ~x21 && x22 && x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s336;
						end
					else if( ~x70 && x66 && ~x21 && x22 && ~x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s107;
						end
					else if( ~x70 && x66 && ~x21 && ~x22 )
						begin
							y8 = 1'b1;	y18 = 1'b1;	
							nx_state = s152;
						end
					else if( ~x70 && ~x66 && x24 && x11 && x26 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x66 && x24 && x11 && ~x26 && x13 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && ~x66 && x24 && x11 && ~x26 && x13 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && ~x66 && x24 && x11 && ~x26 && x13 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && ~x66 && x24 && x11 && ~x26 && x13 && ~x20 )
						nx_state = s1;
					else if( ~x70 && ~x66 && x24 && x11 && ~x26 && ~x13 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s497;
						end
					else if( ~x70 && ~x66 && x24 && ~x11 && x26 && x12 && x13 && x16 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x70 && ~x66 && x24 && ~x11 && x26 && x12 && x13 && x16 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x70 && ~x66 && x24 && ~x11 && x26 && x12 && x13 && x16 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && ~x66 && x24 && ~x11 && x26 && x12 && x13 && x16 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x66 && x24 && ~x11 && x26 && x12 && x13 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x66 && x24 && ~x11 && x26 && x12 && ~x13 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x66 && x24 && ~x11 && x26 && ~x12 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x66 && x24 && ~x11 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && ~x66 && x24 && ~x11 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && ~x66 && x24 && ~x11 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && ~x66 && x24 && ~x11 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x24 && x25 && x26 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x66 && ~x24 && x25 && ~x26 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x70 && ~x66 && ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x70 && ~x66 && ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x66 && ~x24 && ~x25 && ~x26 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else nx_state = s127;
				s128 : if( x70 && x63 && x18 && x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s820;
						end
					else if( x70 && x63 && x18 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s821;
						end
					else if( x70 && x63 && x18 && ~x5 && ~x6 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( x70 && x63 && ~x18 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x70 && x63 && ~x18 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x70 && x63 && ~x18 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x70 && x63 && ~x18 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && x65 && x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x70 && ~x63 && x64 && x65 && x10 && ~x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x70 && ~x63 && x64 && x65 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && x65 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && ~x65 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x63 && x64 && ~x65 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x63 && x64 && ~x65 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && ~x65 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x21 && x22 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( x70 && ~x63 && ~x64 && x21 && ~x22 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( x70 && ~x63 && ~x64 && x21 && ~x22 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && ~x21 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( x70 && ~x63 && ~x64 && ~x21 && ~x23 )
						nx_state = s1;
					else if( ~x70 && x65 && x21 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && x22 && x23 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && x22 && ~x23 && x15 && x9 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( ~x70 && x65 && ~x21 && x22 && ~x23 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && x65 && ~x21 && x22 && ~x23 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && x22 && ~x23 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s495;
						end
					else if( ~x70 && x65 && ~x21 && ~x22 && x23 && x17 && x15 && x9 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && x65 && ~x21 && ~x22 && x23 && x17 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && x65 && ~x21 && ~x22 && x23 && x17 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && ~x22 && x23 && x17 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s495;
						end
					else if( ~x70 && x65 && ~x21 && ~x22 && x23 && ~x17 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x70 && x65 && ~x21 && ~x22 && ~x23 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x70 && ~x65 && x66 && x63 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && ~x63 && x62 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && ~x63 && ~x62 )
						begin
							y21 = 1'b1;	
							nx_state = s822;
						end
					else if( ~x70 && ~x65 && ~x66 && x25 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x25 )
						nx_state = s1;
					else nx_state = s128;
				s129 : if( x21 )
						nx_state = s1;
					else if( ~x21 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else nx_state = s129;
				s130 : if( x70 && x62 && x20 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x70 && x62 && x20 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x70 && x62 && x20 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( x70 && x62 && x20 && ~x21 )
						nx_state = s1;
					else if( x70 && x62 && ~x20 )
						begin
							y5 = 1'b1;	
							nx_state = s791;
						end
					else if( x70 && ~x62 && x63 && x65 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x70 && ~x62 && x63 && x65 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x70 && ~x62 && x63 && x65 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( x70 && ~x62 && x63 && x65 && ~x22 )
						nx_state = s1;
					else if( x70 && ~x62 && x63 && ~x65 && x67 )
						begin
							y22 = 1'b1;	
							nx_state = s823;
						end
					else if( x70 && ~x62 && x63 && ~x65 && ~x67 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x70 && ~x62 && x63 && ~x65 && ~x67 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x70 && ~x62 && x63 && ~x65 && ~x67 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && x63 && ~x65 && ~x67 && ~x14 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && x66 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x66 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x66 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && x66 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x14 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && x66 && x21 && x22 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x66 && x21 && ~x22 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x66 && x21 && ~x22 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && x66 && ~x21 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x66 && ~x21 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x66 && x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x66 && x26 && ~x25 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x66 && x26 && ~x25 && ~x24 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x66 && ~x26 )
						nx_state = s1;
					else if( ~x70 && x68 && x21 && x20 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( ~x70 && x68 && x21 && ~x20 )
						nx_state = s1;
					else if( ~x70 && x68 && ~x21 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s131;
						end
					else if( ~x70 && ~x68 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else nx_state = s130;
				s131 : if( x70 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s824;
						end
					else if( ~x70 && x65 && x21 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s132;
						end
					else if( ~x70 && ~x65 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x20 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x70 && ~x65 && ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x70 && ~x65 && ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x70 && ~x65 && ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x70 && ~x65 && ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else nx_state = s131;
				s132 : if( x70 && x2 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( x70 && ~x2 )
						nx_state = s132;
					else if( ~x70 && x21 && x20 && x2 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s825;
						end
					else if( ~x70 && x21 && x20 && ~x2 && x18 && x15 && x10 && x11 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s600;
						end
					else if( ~x70 && x21 && x20 && ~x2 && x18 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s601;
						end
					else if( ~x70 && x21 && x20 && ~x2 && x18 && x15 && x10 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s776;
						end
					else if( ~x70 && x21 && x20 && ~x2 && x18 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( ~x70 && x21 && x20 && ~x2 && x18 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s602;
						end
					else if( ~x70 && x21 && x20 && ~x2 && x18 && ~x15 && x16 && x10 && x12 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( ~x70 && x21 && x20 && ~x2 && x18 && ~x15 && x16 && x10 && ~x12 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && x21 && x20 && ~x2 && x18 && ~x15 && x16 && ~x10 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( ~x70 && x21 && x20 && ~x2 && x18 && ~x15 && ~x16 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && x21 && x20 && ~x2 && ~x18 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	
							nx_state = s826;
						end
					else if( ~x70 && x21 && ~x20 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	
							nx_state = s826;
						end
					else if( ~x70 && ~x21 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	
							nx_state = s826;
						end
					else nx_state = s132;
				s133 : if( x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( ~x21 )
						nx_state = s1;
					else nx_state = s133;
				s134 : if( x69 && x65 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x69 && ~x65 && x66 && x21 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s18;
						end
					else if( x69 && ~x65 && x66 && ~x21 && x22 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s565;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && x10 && x16 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && x10 && ~x16 && x17 && x15 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && x10 && ~x16 && x17 && ~x15 && x3 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s181;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && x10 && ~x16 && x17 && ~x15 && ~x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s827;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && x10 && ~x16 && ~x17 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && ~x10 && x16 && x15 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s828;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && ~x10 && x16 && ~x15 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s267;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && ~x10 && ~x16 && x17 && x15 && x14 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	
							nx_state = s220;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && ~x10 && ~x16 && x17 && x15 && ~x14 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s149;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && ~x10 && ~x16 && x17 && ~x15 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s149;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && ~x10 && ~x16 && ~x17 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s829;
						end
					else if( x69 && ~x65 && ~x66 && x68 && x21 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && ~x65 && ~x66 && x68 && ~x21 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x65 && ~x66 && ~x68 && x22 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x65 && ~x66 && ~x68 && ~x22 && x21 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x65 && ~x66 && ~x68 && ~x22 && ~x21 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x69 && x45 && x12 && x46 && x14 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && x45 && x12 && x46 && ~x14 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x69 && x45 && x12 && ~x46 && x2 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x69 && x45 && x12 && ~x46 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && x45 && ~x12 && x46 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && x45 && ~x12 && ~x46 && x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && x45 && ~x12 && ~x46 && ~x2 )
						nx_state = s134;
					else if( ~x69 && ~x45 && x46 && x47 && x2 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x45 && x46 && x47 && x2 && ~x8 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x69 && ~x45 && x46 && x47 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x45 && x46 && ~x47 && x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x45 && x46 && ~x47 && ~x2 )
						nx_state = s134;
					else if( ~x69 && ~x45 && ~x46 && x2 && x12 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x45 && ~x46 && x2 && ~x12 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x69 && ~x45 && ~x46 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else nx_state = s134;
				s135 : if( x61 && x60 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x61 && ~x60 && x62 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x61 && ~x60 && ~x62 )
						nx_state = s47;
					else if( ~x61 && x60 )
						nx_state = s47;
					else if( ~x61 && ~x60 && x62 )
						nx_state = s47;
					else if( ~x61 && ~x60 && ~x62 )
						nx_state = s1;
					else nx_state = s135;
				s136 : if( x60 && x61 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else if( x60 && ~x61 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( ~x60 && x62 && x61 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x60 && x62 && x61 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x60 && x62 && x61 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( ~x60 && x62 && x61 && ~x18 )
						nx_state = s1;
					else if( ~x60 && x62 && ~x61 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s830;
						end
					else if( ~x60 && ~x62 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else nx_state = s136;
				s137 : if( x70 && x62 && x12 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && x62 && ~x12 )
						nx_state = s137;
					else if( x70 && ~x62 && x63 && x15 && x14 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x70 && ~x62 && x63 && x15 && ~x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s230;
						end
					else if( x70 && ~x62 && x63 && ~x15 && x12 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && ~x62 && x63 && ~x15 && ~x12 )
						nx_state = s137;
					else if( x70 && ~x62 && ~x63 && x30 && x31 )
						begin
							y33 = 1'b1;	
							nx_state = s589;
						end
					else if( x70 && ~x62 && ~x63 && x30 && ~x31 )
						begin
							y47 = 1'b1;	y49 = 1'b1;	y58 = 1'b1;	
							y61 = 1'b1;	y68 = 1'b1;	
							nx_state = s831;
						end
					else if( x70 && ~x62 && ~x63 && ~x30 )
						begin
							y47 = 1'b1;	y52 = 1'b1;	y61 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s353;
						end
					else if( ~x70 && x65 && x66 && x61 && x60 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && x65 && x66 && x61 && ~x60 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s487;
						end
					else if( ~x70 && x65 && x66 && ~x61 && x60 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s487;
						end
					else if( ~x70 && x65 && x66 && ~x61 && ~x60 )
						nx_state = s47;
					else if( ~x70 && x65 && ~x66 )
						begin
							y15 = 1'b1;	y21 = 1'b1;	y28 = 1'b1;	
							nx_state = s832;
						end
					else if( ~x70 && ~x65 && x66 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && ~x65 && ~x66 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x70 && ~x65 && ~x66 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x70 && ~x65 && ~x66 && x19 && ~x14 && ~x13 )
						nx_state = s137;
					else if( ~x70 && ~x65 && ~x66 && ~x19 )
						nx_state = s1;
					else nx_state = s137;
				s138 : if( x69 && x65 && x60 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s139;
						end
					else if( x69 && x65 && ~x60 && x61 )
						nx_state = s1;
					else if( x69 && x65 && ~x60 && ~x61 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s559;
						end
					else if( x69 && ~x65 && x21 && x3 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	
							nx_state = s758;
						end
					else if( x69 && ~x65 && x21 && ~x3 && x20 && x16 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s233;
						end
					else if( x69 && ~x65 && x21 && ~x3 && x20 && x16 && ~x10 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x65 && x21 && ~x3 && x20 && ~x16 && x17 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x65 && x21 && ~x3 && x20 && ~x16 && ~x17 )
						begin
							y5 = 1'b1;	y17 = 1'b1;	
							nx_state = s721;
						end
					else if( x69 && ~x65 && x21 && ~x3 && ~x20 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( x69 && ~x65 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( x69 && ~x65 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( x69 && ~x65 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x21 && ~x20 )
						nx_state = s1;
					else if( ~x69 && x63 && x55 && x17 && x41 && x19 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x69 && x63 && x55 && x17 && x41 && ~x19 )
						nx_state = s138;
					else if( ~x69 && x63 && x55 && x17 && ~x41 && x19 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x69 && x63 && x55 && x17 && ~x41 && ~x19 )
						nx_state = s138;
					else if( ~x69 && x63 && x55 && ~x17 && x20 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && x63 && x55 && ~x17 && ~x20 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( ~x69 && x63 && x55 && ~x17 && ~x20 && ~x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s503;
						end
					else if( ~x69 && x63 && ~x55 && x10 && x11 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && x63 && ~x55 && x10 && ~x11 && x43 && x4 && x32 )
						nx_state = s138;
					else if( ~x69 && x63 && ~x55 && x10 && ~x11 && x43 && x4 && ~x32 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x69 && x63 && ~x55 && x10 && ~x11 && x43 && ~x4 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( ~x69 && x63 && ~x55 && x10 && ~x11 && ~x43 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && x63 && ~x55 && ~x10 && x42 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y27 = 1'b1;	
							nx_state = s833;
						end
					else if( ~x69 && x63 && ~x55 && ~x10 && ~x42 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && ~x63 && x64 && x40 && x17 && x19 && x10 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x69 && ~x63 && x64 && x40 && x17 && x19 && ~x10 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x69 && ~x63 && x64 && x40 && x17 && ~x19 )
						nx_state = s138;
					else if( ~x69 && ~x63 && x64 && x40 && ~x17 && x20 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && ~x63 && x64 && x40 && ~x17 && ~x20 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && ~x63 && x64 && x40 && ~x17 && ~x20 && ~x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x69 && ~x63 && x64 && ~x40 && x11 && x10 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && ~x63 && x64 && ~x40 && x11 && ~x10 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s638;
						end
					else if( ~x69 && ~x63 && x64 && ~x40 && ~x11 && x10 && x12 && x4 && x1 )
						nx_state = s138;
					else if( ~x69 && ~x63 && x64 && ~x40 && ~x11 && x10 && x12 && x4 && ~x1 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x69 && ~x63 && x64 && ~x40 && ~x11 && x10 && x12 && ~x4 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && ~x63 && x64 && ~x40 && ~x11 && x10 && ~x12 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && ~x63 && x64 && ~x40 && ~x11 && ~x10 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && ~x63 && ~x64 && x44 && x17 && x19 && x10 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x69 && ~x63 && ~x64 && x44 && x17 && x19 && ~x10 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s631;
						end
					else if( ~x69 && ~x63 && ~x64 && x44 && x17 && ~x19 )
						nx_state = s138;
					else if( ~x69 && ~x63 && ~x64 && x44 && ~x17 && x20 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s513;
						end
					else if( ~x69 && ~x63 && ~x64 && x44 && ~x17 && ~x20 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && ~x63 && ~x64 && x44 && ~x17 && ~x20 && ~x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x69 && ~x63 && ~x64 && ~x44 && x11 && x10 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x69 && ~x63 && ~x64 && ~x44 && x11 && ~x10 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s638;
						end
					else if( ~x69 && ~x63 && ~x64 && ~x44 && ~x11 && x10 && x12 && x4 && x1 )
						nx_state = s138;
					else if( ~x69 && ~x63 && ~x64 && ~x44 && ~x11 && x10 && x12 && x4 && ~x1 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s631;
						end
					else if( ~x69 && ~x63 && ~x64 && ~x44 && ~x11 && x10 && x12 && ~x4 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && ~x63 && ~x64 && ~x44 && ~x11 && x10 && ~x12 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else if( ~x69 && ~x63 && ~x64 && ~x44 && ~x11 && ~x10 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else nx_state = s138;
				s139 : if( x60 && x61 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x60 && x61 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x60 && x61 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x60 && x61 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x60 && ~x61 && x15 && x5 && x12 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s834;
						end
					else if( x60 && ~x61 && x15 && x5 && x12 && ~x7 )
						begin
							y4 = 1'b1;	
							nx_state = s834;
						end
					else if( x60 && ~x61 && x15 && x5 && ~x12 && x7 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( x60 && ~x61 && x15 && x5 && ~x12 && ~x7 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s242;
						end
					else if( x60 && ~x61 && x15 && ~x5 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( x60 && ~x61 && ~x15 && x16 && x7 && x12 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( x60 && ~x61 && ~x15 && x16 && x7 && x12 && ~x5 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( x60 && ~x61 && ~x15 && x16 && x7 && ~x12 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( x60 && ~x61 && ~x15 && x16 && ~x7 && x12 && x9 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( x60 && ~x61 && ~x15 && x16 && ~x7 && x12 && ~x9 && x11 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( x60 && ~x61 && ~x15 && x16 && ~x7 && x12 && ~x9 && ~x11 )
						nx_state = s1;
					else if( x60 && ~x61 && ~x15 && x16 && ~x7 && ~x12 && x11 && x10 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( x60 && ~x61 && ~x15 && x16 && ~x7 && ~x12 && x11 && ~x10 )
						nx_state = s1;
					else if( x60 && ~x61 && ~x15 && x16 && ~x7 && ~x12 && ~x11 && x8 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( x60 && ~x61 && ~x15 && x16 && ~x7 && ~x12 && ~x11 && ~x8 )
						nx_state = s1;
					else if( x60 && ~x61 && ~x15 && ~x16 && x5 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s812;
						end
					else if( x60 && ~x61 && ~x15 && ~x16 && x5 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x60 && ~x61 && ~x15 && ~x16 && ~x5 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x60 && x61 && x62 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else if( ~x60 && x61 && ~x62 && x15 && x5 && x12 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s834;
						end
					else if( ~x60 && x61 && ~x62 && x15 && x5 && x12 && ~x7 )
						begin
							y4 = 1'b1;	
							nx_state = s834;
						end
					else if( ~x60 && x61 && ~x62 && x15 && x5 && ~x12 && x7 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x60 && x61 && ~x62 && x15 && x5 && ~x12 && ~x7 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x60 && x61 && ~x62 && x15 && ~x5 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x60 && x61 && ~x62 && ~x15 && x16 && x7 && x12 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x60 && x61 && ~x62 && ~x15 && x16 && x7 && x12 && ~x5 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x60 && x61 && ~x62 && ~x15 && x16 && x7 && ~x12 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x60 && x61 && ~x62 && ~x15 && x16 && ~x7 && x12 && x9 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x60 && x61 && ~x62 && ~x15 && x16 && ~x7 && x12 && ~x9 && x11 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x60 && x61 && ~x62 && ~x15 && x16 && ~x7 && x12 && ~x9 && ~x11 )
						nx_state = s1;
					else if( ~x60 && x61 && ~x62 && ~x15 && x16 && ~x7 && ~x12 && x11 && x10 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x60 && x61 && ~x62 && ~x15 && x16 && ~x7 && ~x12 && x11 && ~x10 )
						nx_state = s1;
					else if( ~x60 && x61 && ~x62 && ~x15 && x16 && ~x7 && ~x12 && ~x11 && x8 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x60 && x61 && ~x62 && ~x15 && x16 && ~x7 && ~x12 && ~x11 && ~x8 )
						nx_state = s1;
					else if( ~x60 && x61 && ~x62 && ~x15 && ~x16 && x5 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s812;
						end
					else if( ~x60 && x61 && ~x62 && ~x15 && ~x16 && x5 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x60 && x61 && ~x62 && ~x15 && ~x16 && ~x5 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x60 && ~x61 && x62 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x60 && ~x61 && ~x62 )
						begin
							y3 = 1'b1;	
							nx_state = s835;
						end
					else nx_state = s139;
				s140 : if( x70 && x62 && x1 && x2 && x3 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x70 && x62 && x1 && x2 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x70 && x62 && x1 && ~x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x70 && x62 && ~x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x70 && ~x62 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s836;
						end
					else if( ~x70 && x65 && x60 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s139;
						end
					else if( ~x70 && x65 && ~x60 && x61 )
						begin
							y2 = 1'b1;	y19 = 1'b1;	y24 = 1'b1;	
							nx_state = s837;
						end
					else if( ~x70 && x65 && ~x60 && ~x61 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && ~x65 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else nx_state = s140;
				s141 : if( x60 )
						nx_state = s331;
					else if( ~x60 && x61 )
						nx_state = s331;
					else if( ~x60 && ~x61 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else nx_state = s141;
				s142 : if( x60 )
						nx_state = s331;
					else if( ~x60 && x61 )
						nx_state = s331;
					else if( ~x60 && ~x61 && x17 && x62 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x60 && ~x61 && x17 && ~x62 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x60 && ~x61 && ~x17 )
						nx_state = s118;
					else nx_state = s142;
				s143 : if( x60 && x15 && x12 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x60 && x15 && x12 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s609;
						end
					else if( x60 && x15 && ~x12 && x7 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x60 && x15 && ~x12 && ~x7 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s565;
						end
					else if( x60 && ~x15 && x16 && x7 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s811;
						end
					else if( x60 && ~x15 && x16 && x7 && ~x12 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x60 && ~x15 && x16 && ~x7 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x60 && ~x15 && ~x16 && x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s764;
						end
					else if( x60 && ~x15 && ~x16 && ~x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x60 && x61 && x15 && x12 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( ~x60 && x61 && x15 && x12 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s609;
						end
					else if( ~x60 && x61 && x15 && ~x12 && x7 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x60 && x61 && x15 && ~x12 && ~x7 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s565;
						end
					else if( ~x60 && x61 && ~x15 && x16 && x7 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s811;
						end
					else if( ~x60 && x61 && ~x15 && x16 && x7 && ~x12 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x60 && x61 && ~x15 && x16 && ~x7 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x60 && x61 && ~x15 && ~x16 && x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s764;
						end
					else if( ~x60 && x61 && ~x15 && ~x16 && ~x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x60 && ~x61 && x62 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y24 = 1'b1;	
							nx_state = s136;
						end
					else if( ~x60 && ~x61 && ~x62 )
						begin
							y25 = 1'b1;	
							nx_state = s838;
						end
					else nx_state = s143;
				s144 : if( x69 && x70 && x65 )
						nx_state = s1;
					else if( x69 && x70 && ~x65 && x17 && x18 && x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	
							nx_state = s20;
						end
					else if( x69 && x70 && ~x65 && x17 && x18 && ~x1 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && x70 && ~x65 && x17 && x18 && ~x1 && ~x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x70 && ~x65 && x17 && ~x18 && x6 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s320;
						end
					else if( x69 && x70 && ~x65 && x17 && ~x18 && ~x6 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s280;
						end
					else if( x69 && x70 && ~x65 && ~x17 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && ~x70 && x61 && x60 && x7 && x15 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x69 && ~x70 && x61 && x60 && x7 && ~x15 && x16 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s811;
						end
					else if( x69 && ~x70 && x61 && x60 && x7 && ~x15 && x16 && ~x12 && x3 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s487;
						end
					else if( x69 && ~x70 && x61 && x60 && x7 && ~x15 && x16 && ~x12 && ~x3 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x69 && ~x70 && x61 && x60 && x7 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s812;
						end
					else if( x69 && ~x70 && x61 && x60 && ~x7 && x15 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s609;
						end
					else if( x69 && ~x70 && x61 && x60 && ~x7 && x15 && ~x12 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && ~x70 && x61 && x60 && ~x7 && ~x15 && x16 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && x61 && x60 && ~x7 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && ~x70 && x61 && ~x60 && x62 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x69 && ~x70 && x61 && ~x60 && ~x62 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x69 && ~x70 && ~x61 && x60 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && x62 && x16 && x15 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && x62 && x16 && ~x15 && x11 && x12 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && x62 && x16 && ~x15 && x11 && ~x12 && x7 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && x62 && x16 && ~x15 && x11 && ~x12 && ~x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && x62 && x16 && ~x15 && ~x11 && x7 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && x62 && x16 && ~x15 && ~x11 && ~x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && x62 && ~x16 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && x15 && x16 && x9 && x11 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && x15 && x16 && x9 && ~x11 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && x15 && x16 && x9 && ~x11 && ~x7 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s564;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && x15 && x16 && ~x9 && x11 && x7 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s565;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && x15 && x16 && ~x9 && x11 && ~x7 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s251;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && x15 && x16 && ~x9 && ~x11 && x7 && x14 )
						nx_state = s331;
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && x15 && x16 && ~x9 && ~x11 && x7 && ~x14 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && x15 && x16 && ~x9 && ~x11 && ~x7 && x13 )
						nx_state = s331;
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && x15 && x16 && ~x9 && ~x11 && ~x7 && ~x13 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && x15 && ~x16 && x9 && x3 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && x15 && ~x16 && x9 && ~x3 && x7 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s738;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && x15 && ~x16 && x9 && ~x3 && ~x7 && x11 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s738;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && x15 && ~x16 && x9 && ~x3 && ~x7 && ~x11 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && x15 && ~x16 && ~x9 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && x15 && ~x16 && ~x9 && ~x3 && x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && x15 && ~x16 && ~x9 && ~x3 && ~x5 && x7 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s839;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && x15 && ~x16 && ~x9 && ~x3 && ~x5 && ~x7 && x11 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && x15 && ~x16 && ~x9 && ~x3 && ~x5 && ~x7 && ~x11 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && ~x15 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && x11 && x9 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && x11 && ~x9 && x7 && x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && x11 && ~x9 && x7 && ~x5 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s839;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && x11 && ~x9 && ~x7 && x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s553;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && x11 && ~x9 && ~x7 && ~x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && x7 && x9 && x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s554;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && x7 && x9 && ~x5 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s707;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && x7 && ~x9 && x8 && x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s554;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && x7 && ~x9 && x8 && ~x5 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s707;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && x7 && ~x9 && ~x8 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && ~x7 && x9 && x10 && x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s554;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && ~x7 && x9 && x10 && ~x5 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s707;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && ~x7 && x9 && ~x10 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && ~x7 && ~x9 && x12 && x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s554;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && ~x7 && ~x9 && x12 && ~x5 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s707;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && ~x7 && ~x9 && ~x12 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && ~x16 && x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x69 && ~x70 && ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && ~x16 && ~x5 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s139;
						end
					else if( ~x69 && x64 && x61 && x35 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( ~x69 && x64 && x61 && ~x35 && x13 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x69 && x64 && x61 && ~x35 && ~x13 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s593;
						end
					else if( ~x69 && x64 && ~x61 && x10 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x64 && ~x61 && ~x10 && x11 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x69 && x64 && ~x61 && ~x10 && ~x11 && x7 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( ~x69 && x64 && ~x61 && ~x10 && ~x11 && ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && ~x64 && x14 && x35 )
						nx_state = s1;
					else if( ~x69 && ~x64 && x14 && ~x35 && x13 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x69 && ~x64 && x14 && ~x35 && ~x13 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s593;
						end
					else if( ~x69 && ~x64 && ~x14 && x10 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && ~x64 && ~x14 && ~x10 && x11 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x69 && ~x64 && ~x14 && ~x10 && ~x11 && x7 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( ~x69 && ~x64 && ~x14 && ~x10 && ~x11 && ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else nx_state = s144;
				s145 : if( x69 && x65 && x60 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x69 && x65 && ~x60 && x61 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x69 && x65 && ~x60 && ~x61 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && ~x65 && x21 && x16 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s233;
						end
					else if( x69 && ~x65 && x21 && x16 && ~x10 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x65 && x21 && ~x16 && x17 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x65 && x21 && ~x16 && ~x17 )
						begin
							y5 = 1'b1;	y17 = 1'b1;	
							nx_state = s721;
						end
					else if( x69 && ~x65 && ~x21 && x3 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( x69 && ~x65 && ~x21 && ~x3 && x19 && x16 && x10 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( x69 && ~x65 && ~x21 && ~x3 && x19 && x16 && ~x10 )
						begin
							y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s233;
						end
					else if( x69 && ~x65 && ~x21 && ~x3 && x19 && ~x16 && x17 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x65 && ~x21 && ~x3 && x19 && ~x16 && ~x17 )
						begin
							y5 = 1'b1;	y17 = 1'b1;	
							nx_state = s721;
						end
					else if( x69 && ~x65 && ~x21 && ~x3 && ~x19 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	
							nx_state = s758;
						end
					else if( ~x69 && x70 && x61 && x7 && x35 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && x70 && x61 && x7 && x35 && ~x1 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s840;
						end
					else if( ~x69 && x70 && x61 && x7 && ~x35 && x1 )
						nx_state = s145;
					else if( ~x69 && x70 && x61 && x7 && ~x35 && ~x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x69 && x70 && x61 && ~x7 )
						nx_state = s145;
					else if( ~x69 && x70 && ~x61 && x3 )
						begin
							y10 = 1'b1;	
							nx_state = s841;
						end
					else if( ~x69 && x70 && ~x61 && ~x3 && x2 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s842;
						end
					else if( ~x69 && x70 && ~x61 && ~x3 && ~x2 && x28 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x69 && x70 && ~x61 && ~x3 && ~x2 && ~x28 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( ~x69 && ~x70 && x10 && x5 && x44 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( ~x69 && ~x70 && x10 && x5 && x44 && ~x3 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x69 && ~x70 && x10 && x5 && x44 && ~x3 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x69 && ~x70 && x10 && x5 && ~x44 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && x10 && ~x5 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && ~x10 && x44 && x11 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && ~x70 && ~x10 && x44 && x11 && ~x1 && x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && ~x70 && ~x10 && x44 && x11 && ~x1 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && ~x10 && x44 && ~x11 )
						nx_state = s145;
					else if( ~x69 && ~x70 && ~x10 && ~x44 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && ~x70 && ~x10 && ~x44 && ~x1 && x3 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( ~x69 && ~x70 && ~x10 && ~x44 && ~x1 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else nx_state = s145;
				s146 : if( x70 && x62 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x70 && ~x62 && x5 )
						begin
							y8 = 1'b1;	
							nx_state = s744;
						end
					else if( x70 && ~x62 && ~x5 && x21 && x22 && x10 && x14 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( x70 && ~x62 && ~x5 && x21 && x22 && x10 && ~x14 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x70 && ~x62 && ~x5 && x21 && x22 && ~x10 && x11 && x14 && x8 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( x70 && ~x62 && ~x5 && x21 && x22 && ~x10 && x11 && x14 && ~x8 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x5 && x21 && x22 && ~x10 && x11 && x14 && ~x8 && x6 && ~x7 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x5 && x21 && x22 && ~x10 && x11 && x14 && ~x8 && ~x6 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x5 && x21 && x22 && ~x10 && x11 && ~x14 && x7 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( x70 && ~x62 && ~x5 && x21 && x22 && ~x10 && x11 && ~x14 && ~x7 && x6 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x5 && x21 && x22 && ~x10 && x11 && ~x14 && ~x7 && x6 && ~x8 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x5 && x21 && x22 && ~x10 && x11 && ~x14 && ~x7 && ~x6 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x5 && x21 && x22 && ~x10 && ~x11 && x14 )
						begin
							y60 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y67 = 1'b1;	y68 = 1'b1;	
							nx_state = s516;
						end
					else if( x70 && ~x62 && ~x5 && x21 && x22 && ~x10 && ~x11 && ~x14 )
						begin
							y58 = 1'b1;	y59 = 1'b1;	y60 = 1'b1;	
							y62 = 1'b1;	
							nx_state = s516;
						end
					else if( x70 && ~x62 && ~x5 && x21 && ~x22 && x9 )
						begin
							y9 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y94 = 1'b1;	
							nx_state = s844;
						end
					else if( x70 && ~x62 && ~x5 && x21 && ~x22 && ~x9 && x11 && x14 && x10 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x70 && ~x62 && ~x5 && x21 && ~x22 && ~x9 && x11 && x14 && ~x10 )
						begin
							y62 = 1'b1;	y65 = 1'b1;	y90 = 1'b1;	
							y95 = 1'b1;	
							nx_state = s516;
						end
					else if( x70 && ~x62 && ~x5 && x21 && ~x22 && ~x9 && x11 && ~x14 && x10 )
						begin
							y38 = 1'b1;	
							nx_state = s845;
						end
					else if( x70 && ~x62 && ~x5 && x21 && ~x22 && ~x9 && x11 && ~x14 && ~x10 )
						begin
							y62 = 1'b1;	y65 = 1'b1;	y93 = 1'b1;	
							y94 = 1'b1;	
							nx_state = s516;
						end
					else if( x70 && ~x62 && ~x5 && x21 && ~x22 && ~x9 && ~x11 && x14 && x10 )
						begin
							y100 = 1'b1;	
							nx_state = s516;
						end
					else if( x70 && ~x62 && ~x5 && x21 && ~x22 && ~x9 && ~x11 && x14 && ~x10 )
						begin
							y46 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y73 = 1'b1;	y95 = 1'b1;	
							nx_state = s846;
						end
					else if( x70 && ~x62 && ~x5 && x21 && ~x22 && ~x9 && ~x11 && ~x14 && x10 )
						begin
							y62 = 1'b1;	y65 = 1'b1;	y78 = 1'b1;	
							y90 = 1'b1;	
							nx_state = s516;
						end
					else if( x70 && ~x62 && ~x5 && x21 && ~x22 && ~x9 && ~x11 && ~x14 && ~x10 )
						begin
							y74 = 1'b1;	
							nx_state = s847;
						end
					else if( x70 && ~x62 && ~x5 && ~x21 && x22 )
						begin
							y9 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y94 = 1'b1;	
							nx_state = s844;
						end
					else if( x70 && ~x62 && ~x5 && ~x21 && ~x22 && x10 && x11 && x9 )
						begin
							y9 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y90 = 1'b1;	
							nx_state = s848;
						end
					else if( x70 && ~x62 && ~x5 && ~x21 && ~x22 && x10 && x11 && ~x9 )
						begin
							y65 = 1'b1;	y90 = 1'b1;	y92 = 1'b1;	
							y93 = 1'b1;	
							nx_state = s516;
						end
					else if( x70 && ~x62 && ~x5 && ~x21 && ~x22 && x10 && ~x11 && x9 )
						begin
							y9 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y94 = 1'b1;	
							nx_state = s844;
						end
					else if( x70 && ~x62 && ~x5 && ~x21 && ~x22 && x10 && ~x11 && ~x9 )
						begin
							y65 = 1'b1;	y92 = 1'b1;	y94 = 1'b1;	
							y95 = 1'b1;	
							nx_state = s516;
						end
					else if( x70 && ~x62 && ~x5 && ~x21 && ~x22 && ~x10 && x9 )
						begin
							y9 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y94 = 1'b1;	
							nx_state = s849;
						end
					else if( x70 && ~x62 && ~x5 && ~x21 && ~x22 && ~x10 && ~x9 )
						begin
							y65 = 1'b1;	y90 = 1'b1;	y91 = 1'b1;	
							y92 = 1'b1;	y93 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x70 && x65 && x61 && x60 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x65 && x61 && x60 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x65 && x61 && x60 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( ~x70 && x65 && x61 && x60 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( ~x70 && x65 && x61 && ~x60 && x62 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && x16 && x7 && x12 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && x16 && x7 && ~x12 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && x16 && ~x7 && x12 && x14 && x11 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s251;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && x16 && ~x7 && x12 && x14 && ~x11 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && x16 && ~x7 && x12 && ~x14 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && x16 && ~x7 && x12 && ~x14 && x18 && ~x13 )
						nx_state = s118;
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && x16 && ~x7 && x12 && ~x14 && ~x18 )
						nx_state = s118;
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && x16 && ~x7 && ~x12 && x13 && x11 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s564;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && x16 && ~x7 && ~x12 && x13 && ~x11 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && x16 && ~x7 && ~x12 && ~x13 && x18 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && x16 && ~x7 && ~x12 && ~x13 && x18 && ~x14 )
						nx_state = s118;
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && x16 && ~x7 && ~x12 && ~x13 && ~x18 )
						nx_state = s118;
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && ~x16 && x11 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s689;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && ~x16 && x11 && ~x7 && x12 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && ~x16 && x11 && ~x7 && ~x12 )
						begin
							y4 = 1'b1;	
							nx_state = s834;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && ~x16 && ~x11 && x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s384;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && ~x16 && ~x11 && ~x4 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && ~x16 && ~x11 && ~x4 && ~x2 && x12 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s850;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && ~x16 && ~x11 && ~x4 && ~x2 && x12 && ~x7 )
						begin
							y4 = 1'b1;	
							nx_state = s834;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && ~x16 && ~x11 && ~x4 && ~x2 && ~x12 && x7 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s566;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && x15 && ~x16 && ~x11 && ~x4 && ~x2 && ~x12 && ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && ~x15 && x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s384;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && x7 && x12 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && x7 && x12 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s834;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && x7 && ~x12 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && x12 && x11 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && x12 && x11 && ~x2 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && x12 && ~x11 && x9 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && x12 && ~x11 && x9 && ~x2 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && x12 && ~x11 && ~x9 )
						nx_state = s1;
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && x11 && x10 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && x11 && x10 && ~x2 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && x11 && ~x10 )
						nx_state = s1;
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && ~x11 && x8 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && ~x11 && x8 && ~x2 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && ~x11 && ~x8 )
						nx_state = s1;
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && ~x16 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && ~x16 && ~x2 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s834;
						end
					else if( ~x70 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && ~x16 && ~x2 && ~x7 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( ~x70 && x65 && ~x61 && x60 && x15 && x16 && x7 && x12 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x70 && x65 && ~x61 && x60 && x15 && x16 && x7 && ~x12 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && x65 && ~x61 && x60 && x15 && x16 && ~x7 && x12 && x14 && x11 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s251;
						end
					else if( ~x70 && x65 && ~x61 && x60 && x15 && x16 && ~x7 && x12 && x14 && ~x11 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x70 && x65 && ~x61 && x60 && x15 && x16 && ~x7 && x12 && ~x14 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x61 && x60 && x15 && x16 && ~x7 && x12 && ~x14 && x18 && ~x13 )
						nx_state = s118;
					else if( ~x70 && x65 && ~x61 && x60 && x15 && x16 && ~x7 && x12 && ~x14 && ~x18 )
						nx_state = s118;
					else if( ~x70 && x65 && ~x61 && x60 && x15 && x16 && ~x7 && ~x12 && x13 && x11 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s564;
						end
					else if( ~x70 && x65 && ~x61 && x60 && x15 && x16 && ~x7 && ~x12 && x13 && ~x11 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x70 && x65 && ~x61 && x60 && x15 && x16 && ~x7 && ~x12 && ~x13 && x18 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x61 && x60 && x15 && x16 && ~x7 && ~x12 && ~x13 && x18 && ~x14 )
						nx_state = s118;
					else if( ~x70 && x65 && ~x61 && x60 && x15 && x16 && ~x7 && ~x12 && ~x13 && ~x18 )
						nx_state = s118;
					else if( ~x70 && x65 && ~x61 && x60 && x15 && ~x16 && x11 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s689;
						end
					else if( ~x70 && x65 && ~x61 && x60 && x15 && ~x16 && x11 && ~x7 && x12 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && x65 && ~x61 && x60 && x15 && ~x16 && x11 && ~x7 && ~x12 )
						begin
							y4 = 1'b1;	
							nx_state = s834;
						end
					else if( ~x70 && x65 && ~x61 && x60 && x15 && ~x16 && ~x11 && x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s384;
						end
					else if( ~x70 && x65 && ~x61 && x60 && x15 && ~x16 && ~x11 && ~x4 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && ~x61 && x60 && x15 && ~x16 && ~x11 && ~x4 && ~x2 && x12 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s850;
						end
					else if( ~x70 && x65 && ~x61 && x60 && x15 && ~x16 && ~x11 && ~x4 && ~x2 && x12 && ~x7 )
						begin
							y4 = 1'b1;	
							nx_state = s834;
						end
					else if( ~x70 && x65 && ~x61 && x60 && x15 && ~x16 && ~x11 && ~x4 && ~x2 && ~x12 && x7 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s566;
						end
					else if( ~x70 && x65 && ~x61 && x60 && x15 && ~x16 && ~x11 && ~x4 && ~x2 && ~x12 && ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x61 && x60 && ~x15 && x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s384;
						end
					else if( ~x70 && x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && x7 && x12 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && x7 && x12 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s834;
						end
					else if( ~x70 && x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && x7 && ~x12 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x70 && x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && x12 && x11 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && x12 && x11 && ~x2 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && x12 && ~x11 && x9 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && x12 && ~x11 && x9 && ~x2 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && x12 && ~x11 && ~x9 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && x11 && x10 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && x11 && x10 && ~x2 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && x11 && ~x10 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && ~x11 && x8 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && ~x11 && x8 && ~x2 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && ~x11 && ~x8 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x61 && x60 && ~x15 && ~x4 && ~x16 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && ~x61 && x60 && ~x15 && ~x4 && ~x16 && ~x2 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s834;
						end
					else if( ~x70 && x65 && ~x61 && x60 && ~x15 && ~x4 && ~x16 && ~x2 && ~x7 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( ~x70 && x65 && ~x61 && ~x60 && x62 )
						nx_state = s47;
					else if( ~x70 && x65 && ~x61 && ~x60 && ~x62 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x70 && ~x65 && x15 && x66 && x21 && x10 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s274;
						end
					else if( ~x70 && ~x65 && x15 && x66 && x21 && ~x10 && x12 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x70 && ~x65 && x15 && x66 && x21 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s124;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && x10 && x23 && x16 && x12 )
						begin
							y14 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && x10 && x23 && x16 && ~x12 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && x10 && x23 && ~x16 && x11 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s851;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && x10 && x23 && ~x16 && ~x11 && x12 )
						begin
							y14 = 1'b1;	
							nx_state = s124;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && x10 && x23 && ~x16 && ~x11 && ~x12 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && x10 && x23 && ~x16 && ~x11 && ~x12 && ~x2 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && x10 && x23 && ~x16 && ~x11 && ~x12 && ~x2 && ~x4 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s275;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && x10 && ~x23 && x11 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && x10 && ~x23 && ~x11 && x12 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && x10 && ~x23 && ~x11 && ~x12 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && x11 && x16 && x12 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s274;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && x11 && x16 && ~x12 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && x11 && ~x16 && x12 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && x11 && ~x16 && ~x12 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && x16 && x12 && x13 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s852;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && x16 && x12 && ~x13 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && x16 && x12 && ~x13 && x17 && ~x14 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && x16 && x12 && ~x13 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && x16 && ~x12 && x14 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s852;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && x16 && ~x12 && ~x14 && x17 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && x16 && ~x12 && ~x14 && x17 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && x16 && ~x12 && ~x14 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && ~x16 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && ~x16 && ~x2 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && ~x16 && ~x2 && ~x4 && x12 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && ~x16 && ~x2 && ~x4 && ~x12 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s367;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && ~x23 && x12 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && ~x23 && x12 && ~x11 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && ~x23 && ~x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && x9 && x7 && x23 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && x9 && x7 && ~x23 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && x9 && ~x7 && x8 && x23 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && x9 && ~x7 && x8 && ~x23 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s358;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && x9 && ~x7 && ~x8 && x13 && x23 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s853;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && x9 && ~x7 && ~x8 && x13 && ~x23 )
						begin
							y7 = 1'b1;	
							nx_state = s747;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && x9 && ~x7 && ~x8 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && ~x9 && x7 && x23 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && ~x9 && x7 && ~x23 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && ~x9 && ~x7 && x8 && x23 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s358;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && ~x9 && ~x7 && x8 && ~x23 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s851;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && ~x9 && ~x7 && ~x8 && x14 && x23 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s853;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && ~x9 && ~x7 && ~x8 && x14 && ~x23 )
						begin
							y7 = 1'b1;	
							nx_state = s747;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && ~x9 && ~x7 && ~x8 && ~x14 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && x7 && x9 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && x7 && ~x9 && x8 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && x7 && ~x9 && ~x8 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && x7 && ~x9 && ~x8 && ~x2 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && x7 && ~x9 && ~x8 && ~x2 && ~x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s357;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && ~x7 && x8 && x9 && x23 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s363;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && ~x7 && x8 && x9 && ~x23 )
						begin
							y14 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && ~x7 && x8 && ~x9 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && ~x7 && ~x8 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && ~x7 && ~x8 && ~x2 && x3 && x23 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && ~x7 && ~x8 && ~x2 && x3 && ~x23 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && ~x7 && ~x8 && ~x2 && ~x3 && x9 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && ~x7 && ~x8 && ~x2 && ~x3 && ~x9 && x23 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s365;
						end
					else if( ~x70 && ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && ~x7 && ~x8 && ~x2 && ~x3 && ~x9 && ~x23 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x65 && x15 && ~x66 && x8 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x65 && x15 && ~x66 && ~x8 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s781;
						end
					else if( ~x70 && ~x65 && x15 && ~x66 && ~x8 && ~x6 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && x21 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && x12 && x8 && x2 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s365;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && x12 && x8 && ~x2 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && x12 && x8 && ~x2 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && x12 && x8 && ~x2 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && x12 && x8 && ~x2 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && x12 && ~x8 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && x12 && ~x8 && ~x2 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && x12 && ~x8 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && ~x12 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && ~x12 && ~x2 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && ~x12 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && ~x23 && x12 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && ~x23 && ~x12 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s365;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && x7 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && x7 && ~x2 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && x7 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && ~x7 && x11 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && ~x7 && x11 && ~x2 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && ~x7 && x11 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && ~x7 && ~x11 && x2 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s365;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && ~x7 && ~x11 && ~x2 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && ~x7 && ~x11 && ~x2 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && ~x7 && ~x11 && ~x2 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && ~x7 && ~x11 && ~x2 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && x11 && x9 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && x11 && x9 && ~x2 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && x11 && x9 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && x11 && ~x9 && x2 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s365;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && x11 && ~x9 && ~x2 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && x11 && ~x9 && ~x2 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && x11 && ~x9 && ~x2 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && x11 && ~x9 && ~x2 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && ~x11 && x8 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && ~x11 && x8 && ~x2 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && ~x11 && x8 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && ~x11 && ~x8 && x2 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s365;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && ~x11 && ~x8 && ~x2 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && ~x11 && ~x8 && ~x2 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && ~x11 && ~x8 && ~x2 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && ~x11 && ~x8 && ~x2 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && ~x23 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && x7 && x11 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && x7 && ~x11 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && x7 && ~x11 && ~x2 && x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && x7 && ~x11 && ~x2 && x23 && ~x3 )
						begin
							y14 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && x7 && ~x11 && ~x2 && ~x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && x7 && ~x11 && ~x2 && ~x23 && ~x3 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && x10 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && x10 && ~x2 && x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && x10 && ~x2 && x23 && ~x3 )
						begin
							y14 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && x10 && ~x2 && ~x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && x10 && ~x2 && ~x23 && ~x3 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && ~x10 && x8 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && ~x10 && x8 && ~x2 && x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && ~x10 && x8 && ~x2 && x23 && ~x3 )
						begin
							y14 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && ~x10 && x8 && ~x2 && ~x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && ~x10 && x8 && ~x2 && ~x23 && ~x3 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && ~x10 && ~x8 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && x7 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && x7 && ~x2 && x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && x7 && ~x2 && x23 && ~x3 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && x7 && ~x2 && ~x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && x7 && ~x2 && ~x23 && ~x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && x8 && x12 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && x8 && x12 && ~x2 && x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && x8 && x12 && ~x2 && x23 && ~x3 )
						begin
							y14 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && x8 && x12 && ~x2 && ~x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && x8 && x12 && ~x2 && ~x23 && ~x3 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && x8 && ~x12 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && x8 && ~x12 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && x8 && ~x12 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && x8 && ~x12 && x23 && ~x19 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && x8 && ~x12 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && ~x8 && x11 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && ~x8 && x11 && ~x2 && x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && ~x8 && x11 && ~x2 && x23 && ~x3 )
						begin
							y14 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && ~x8 && x11 && ~x2 && ~x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && ~x8 && x11 && ~x2 && ~x23 && ~x3 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && ~x8 && ~x11 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x15 && x16 && ~x66 && x8 && x7 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && ~x66 && x8 && ~x7 && x9 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && ~x66 && x8 && ~x7 && ~x9 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && ~x66 && x8 && ~x7 && ~x9 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && ~x66 && x8 && ~x7 && ~x9 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x15 && x16 && ~x66 && x8 && ~x7 && ~x9 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x15 && x16 && ~x66 && ~x8 && x7 && x11 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && ~x66 && ~x8 && x7 && ~x11 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && ~x66 && ~x8 && x7 && ~x11 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && ~x66 && ~x8 && x7 && ~x11 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x15 && x16 && ~x66 && ~x8 && x7 && ~x11 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x15 && x16 && ~x66 && ~x8 && ~x7 && x10 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && ~x66 && ~x8 && ~x7 && ~x10 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && ~x66 && ~x8 && ~x7 && ~x10 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x70 && ~x65 && ~x15 && x16 && ~x66 && ~x8 && ~x7 && ~x10 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x15 && x16 && ~x66 && ~x8 && ~x7 && ~x10 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x15 && ~x16 && x66 && x21 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s357;
						end
					else if( ~x70 && ~x65 && ~x15 && ~x16 && x66 && ~x21 && x22 && x23 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( ~x70 && ~x65 && ~x15 && ~x16 && x66 && ~x21 && x22 && x23 && ~x2 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x70 && ~x65 && ~x15 && ~x16 && x66 && ~x21 && x22 && x23 && ~x2 && ~x4 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x65 && ~x15 && ~x16 && x66 && ~x21 && x22 && ~x23 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s151;
						end
					else if( ~x70 && ~x65 && ~x15 && ~x16 && x66 && ~x21 && ~x22 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( ~x70 && ~x65 && ~x15 && ~x16 && x66 && ~x21 && ~x22 && ~x2 && x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x70 && ~x65 && ~x15 && ~x16 && x66 && ~x21 && ~x22 && ~x2 && x23 && ~x3 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s851;
						end
					else if( ~x70 && ~x65 && ~x15 && ~x16 && x66 && ~x21 && ~x22 && ~x2 && ~x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x65 && ~x15 && ~x16 && x66 && ~x21 && ~x22 && ~x2 && ~x23 && ~x3 )
						begin
							y14 = 1'b1;	
							nx_state = s124;
						end
					else if( ~x70 && ~x65 && ~x15 && ~x16 && ~x66 && x6 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x70 && ~x65 && ~x15 && ~x16 && ~x66 && ~x6 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else nx_state = s146;
				s147 : if( x70 && x63 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x70 && x63 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x70 && x63 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x70 && x63 && ~x1 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && x66 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x70 && ~x63 && x64 && x66 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x70 && ~x63 && x64 && x66 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && x66 && ~x14 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && ~x66 && x12 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x70 && ~x63 && x64 && ~x66 && x12 && ~x8 && x7 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x70 && ~x63 && x64 && ~x66 && x12 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && ~x66 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x67 && x24 && x23 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x67 && x24 && ~x23 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x70 && ~x63 && ~x64 && x67 && x24 && ~x23 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x70 && ~x63 && ~x64 && x67 && x24 && ~x23 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x67 && x24 && ~x23 && ~x20 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x67 && ~x24 && x11 && x12 && x23 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x63 && ~x64 && x67 && ~x24 && x11 && x12 && ~x23 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x70 && ~x63 && ~x64 && x67 && ~x24 && x11 && ~x12 && x13 && x23 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x63 && ~x64 && x67 && ~x24 && x11 && ~x12 && x13 && ~x23 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x70 && ~x63 && ~x64 && x67 && ~x24 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x67 && ~x24 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && ~x67 && x28 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x63 && ~x64 && ~x67 && x28 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x63 && ~x64 && ~x67 && x28 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && ~x67 && x28 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && ~x67 && ~x28 )
						begin
							y8 = 1'b1;	
							nx_state = s783;
						end
					else if( ~x70 && x65 && x66 && x67 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && x66 && x67 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && x66 && x67 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && x67 && x22 && ~x17 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && x67 && ~x22 && x18 && x13 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && x65 && x66 && x67 && ~x22 && x18 && x13 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x65 && x66 && x67 && ~x22 && x18 && ~x13 && x12 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && x65 && x66 && x67 && ~x22 && x18 && ~x13 && x12 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x65 && x66 && x67 && ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && x67 && ~x22 && ~x18 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && ~x67 && x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && x66 && ~x67 && x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && x66 && ~x67 && x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && ~x67 && x21 && x20 && ~x17 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && ~x67 && x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x65 && x66 && ~x67 && x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x65 && x66 && ~x67 && x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && ~x67 && x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && ~x67 && ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x65 && x66 && ~x67 && ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && ~x67 && ~x21 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && x65 && ~x66 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x22 && x23 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x22 && x23 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x22 && x23 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x22 && x23 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x22 && x23 && ~x19 && ~x17 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x22 && ~x23 && x18 && x14 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x22 && ~x23 && x18 && ~x14 && x13 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x22 && x23 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x22 && x23 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x22 && x23 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x22 && x23 && ~x20 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x22 && ~x23 && x15 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x70 && x65 && ~x66 && ~x21 && ~x22 && ~x23 && ~x15 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s495;
						end
					else if( ~x70 && ~x65 && x66 && x67 && x68 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x65 && x66 && x67 && x68 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x65 && x66 && x67 && x68 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && x67 && x68 && x21 && ~x19 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && x67 && x68 && ~x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s224;
						end
					else if( ~x70 && ~x65 && x66 && x67 && ~x68 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && ~x65 && x66 && x67 && ~x68 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && ~x65 && x66 && x67 && ~x68 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && x67 && ~x68 && x62 && ~x61 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && ~x67 && x21 && x68 )
						begin
							y8 = 1'b1;	y18 = 1'b1;	
							nx_state = s152;
						end
					else if( ~x70 && ~x65 && x66 && ~x67 && x21 && ~x68 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( ~x70 && ~x65 && x66 && ~x67 && ~x21 && x68 && x22 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x70 && ~x65 && x66 && ~x67 && ~x21 && x68 && x22 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x70 && ~x65 && x66 && ~x67 && ~x21 && x68 && x22 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && ~x67 && ~x21 && x68 && x22 && ~x7 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && ~x67 && ~x21 && x68 && ~x22 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x70 && ~x65 && x66 && ~x67 && ~x21 && x68 && ~x22 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x70 && ~x65 && x66 && ~x67 && ~x21 && x68 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && ~x67 && ~x21 && x68 && ~x22 && ~x4 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && ~x67 && ~x21 && ~x68 && x23 && x22 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && ~x65 && x66 && ~x67 && ~x21 && ~x68 && x23 && ~x22 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x70 && ~x65 && x66 && ~x67 && ~x21 && ~x68 && x23 && ~x22 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x70 && ~x65 && x66 && ~x67 && ~x21 && ~x68 && x23 && ~x22 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && ~x67 && ~x21 && ~x68 && x23 && ~x22 && ~x19 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && ~x67 && ~x21 && ~x68 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x65 && ~x66 && x68 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && ~x66 && x68 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && ~x66 && x68 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && x68 && x20 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && x68 && ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x70 && ~x65 && ~x66 && x68 && ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x70 && ~x65 && ~x66 && x68 && ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && x68 && ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && x68 && ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x70 && ~x65 && ~x66 && x68 && ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x70 && ~x65 && ~x66 && x68 && ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && x68 && ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && ~x68 && x24 && x26 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x68 && x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x68 && x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x68 && x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && ~x68 && x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && x25 && x19 && ~x14 && ~x13 && x26 )
						nx_state = s147;
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && x25 && x19 && ~x14 && ~x13 && ~x26 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && x4 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && x19 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && x20 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && ~x20 && x21 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && ~x20 && ~x21 && x22 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && ~x20 && ~x21 && ~x22 && x16 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && ~x20 && ~x21 && ~x22 && x16 && ~x11 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && ~x20 && ~x21 && ~x22 && x16 && ~x11 && ~x12 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && ~x20 && ~x21 && ~x22 && x16 && ~x11 && ~x12 && ~x10 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && ~x20 && ~x21 && ~x22 && ~x16 && x17 && x10 && x12 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && ~x20 && ~x21 && ~x22 && ~x16 && x17 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && ~x20 && ~x21 && ~x22 && ~x16 && x17 && ~x10 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && ~x20 && ~x21 && ~x22 && ~x16 && ~x17 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else nx_state = s147;
				s148 : if( x70 && x64 && x21 && x17 && x16 && x19 && x11 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x70 && x64 && x21 && x17 && x16 && x19 && ~x11 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && x64 && x21 && x17 && x16 && ~x19 && x18 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x70 && x64 && x21 && x17 && x16 && ~x19 && ~x18 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && x64 && x21 && x17 && ~x16 && x11 )
						begin
							y3 = 1'b1;	
							nx_state = s788;
						end
					else if( x70 && x64 && x21 && x17 && ~x16 && ~x11 )
						begin
							y32 = 1'b1;	
							nx_state = s854;
						end
					else if( x70 && x64 && x21 && ~x17 && x16 && x19 && x14 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x70 && x64 && x21 && ~x17 && x16 && x19 && ~x14 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && x64 && x21 && ~x17 && x16 && ~x19 && x13 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x70 && x64 && x21 && ~x17 && x16 && ~x19 && ~x13 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && x64 && x21 && ~x17 && ~x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && x64 && ~x21 )
						begin
							y30 = 1'b1;	
							nx_state = s416;
						end
					else if( x70 && ~x64 && x30 && x31 && x14 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && ~x64 && x30 && x31 && ~x14 )
						begin
							y47 = 1'b1;	y54 = 1'b1;	y61 = 1'b1;	
							y68 = 1'b1;	
							nx_state = s855;
						end
					else if( x70 && ~x64 && x30 && ~x31 && x14 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x64 && x30 && ~x31 && x14 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x64 && x30 && ~x31 && x14 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x70 && ~x64 && x30 && ~x31 && x14 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x64 && x30 && ~x31 && ~x14 )
						begin
							y47 = 1'b1;	y53 = 1'b1;	y61 = 1'b1;	
							y72 = 1'b1;	
							nx_state = s856;
						end
					else if( x70 && ~x64 && ~x30 )
						begin
							y47 = 1'b1;	y49 = 1'b1;	y58 = 1'b1;	
							y61 = 1'b1;	y68 = 1'b1;	
							nx_state = s857;
						end
					else if( ~x70 && x65 && x66 && x61 && x60 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x65 && x66 && x61 && x60 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x65 && x66 && x61 && x60 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( ~x70 && x65 && x66 && x61 && x60 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( ~x70 && x65 && x66 && x61 && ~x60 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && x66 && x61 && ~x60 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && x66 && x61 && ~x60 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && x61 && ~x60 && x62 && ~x18 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && x61 && ~x60 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && x66 && x61 && ~x60 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && x66 && x61 && ~x60 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( ~x70 && x65 && x66 && x61 && ~x60 && ~x62 && ~x18 )
						nx_state = s118;
					else if( ~x70 && x65 && x66 && ~x61 && x60 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && x66 && ~x61 && x60 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && x66 && ~x61 && x60 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( ~x70 && x65 && x66 && ~x61 && x60 && ~x18 )
						nx_state = s118;
					else if( ~x70 && x65 && x66 && ~x61 && ~x60 && x62 )
						nx_state = s47;
					else if( ~x70 && x65 && x66 && ~x61 && ~x60 && ~x62 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s566;
						end
					else if( ~x70 && x65 && ~x66 && x67 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x67 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x67 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x67 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && x22 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && ~x22 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x70 && ~x65 && x21 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x70 && ~x65 && ~x21 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x70 && ~x65 && ~x21 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && ~x7 )
						nx_state = s1;
					else nx_state = s148;
				s149 : if( x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x21 && x22 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x10 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s792;
						end
					else if( ~x21 && ~x22 && ~x10 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x21 && ~x22 && ~x10 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x21 && ~x22 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x10 && ~x4 )
						nx_state = s1;
					else nx_state = s149;
				s150 : if( x22 )
						nx_state = s1;
					else if( ~x22 && x21 )
						nx_state = s1;
					else if( ~x22 && ~x21 && x23 && x15 && x7 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s151;
						end
					else if( ~x22 && ~x21 && x23 && x15 && ~x7 && x9 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x22 && ~x21 && x23 && x15 && ~x7 && ~x9 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x22 && ~x21 && x23 && ~x15 && x7 && x9 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s274;
						end
					else if( ~x22 && ~x21 && x23 && ~x15 && x7 && ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x22 && ~x21 && x23 && ~x15 && ~x7 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s274;
						end
					else if( ~x22 && ~x21 && ~x23 )
						begin
							y14 = 1'b1;	
							nx_state = s366;
						end
					else nx_state = s150;
				s151 : if( x21 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s367;
						end
					else if( ~x21 && x22 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x19 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else nx_state = s151;
				s152 : if( x21 && x66 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( x21 && ~x66 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x21 && ~x66 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x21 && ~x66 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x21 && ~x66 && ~x3 )
						nx_state = s1;
					else if( ~x21 && x66 && x22 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x21 && x66 && ~x22 && x16 && x15 && x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s336;
						end
					else if( ~x21 && x66 && ~x22 && x16 && x15 && ~x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s828;
						end
					else if( ~x21 && x66 && ~x22 && x16 && ~x15 && x10 )
						begin
							y2 = 1'b1;	y16 = 1'b1;	y24 = 1'b1;	
							nx_state = s270;
						end
					else if( ~x21 && x66 && ~x22 && x16 && ~x15 && ~x10 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s267;
						end
					else if( ~x21 && x66 && ~x22 && ~x16 && x17 && x10 && x15 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s336;
						end
					else if( ~x21 && x66 && ~x22 && ~x16 && x17 && x10 && ~x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s827;
						end
					else if( ~x21 && x66 && ~x22 && ~x16 && x17 && ~x10 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x66 && ~x22 && ~x16 && ~x17 && x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s336;
						end
					else if( ~x21 && x66 && ~x22 && ~x16 && ~x17 && ~x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s829;
						end
					else if( ~x21 && ~x66 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x21 && ~x66 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x21 && ~x66 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && ~x66 && ~x8 )
						nx_state = s1;
					else nx_state = s152;
				s153 : if( x70 && x62 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x70 && x62 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x70 && x62 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( x70 && x62 && ~x27 )
						nx_state = s1;
					else if( x70 && ~x62 && x65 && x64 && x63 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x70 && ~x62 && x65 && x64 && x63 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x70 && ~x62 && x65 && x64 && x63 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( x70 && ~x62 && x65 && x64 && x63 && ~x22 )
						nx_state = s1;
					else if( x70 && ~x62 && x65 && x64 && ~x63 && x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x70 && ~x62 && x65 && x64 && ~x63 && x10 && ~x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x70 && ~x62 && x65 && x64 && ~x63 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x62 && x65 && x64 && ~x63 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x62 && x65 && ~x64 && x63 && x66 && x30 && x8 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( x70 && ~x62 && x65 && ~x64 && x63 && x66 && x30 && ~x8 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x70 && ~x62 && x65 && ~x64 && x63 && x66 && ~x30 )
						begin
							y17 = 1'b1;	
							nx_state = s3;
						end
					else if( x70 && ~x62 && x65 && ~x64 && x63 && ~x66 )
						nx_state = s1;
					else if( x70 && ~x62 && x65 && ~x64 && ~x63 && x66 && x23 && x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x62 && x65 && ~x64 && ~x63 && x66 && x23 && x11 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x62 && x65 && ~x64 && ~x63 && x66 && x23 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x70 && ~x62 && x65 && ~x64 && ~x63 && x66 && x23 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && x65 && ~x64 && ~x63 && x66 && ~x23 && x24 )
						nx_state = s1;
					else if( x70 && ~x62 && x65 && ~x64 && ~x63 && x66 && ~x23 && ~x24 && x11 && x12 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x70 && ~x62 && x65 && ~x64 && ~x63 && x66 && ~x23 && ~x24 && x11 && ~x12 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x70 && ~x62 && x65 && ~x64 && ~x63 && x66 && ~x23 && ~x24 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x70 && ~x62 && x65 && ~x64 && ~x63 && x66 && ~x23 && ~x24 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && x65 && ~x64 && ~x63 && ~x66 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x62 && x65 && ~x64 && ~x63 && ~x66 && x20 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x62 && x65 && ~x64 && ~x63 && ~x66 && x20 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x62 && x65 && ~x64 && ~x63 && ~x66 && ~x20 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x65 && x64 && x63 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x70 && ~x62 && ~x65 && x64 && x63 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x70 && ~x62 && ~x65 && x64 && x63 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x65 && x64 && x63 && ~x14 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x65 && x64 && ~x63 && x66 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x65 && x64 && ~x63 && x66 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x65 && x64 && ~x63 && x66 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x65 && x64 && ~x63 && x66 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x65 && x64 && ~x63 && ~x66 && x67 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x70 && ~x62 && ~x65 && x64 && ~x63 && ~x66 && x67 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x70 && ~x62 && ~x65 && x64 && ~x63 && ~x66 && x67 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x65 && x64 && ~x63 && ~x66 && x67 && ~x14 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x65 && x64 && ~x63 && ~x66 && ~x67 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x70 && ~x62 && ~x65 && x64 && ~x63 && ~x66 && ~x67 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x70 && ~x62 && ~x65 && x64 && ~x63 && ~x66 && ~x67 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x65 && x64 && ~x63 && ~x66 && ~x67 && ~x18 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x65 && ~x64 && x63 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x70 && ~x62 && ~x65 && ~x64 && ~x63 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && x68 && x21 && x20 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 && x18 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y21 = 1'b1;	
							nx_state = s599;
						end
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 && ~x18 && x15 && x10 && x11 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s600;
						end
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 && ~x18 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s601;
						end
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 && ~x18 && x15 && x10 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y13 = 1'b1;	
							nx_state = s600;
						end
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 && ~x18 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 && ~x18 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s602;
						end
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && x10 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && x10 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && x10 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && x10 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && ~x10 && x12 && x11 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s603;
						end
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && ~x10 && x12 && ~x11 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && ~x10 && x12 && ~x11 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && ~x10 && x12 && ~x11 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && ~x10 && x12 && ~x11 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && ~x10 && ~x12 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && ~x10 && ~x12 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && ~x10 && ~x12 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && ~x10 && ~x12 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s604;
						end
					else if( ~x70 && x65 && x66 && x68 && ~x21 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && ~x68 && x60 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && x16 && x4 && x11 && x12 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s97;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && x16 && x4 && x11 && ~x12 && x13 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s858;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && x16 && x4 && x11 && ~x12 && ~x13 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && x16 && x4 && ~x11 && x13 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && x16 && x4 && ~x11 && ~x13 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && x16 && ~x4 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && x11 && x9 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && x11 && ~x9 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && x11 && ~x9 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && x11 && ~x9 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && x11 && ~x9 && ~x18 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && ~x11 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && ~x11 && ~x8 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && ~x11 && ~x8 && ~x12 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && ~x11 && ~x8 && ~x12 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && ~x11 && ~x8 && ~x12 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && ~x11 && ~x8 && ~x12 && ~x18 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && x11 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && ~x11 && x12 && x10 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && ~x11 && x12 && ~x10 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && ~x11 && x12 && ~x10 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && ~x11 && x12 && ~x10 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && ~x11 && x12 && ~x10 && ~x18 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && ~x11 && ~x12 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && ~x11 && ~x12 && ~x7 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && ~x11 && ~x12 && ~x7 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && ~x11 && ~x12 && ~x7 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && ~x11 && ~x12 && ~x7 && ~x18 )
						nx_state = s1;
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && ~x17 && x45 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && ~x17 && ~x45 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x65 && x66 && ~x68 && ~x60 && ~x61 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x67 && x21 && x68 && x18 )
						begin
							y14 = 1'b1;	y19 = 1'b1;	
							nx_state = s723;
						end
					else if( ~x70 && x65 && ~x66 && x67 && x21 && x68 && ~x18 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s724;
						end
					else if( ~x70 && x65 && ~x66 && x67 && x21 && ~x68 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x67 && x21 && ~x68 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x67 && x21 && ~x68 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x67 && x21 && ~x68 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && x22 && x68 && x8 && x23 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && x22 && x68 && x8 && x23 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && x22 && x68 && x8 && x23 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && x22 && x68 && x8 && ~x23 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && x22 && x68 && x8 && ~x23 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && x22 && x68 && x8 && ~x23 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && x22 && x68 && ~x8 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && x22 && ~x68 && x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && x22 && ~x68 && x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && x22 && ~x68 && x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && x22 && ~x68 && x19 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && x22 && ~x68 && ~x19 && x18 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && x22 && ~x68 && ~x19 && x18 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && x22 && ~x68 && ~x19 && x18 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && x22 && ~x68 && ~x19 && x18 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && x22 && ~x68 && ~x19 && ~x18 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && ~x22 && x68 && x23 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && ~x22 && x68 && x23 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && ~x22 && x68 && x23 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && ~x22 && x68 && x23 && ~x9 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && ~x22 && x68 && ~x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && ~x22 && x68 && ~x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && ~x22 && x68 && ~x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && ~x22 && x68 && ~x23 && ~x8 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && ~x22 && ~x68 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && ~x22 && ~x68 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && ~x22 && ~x68 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x67 && ~x21 && ~x22 && ~x68 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && x17 && x20 && x16 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && x17 && x20 && ~x16 )
						begin
							y24 = 1'b1;	
							nx_state = s259;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && x17 && ~x20 && x16 )
						begin
							y13 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	y29 = 1'b1;	y30 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s859;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && x17 && ~x20 && ~x16 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && ~x17 && x16 && x4 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s860;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && ~x17 && x16 && ~x4 )
						begin
							y10 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s861;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && ~x17 && ~x16 && x20 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && ~x17 && ~x16 && x20 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && ~x17 && ~x16 && x20 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && ~x17 && ~x16 && x20 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && ~x17 && ~x16 && ~x20 )
						begin
							y15 = 1'b1;	y28 = 1'b1;	
							nx_state = s862;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && x15 && x17 && x20 && x16 )
						begin
							y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && x15 && x17 && x20 && ~x16 )
						begin
							y4 = 1'b1;	y12 = 1'b1;	y27 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && x15 && x17 && ~x20 && x16 )
						begin
							y24 = 1'b1;	
							nx_state = s259;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && x15 && x17 && ~x20 && ~x16 )
						begin
							y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && x15 && ~x17 && x16 )
						begin
							y15 = 1'b1;	y28 = 1'b1;	
							nx_state = s862;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && x15 && ~x17 && ~x16 && x13 )
						begin
							y15 = 1'b1;	y28 = 1'b1;	
							nx_state = s862;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && x15 && ~x17 && ~x16 && ~x13 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && x15 && ~x17 && ~x16 && ~x13 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && x15 && ~x17 && ~x16 && ~x13 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && x15 && ~x17 && ~x16 && ~x13 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && x17 && x6 && x16 && x7 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && x17 && x6 && x16 && ~x7 && x5 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && x17 && x6 && x16 && ~x7 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && x17 && x6 && ~x16 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && x17 && ~x6 && x7 && x16 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && x17 && ~x6 && x7 && ~x16 && x5 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && x17 && ~x6 && x7 && ~x16 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && x17 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && ~x17 && x16 && x12 )
						begin
							y15 = 1'b1;	y28 = 1'b1;	
							nx_state = s862;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && ~x17 && x16 && ~x12 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && ~x17 && x16 && ~x12 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && ~x17 && x16 && ~x12 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && ~x17 && x16 && ~x12 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && ~x17 && ~x16 && x11 )
						begin
							y15 = 1'b1;	y28 = 1'b1;	
							nx_state = s862;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && ~x17 && ~x16 && ~x11 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && ~x17 && ~x16 && ~x11 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && ~x17 && ~x16 && ~x11 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && ~x17 && ~x16 && ~x11 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && x20 && x14 && x13 )
						begin
							y10 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s861;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && x20 && x14 && ~x13 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && x20 && ~x14 && x13 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	y19 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s861;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && x20 && ~x14 && ~x13 && x6 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && x20 && ~x14 && ~x13 && ~x6 && x5 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && x20 && ~x14 && ~x13 && ~x6 && x5 && ~x7 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && x20 && ~x14 && ~x13 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && ~x20 && x15 && x14 )
						begin
							y10 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s861;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && ~x20 && x15 && ~x14 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && ~x20 && ~x15 && x14 )
						begin
							y15 = 1'b1;	y28 = 1'b1;	
							nx_state = s862;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && ~x20 && ~x15 && ~x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && x13 && x12 && x14 )
						begin
							y15 = 1'b1;	y28 = 1'b1;	
							nx_state = s862;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && x13 && x12 && ~x14 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && x13 && x12 && ~x14 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && x13 && x12 && ~x14 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && x13 && x12 && ~x14 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && x13 && ~x12 )
						begin
							y15 = 1'b1;	y28 = 1'b1;	
							nx_state = s862;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && ~x13 && x11 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && ~x13 && x11 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && ~x13 && x11 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && ~x13 && x11 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && ~x13 && ~x11 )
						begin
							y15 = 1'b1;	y28 = 1'b1;	
							nx_state = s862;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && x14 && x13 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s860;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && x14 && ~x13 && x15 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s860;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && x14 && ~x13 && ~x15 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && x14 && ~x13 && ~x15 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && x14 && ~x13 && ~x15 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && x14 && ~x13 && ~x15 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && ~x14 && x15 && x12 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s860;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && ~x14 && x15 && ~x12 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && ~x14 && x15 && ~x12 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && ~x14 && x15 && ~x12 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && ~x14 && x15 && ~x12 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && ~x14 && ~x15 && x11 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s860;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && ~x14 && ~x15 && ~x11 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && ~x14 && ~x15 && ~x11 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && ~x14 && ~x15 && ~x11 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && ~x14 && ~x15 && ~x11 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && x14 && x15 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && x14 && ~x15 && x16 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && x14 && ~x15 && ~x16 && x4 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s860;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && x14 && ~x15 && ~x16 && ~x4 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s864;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && ~x14 && x16 && x15 && x13 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && ~x14 && x16 && x15 && ~x13 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	y32 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && ~x14 && x16 && ~x15 && x4 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s860;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && ~x14 && x16 && ~x15 && ~x4 )
						begin
							y4 = 1'b1;	y17 = 1'b1;	y29 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && ~x14 && ~x16 && x15 )
						begin
							y4 = 1'b1;	y29 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && ~x14 && ~x16 && ~x15 && x4 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	y21 = 1'b1;	y28 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && ~x14 && ~x16 && ~x15 && ~x4 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && ~x19 && x16 && x14 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	y21 = 1'b1;	y28 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && ~x19 && x16 && ~x14 && x4 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && ~x19 && x16 && ~x14 && ~x4 )
						begin
							y16 = 1'b1;	y28 = 1'b1;	
							nx_state = s865;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && ~x19 && ~x16 && x13 && x14 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	y21 = 1'b1;	y28 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && ~x19 && ~x16 && x13 && x14 && ~x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && ~x19 && ~x16 && x13 && ~x14 && x4 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && ~x19 && ~x16 && x13 && ~x14 && ~x4 )
						begin
							y4 = 1'b1;	y12 = 1'b1;	y27 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && ~x19 && ~x16 && ~x13 && x4 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && ~x19 && ~x16 && ~x13 && ~x4 )
						begin
							y24 = 1'b1;	
							nx_state = s259;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && x14 && x19 && x15 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && x14 && x19 && ~x15 && x16 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && x14 && x19 && ~x15 && ~x16 && x4 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s860;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && x14 && x19 && ~x15 && ~x16 && ~x4 )
						begin
							y4 = 1'b1;	y29 = 1'b1;	y32 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && x14 && ~x19 && x16 )
						begin
							y24 = 1'b1;	
							nx_state = s259;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && x14 && ~x19 && ~x16 && x15 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && x14 && ~x19 && ~x16 && x15 && ~x13 )
						begin
							y4 = 1'b1;	y12 = 1'b1;	y27 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && x14 && ~x19 && ~x16 && ~x15 )
						begin
							y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && x15 && x16 && x19 && x13 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && x15 && x16 && x19 && ~x13 )
						begin
							y4 = 1'b1;	y29 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && x15 && x16 && ~x19 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && x15 && ~x16 && x4 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s860;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && x15 && ~x16 && ~x4 && x19 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && x15 && ~x16 && ~x4 && ~x19 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && ~x15 && x4 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s860;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && ~x15 && ~x4 && x19 && x16 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && ~x15 && ~x4 && x19 && ~x16 )
						begin
							y4 = 1'b1;	y12 = 1'b1;	y27 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && ~x15 && ~x4 && ~x19 && x16 )
						begin
							y16 = 1'b1;	y28 = 1'b1;	
							nx_state = s865;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && ~x15 && ~x4 && ~x19 && ~x16 )
						begin
							y13 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	y29 = 1'b1;	y30 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s859;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && ~x17 && x4 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s860;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && ~x17 && ~x4 )
						begin
							y4 = 1'b1;	y17 = 1'b1;	
							nx_state = s235;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && ~x21 && x23 && x22 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && ~x21 && x23 && x22 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && ~x21 && x23 && x22 && ~x19 && ~x17 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && ~x21 && x23 && ~x22 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && ~x21 && x23 && ~x22 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && ~x21 && x23 && ~x22 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && ~x21 && x23 && ~x22 && ~x20 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x23 && x18 && x14 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x23 && x18 && x14 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x23 && x18 && ~x14 && x13 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x23 && x18 && ~x14 && x13 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x67 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && ~x65 && x67 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && ~x65 && x67 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x67 && x62 && ~x61 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x67 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x65 && x67 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && ~x65 && x67 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x65 && x67 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && ~x65 && x67 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x67 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x67 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && x67 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x65 && x67 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && x67 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x65 && x67 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x67 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x67 )
						nx_state = s1;
					else nx_state = s153;
				s154 : if( x69 && x21 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( x69 && ~x21 && x23 && x22 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s866;
						end
					else if( x69 && ~x21 && x23 && ~x22 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s150;
						end
					else if( x69 && ~x21 && ~x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s150;
						end
					else if( ~x69 && x44 && x10 && x12 && x23 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x69 && x44 && x10 && x12 && ~x23 && x4 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s867;
						end
					else if( ~x69 && x44 && x10 && x12 && ~x23 && ~x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && x44 && x10 && ~x12 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s868;
						end
					else if( ~x69 && x44 && ~x10 && x37 && x22 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							nx_state = s869;
						end
					else if( ~x69 && x44 && ~x10 && x37 && ~x22 && x2 && x11 && x42 )
						nx_state = s154;
					else if( ~x69 && x44 && ~x10 && x37 && ~x22 && x2 && x11 && ~x42 && x5 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && x44 && ~x10 && x37 && ~x22 && x2 && x11 && ~x42 && ~x5 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s870;
						end
					else if( ~x69 && x44 && ~x10 && x37 && ~x22 && x2 && ~x11 && x42 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( ~x69 && x44 && ~x10 && x37 && ~x22 && x2 && ~x11 && ~x42 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s867;
						end
					else if( ~x69 && x44 && ~x10 && x37 && ~x22 && ~x2 )
						begin
							y11 = 1'b1;	
							nx_state = s250;
						end
					else if( ~x69 && x44 && ~x10 && ~x37 && x11 && x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && x44 && ~x10 && ~x37 && x11 && ~x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( ~x69 && x44 && ~x10 && ~x37 && ~x11 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && ~x44 && x10 && x39 && x46 && x51 && x36 )
						nx_state = s154;
					else if( ~x69 && ~x44 && x10 && x39 && x46 && x51 && ~x36 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x69 && ~x44 && x10 && x39 && x46 && ~x51 && x36 )
						nx_state = s154;
					else if( ~x69 && ~x44 && x10 && x39 && x46 && ~x51 && ~x36 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && ~x44 && x10 && x39 && ~x46 && x36 )
						nx_state = s154;
					else if( ~x69 && ~x44 && x10 && x39 && ~x46 && ~x36 )
						begin
							y11 = 1'b1;	
							nx_state = s250;
						end
					else if( ~x69 && ~x44 && x10 && ~x39 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s871;
						end
					else if( ~x69 && ~x44 && ~x10 && x11 && x34 && x8 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( ~x69 && ~x44 && ~x10 && x11 && x34 && ~x8 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x69 && ~x44 && ~x10 && x11 && x34 && ~x8 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( ~x69 && ~x44 && ~x10 && x11 && ~x34 && x32 && x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( ~x69 && ~x44 && ~x10 && x11 && ~x34 && x32 && ~x7 && x54 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x69 && ~x44 && ~x10 && x11 && ~x34 && x32 && ~x7 && x54 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( ~x69 && ~x44 && ~x10 && x11 && ~x34 && x32 && ~x7 && ~x54 )
						begin
							y11 = 1'b1;	
							nx_state = s250;
						end
					else if( ~x69 && ~x44 && ~x10 && x11 && ~x34 && ~x32 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s870;
						end
					else if( ~x69 && ~x44 && ~x10 && ~x11 && x12 && x20 )
						begin
							y11 = 1'b1;	
							nx_state = s250;
						end
					else if( ~x69 && ~x44 && ~x10 && ~x11 && x12 && ~x20 && x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && ~x44 && ~x10 && ~x11 && x12 && ~x20 && ~x2 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s867;
						end
					else if( ~x69 && ~x44 && ~x10 && ~x11 && ~x12 && x13 && x36 && x3 && x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s868;
						end
					else if( ~x69 && ~x44 && ~x10 && ~x11 && ~x12 && x13 && x36 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( ~x69 && ~x44 && ~x10 && ~x11 && ~x12 && x13 && x36 && ~x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( ~x69 && ~x44 && ~x10 && ~x11 && ~x12 && x13 && ~x36 )
						begin
							y11 = 1'b1;	
							nx_state = s250;
						end
					else if( ~x69 && ~x44 && ~x10 && ~x11 && ~x12 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else nx_state = s154;
				s155 : if( x69 && x70 && x62 && x24 && x2 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && x70 && x62 && x24 && x2 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x69 && x70 && x62 && x24 && ~x2 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x69 && x70 && x62 && ~x24 && x2 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( x69 && x70 && x62 && ~x24 && ~x2 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( x69 && x70 && x62 && ~x24 && ~x2 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x69 && x70 && ~x62 && x19 && x18 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s873;
						end
					else if( x69 && x70 && ~x62 && x19 && ~x18 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s872;
						end
					else if( x69 && x70 && ~x62 && ~x19 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s873;
						end
					else if( x69 && ~x70 && x65 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && ~x70 && ~x65 && x22 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s357;
						end
					else if( x69 && ~x70 && ~x65 && ~x22 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s853;
						end
					else if( ~x69 && x70 && x61 && x16 && x19 && x33 )
						begin
							y10 = 1'b1;	
							nx_state = s841;
						end
					else if( ~x69 && x70 && x61 && x16 && x19 && ~x33 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( ~x69 && x70 && x61 && x16 && x19 && ~x33 && ~x13 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s840;
						end
					else if( ~x69 && x70 && x61 && x16 && ~x19 && x30 && x26 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s874;
						end
					else if( ~x69 && x70 && x61 && x16 && ~x19 && x30 && x26 && ~x1 && x9 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x69 && x70 && x61 && x16 && ~x19 && x30 && x26 && ~x1 && x9 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s875;
						end
					else if( ~x69 && x70 && x61 && x16 && ~x19 && x30 && x26 && ~x1 && ~x9 )
						nx_state = s155;
					else if( ~x69 && x70 && x61 && x16 && ~x19 && x30 && ~x26 && x3 )
						nx_state = s155;
					else if( ~x69 && x70 && x61 && x16 && ~x19 && x30 && ~x26 && ~x3 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s874;
						end
					else if( ~x69 && x70 && x61 && x16 && ~x19 && x30 && ~x26 && ~x3 && ~x1 && x9 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x69 && x70 && x61 && x16 && ~x19 && x30 && ~x26 && ~x3 && ~x1 && x9 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s875;
						end
					else if( ~x69 && x70 && x61 && x16 && ~x19 && x30 && ~x26 && ~x3 && ~x1 && ~x9 )
						nx_state = s155;
					else if( ~x69 && x70 && x61 && x16 && ~x19 && ~x30 )
						nx_state = s155;
					else if( ~x69 && x70 && x61 && ~x16 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( ~x69 && x70 && ~x61 && x28 && x57 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s733;
						end
					else if( ~x69 && x70 && ~x61 && x28 && ~x57 )
						nx_state = s155;
					else if( ~x69 && x70 && ~x61 && ~x28 && x27 && x8 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s733;
						end
					else if( ~x69 && x70 && ~x61 && ~x28 && x27 && ~x8 && x37 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( ~x69 && x70 && ~x61 && ~x28 && x27 && ~x8 && ~x37 )
						begin
							y10 = 1'b1;	
							nx_state = s841;
						end
					else if( ~x69 && x70 && ~x61 && ~x28 && ~x27 && x50 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x69 && x70 && ~x61 && ~x28 && ~x27 && ~x50 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x10 && x6 && x7 && x2 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x10 && x6 && x7 && x2 && ~x3 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x10 && x6 && x7 && x2 && ~x3 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x10 && x6 && x7 && ~x2 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x10 && x6 && ~x7 && x8 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x10 && x6 && ~x7 && ~x8 && x2 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x10 && x6 && ~x7 && ~x8 && x2 && ~x3 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x10 && x6 && ~x7 && ~x8 && x2 && ~x3 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x10 && x6 && ~x7 && ~x8 && ~x2 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x10 && ~x6 && x2 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x10 && ~x6 && ~x2 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x44 && x45 && ~x10 && x11 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x10 && x11 && ~x5 && x6 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x10 && x11 && ~x5 && ~x6 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x44 && ~x45 && x9 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x9 && x7 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x9 && ~x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							nx_state = s38;
						end
					else if( ~x69 && ~x70 && ~x44 && x10 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x44 && ~x10 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 && ~x5 && x6 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 && ~x5 && ~x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else nx_state = s155;
				s156 : if( x21 && x19 && x15 && x10 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s274;
						end
					else if( x21 && x19 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x21 && x19 && x15 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s124;
						end
					else if( x21 && x19 && ~x15 && x16 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x21 && x19 && ~x15 && ~x16 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s357;
						end
					else if( x21 && ~x19 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x21 && x23 )
						nx_state = s1;
					else if( ~x21 && ~x23 && x22 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x21 && ~x23 && ~x22 )
						nx_state = s1;
					else nx_state = s156;
				s157 : if( x21 && x66 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x21 && x66 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x21 && x66 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x21 && x66 && ~x9 )
						nx_state = s1;
					else if( x21 && ~x66 && x19 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s574;
						end
					else if( x21 && ~x66 && x19 && ~x12 && x17 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s574;
						end
					else if( x21 && ~x66 && x19 && ~x12 && ~x17 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s377;
						end
					else if( x21 && ~x66 && ~x19 && x20 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s574;
						end
					else if( x21 && ~x66 && ~x19 && x20 && ~x12 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s377;
						end
					else if( x21 && ~x66 && ~x19 && ~x20 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s573;
						end
					else if( x21 && ~x66 && ~x19 && ~x20 && ~x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x21 && x66 )
						nx_state = s1;
					else if( ~x21 && ~x66 && x22 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x21 && ~x66 && ~x22 )
						nx_state = s1;
					else nx_state = s157;
				s158 : if( x69 && x70 && x63 && x64 )
						begin
							y21 = 1'b1;	y27 = 1'b1;	y48 = 1'b1;	
							nx_state = s877;
						end
					else if( x69 && x70 && x63 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && ~x63 )
						begin
							y47 = 1'b1;	y51 = 1'b1;	y61 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s878;
						end
					else if( x69 && ~x70 && x66 && x65 && x61 && x60 )
						nx_state = s47;
					else if( x69 && ~x70 && x66 && x65 && x61 && ~x60 && x62 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && x61 && ~x60 && ~x62 && x15 && x12 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x69 && ~x70 && x66 && x65 && x61 && ~x60 && ~x62 && x15 && x12 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s609;
						end
					else if( x69 && ~x70 && x66 && x65 && x61 && ~x60 && ~x62 && x15 && ~x12 && x7 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x69 && ~x70 && x66 && x65 && x61 && ~x60 && ~x62 && x15 && ~x12 && ~x7 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s565;
						end
					else if( x69 && ~x70 && x66 && x65 && x61 && ~x60 && ~x62 && ~x15 && x16 && x7 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s811;
						end
					else if( x69 && ~x70 && x66 && x65 && x61 && ~x60 && ~x62 && ~x15 && x16 && x7 && ~x12 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s707;
						end
					else if( x69 && ~x70 && x66 && x65 && x61 && ~x60 && ~x62 && ~x15 && x16 && ~x7 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s707;
						end
					else if( x69 && ~x70 && x66 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x16 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s812;
						end
					else if( x69 && ~x70 && x66 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x16 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x61 && x60 && x15 && x12 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x61 && x60 && x15 && x12 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s609;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x61 && x60 && x15 && ~x12 && x7 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x61 && x60 && x15 && ~x12 && ~x7 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s565;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x61 && x60 && ~x15 && x16 && x7 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s811;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x61 && x60 && ~x15 && x16 && x7 && ~x12 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s707;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x61 && x60 && ~x15 && x16 && ~x7 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s707;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x61 && x60 && ~x15 && ~x16 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s812;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x61 && x60 && ~x15 && ~x16 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x61 && ~x60 && x62 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x61 && ~x60 && ~x62 )
						nx_state = s47;
					else if( x69 && ~x70 && x66 && ~x65 && x67 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && x67 && x62 && ~x61 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && x21 && x68 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && x21 && x68 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && x21 && x68 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && x21 && x68 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && x21 && ~x68 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && x21 && ~x68 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && x21 && ~x68 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && x21 && ~x68 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x22 && x68 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x22 && x68 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x22 && x68 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x7 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x22 && ~x68 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x22 && ~x68 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x22 && ~x68 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x22 && ~x68 && x23 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && x18 && x14 )
						nx_state = s47;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s47;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x22 && ~x68 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x22 && ~x68 && ~x23 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && x26 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && x26 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && x26 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && x26 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && x25 && x26 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && x25 && x26 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && x25 && x26 && x19 && ~x14 && ~x13 )
						nx_state = s158;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && x25 && x26 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && x25 && ~x26 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && x21 && x19 && x17 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s574;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && x21 && x19 && x17 && ~x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s574;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && x21 && x19 && ~x17 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && x21 && x19 && ~x17 && ~x12 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s377;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && x21 && ~x19 && x20 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s574;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && x21 && ~x19 && x20 && ~x12 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s171;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && x21 && ~x19 && ~x20 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s573;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && x21 && ~x19 && ~x20 && ~x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s175;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && x12 && x4 && x18 && x17 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && x12 && x4 && x18 && ~x17 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s576;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && x12 && x4 && ~x18 && x19 && x17 )
						begin
							y18 = 1'b1;	
							nx_state = s574;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && x12 && x4 && ~x18 && x19 && ~x17 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s576;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && x12 && x4 && ~x18 && ~x19 )
						begin
							y18 = 1'b1;	
							nx_state = s574;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && x12 && ~x4 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s576;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && x18 && x4 && x17 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && x18 && x4 && ~x17 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s377;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && x18 && ~x4 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s576;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && x17 && x14 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s576;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && x17 && ~x14 && x16 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s576;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && x17 && ~x14 && ~x16 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && x17 && ~x14 && ~x16 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && x17 && ~x14 && ~x16 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && x17 && ~x14 && ~x16 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && ~x17 && x16 && x15 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s576;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && ~x17 && x16 && ~x15 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && ~x17 && x16 && ~x15 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && ~x17 && x16 && ~x15 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && ~x17 && x16 && ~x15 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && ~x17 && ~x16 && x13 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && ~x17 && ~x16 && x13 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && ~x17 && ~x16 && x13 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && ~x17 && ~x16 && x13 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && ~x17 && ~x16 && ~x13 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s576;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && ~x19 && x4 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && ~x19 && ~x4 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s576;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && x15 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && ~x15 && x19 && x18 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && ~x15 && x19 && ~x18 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && ~x15 && ~x19 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x69 && x44 && x45 && x40 && x24 && x5 && x36 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && x44 && x45 && x40 && x24 && x5 && ~x36 )
						begin
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x69 && x44 && x45 && x40 && x24 && ~x5 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && x44 && x45 && x40 && ~x24 && x31 && x29 )
						begin
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x69 && x44 && x45 && x40 && ~x24 && x31 && ~x29 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && x44 && x45 && x40 && ~x24 && ~x31 )
						begin
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x69 && x44 && x45 && ~x40 && x11 && x35 && x5 )
						begin
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x69 && x44 && x45 && ~x40 && x11 && x35 && ~x5 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && x44 && x45 && ~x40 && x11 && ~x35 && x14 )
						nx_state = s1;
					else if( ~x69 && x44 && x45 && ~x40 && x11 && ~x35 && ~x14 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && x44 && x45 && ~x40 && ~x11 && x30 && x35 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && x44 && x45 && ~x40 && ~x11 && x30 && ~x35 && x14 )
						nx_state = s1;
					else if( ~x69 && x44 && x45 && ~x40 && ~x11 && x30 && ~x35 && ~x14 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && x44 && x45 && ~x40 && ~x11 && ~x30 && x3 && x6 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && x44 && x45 && ~x40 && ~x11 && ~x30 && x3 && ~x6 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && x44 && x45 && ~x40 && ~x11 && ~x30 && ~x3 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && x44 && ~x45 && x46 && x3 )
						nx_state = s1;
					else if( ~x69 && x44 && ~x45 && x46 && ~x3 && x1 )
						begin
							y11 = 1'b1;	
							nx_state = s272;
						end
					else if( ~x69 && x44 && ~x45 && x46 && ~x3 && ~x1 )
						begin
							y8 = 1'b1;	y12 = 1'b1;	
							nx_state = s879;
						end
					else if( ~x69 && x44 && ~x45 && ~x46 && x16 && x14 && x5 )
						begin
							y7 = 1'b1;	
							nx_state = s82;
						end
					else if( ~x69 && x44 && ~x45 && ~x46 && x16 && x14 && ~x5 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && x44 && ~x45 && ~x46 && x16 && ~x14 && x11 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && x44 && ~x45 && ~x46 && x16 && ~x14 && ~x11 && x3 )
						nx_state = s1;
					else if( ~x69 && x44 && ~x45 && ~x46 && x16 && ~x14 && ~x11 && ~x3 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && x44 && ~x45 && ~x46 && ~x16 && x11 && x5 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && x44 && ~x45 && ~x46 && ~x16 && x11 && ~x5 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && x44 && ~x45 && ~x46 && ~x16 && ~x11 && x3 )
						nx_state = s1;
					else if( ~x69 && x44 && ~x45 && ~x46 && ~x16 && ~x11 && ~x3 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x44 && x10 && x11 && x5 && x12 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x44 && x10 && x11 && x5 && ~x12 && x13 )
						begin
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x69 && ~x44 && x10 && x11 && x5 && ~x12 && ~x13 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x69 && ~x44 && x10 && x11 && ~x5 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x44 && x10 && ~x11 && x8 && x1 )
						begin
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x69 && ~x44 && x10 && ~x11 && x8 && ~x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x44 && x10 && ~x11 && ~x8 )
						begin
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x69 && ~x44 && ~x10 && x11 && x13 && x5 )
						begin
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x69 && ~x44 && ~x10 && x11 && x13 && ~x5 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x44 && ~x10 && x11 && ~x13 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x44 && ~x10 && x11 && ~x13 && ~x1 && x3 )
						nx_state = s1;
					else if( ~x69 && ~x44 && ~x10 && x11 && ~x13 && ~x1 && ~x3 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x44 && ~x10 && ~x11 && x12 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x44 && ~x10 && ~x11 && x12 && ~x1 && x3 )
						nx_state = s1;
					else if( ~x69 && ~x44 && ~x10 && ~x11 && x12 && ~x1 && ~x3 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x44 && ~x10 && ~x11 && ~x12 && x3 && x6 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && ~x44 && ~x10 && ~x11 && ~x12 && x3 && ~x6 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x44 && ~x10 && ~x11 && ~x12 && ~x3 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else nx_state = s158;
				s159 : if( 1'b1 )
						begin
							y2 = 1'b1;	y21 = 1'b1;	
							nx_state = s880;
						end
					else nx_state = s159;
				s160 : if( x69 && x70 && x62 && x65 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x69 && x70 && x62 && x65 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x69 && x70 && x62 && x65 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( x69 && x70 && x62 && x65 && ~x27 )
						nx_state = s1;
					else if( x69 && x70 && x62 && ~x65 && x17 && x11 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x69 && x70 && x62 && ~x65 && x17 && x11 && ~x8 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && x70 && x62 && ~x65 && x17 && ~x11 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x17 && x18 && x8 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x17 && x18 && ~x8 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s280;
						end
					else if( x69 && x70 && x62 && ~x65 && ~x17 && ~x18 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && x70 && ~x62 && x63 && x2 && x3 && x11 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( x69 && x70 && ~x62 && x63 && x2 && x3 && ~x11 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s504;
						end
					else if( x69 && x70 && ~x62 && x63 && x2 && ~x3 && x4 && x11 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s670;
						end
					else if( x69 && x70 && ~x62 && x63 && x2 && ~x3 && x4 && ~x11 && x12 && x13 && x14 )
						begin
							y3 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s881;
						end
					else if( x69 && x70 && ~x62 && x63 && x2 && ~x3 && x4 && ~x11 && x12 && x13 && ~x14 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s882;
						end
					else if( x69 && x70 && ~x62 && x63 && x2 && ~x3 && x4 && ~x11 && x12 && ~x13 )
						begin
							y3 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s883;
						end
					else if( x69 && x70 && ~x62 && x63 && x2 && ~x3 && x4 && ~x11 && ~x12 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							y16 = 1'b1;	y21 = 1'b1;	
							nx_state = s884;
						end
					else if( x69 && x70 && ~x62 && x63 && x2 && ~x3 && ~x4 && x6 && x5 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s456;
						end
					else if( x69 && x70 && ~x62 && x63 && x2 && ~x3 && ~x4 && x6 && ~x5 && x9 && x7 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s456;
						end
					else if( x69 && x70 && ~x62 && x63 && x2 && ~x3 && ~x4 && x6 && ~x5 && x9 && ~x7 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && x63 && x2 && ~x3 && ~x4 && x6 && ~x5 && ~x9 && x7 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && x63 && x2 && ~x3 && ~x4 && x6 && ~x5 && ~x9 && ~x7 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s456;
						end
					else if( x69 && x70 && ~x62 && x63 && x2 && ~x3 && ~x4 && ~x6 && x7 && x5 && x8 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s456;
						end
					else if( x69 && x70 && ~x62 && x63 && x2 && ~x3 && ~x4 && ~x6 && x7 && x5 && ~x8 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && x63 && x2 && ~x3 && ~x4 && ~x6 && x7 && ~x5 && x10 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s456;
						end
					else if( x69 && x70 && ~x62 && x63 && x2 && ~x3 && ~x4 && ~x6 && x7 && ~x5 && ~x10 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && x63 && x2 && ~x3 && ~x4 && ~x6 && ~x7 && x5 && x8 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && x63 && x2 && ~x3 && ~x4 && ~x6 && ~x7 && x5 && ~x8 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s456;
						end
					else if( x69 && x70 && ~x62 && x63 && x2 && ~x3 && ~x4 && ~x6 && ~x7 && ~x5 && x10 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && x63 && x2 && ~x3 && ~x4 && ~x6 && ~x7 && ~x5 && ~x10 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s456;
						end
					else if( x69 && x70 && ~x62 && x63 && ~x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x65 && x20 && x3 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x65 && x20 && ~x3 )
						begin
							y11 = 1'b1;	
							nx_state = s91;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x65 && ~x20 && x21 && x3 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x65 && ~x20 && x21 && ~x3 )
						begin
							y31 = 1'b1;	
							nx_state = s886;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x65 && ~x20 && ~x21 && x3 )
						begin
							y14 = 1'b1;	
							nx_state = s5;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x65 && ~x20 && ~x21 && ~x3 )
						begin
							y31 = 1'b1;	
							nx_state = s887;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && x19 && x12 )
						begin
							y54 = 1'b1;	
							nx_state = s525;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && x19 && ~x12 )
						begin
							y55 = 1'b1;	
							nx_state = s526;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && x12 && x6 )
						begin
							y16 = 1'b1;	y50 = 1'b1;	
							nx_state = s527;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && x12 && ~x6 && x16 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && x12 && ~x6 && ~x16 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && x12 && ~x6 && ~x16 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && x12 && ~x6 && ~x16 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && x12 && ~x6 && ~x16 && ~x9 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && ~x12 && x6 )
						begin
							y12 = 1'b1;	y48 = 1'b1;	
							nx_state = s529;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && ~x12 && ~x6 && x15 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && ~x12 && ~x6 && ~x15 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && ~x12 && ~x6 && ~x15 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && ~x12 && ~x6 && ~x15 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && x18 && ~x19 && ~x12 && ~x6 && ~x15 && ~x9 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && ~x18 && x19 )
						begin
							y27 = 1'b1;	y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s284;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && ~x18 && ~x19 && x6 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && x5 && ~x18 && ~x19 && ~x6 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && x19 && x6 && x12 && x11 )
						begin
							y46 = 1'b1;	
							nx_state = s531;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && x19 && x6 && x12 && ~x11 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && x19 && x6 && x12 && ~x11 && x9 && ~x10 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && x19 && x6 && x12 && ~x11 && ~x9 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && x19 && x6 && ~x12 && x10 )
						begin
							y46 = 1'b1;	
							nx_state = s531;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && x19 && x6 && ~x12 && ~x10 && x9 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && x19 && x6 && ~x12 && ~x10 && x9 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && x19 && x6 && ~x12 && ~x10 && ~x9 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && x19 && ~x6 && x12 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && x19 && ~x6 && ~x12 )
						begin
							y56 = 1'b1;	y57 = 1'b1;	
							nx_state = s284;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && x6 && x12 && x14 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && x6 && x12 && ~x14 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && x6 && x12 && ~x14 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && x6 && x12 && ~x14 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && x6 && x12 && ~x14 && ~x9 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && x6 && ~x12 && x13 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && x6 && ~x12 && ~x13 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && x6 && ~x12 && ~x13 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && x6 && ~x12 && ~x13 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && x6 && ~x12 && ~x13 && ~x9 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && x18 && ~x19 && ~x6 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && ~x18 && x19 && x12 && x6 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && ~x18 && x19 && x12 && ~x6 )
						begin
							y38 = 1'b1;	
							nx_state = s532;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && ~x18 && x19 && ~x12 && x6 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && ~x18 && x19 && ~x12 && ~x6 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x65 && ~x5 && ~x18 && ~x19 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 )
						begin
							y37 = 1'b1;	
							nx_state = s888;
						end
					else if( x69 && ~x70 && x65 && x67 && x21 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s889;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x23 && x22 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x23 && x22 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x23 && x22 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x23 && x22 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x23 && ~x22 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x23 && ~x22 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x23 && ~x22 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x21 && x23 && ~x22 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x23 && x8 && x22 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x23 && x8 && x22 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x23 && x8 && x22 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x23 && x8 && ~x22 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x23 && x8 && ~x22 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x23 && x8 && ~x22 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && x67 && ~x21 && ~x23 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && x68 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x68 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && x65 && ~x67 && x68 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && x68 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && x21 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && x23 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && x23 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && x23 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && x23 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && x23 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && x7 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && x7 && ~x9 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && ~x7 && x8 && x9 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s296;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && ~x7 && x8 && ~x9 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s297;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && ~x7 && ~x8 && x9 && x13 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && ~x7 && ~x8 && x9 && ~x13 && x18 && x14 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && ~x7 && ~x8 && x9 && ~x13 && x18 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && ~x7 && ~x8 && x9 && ~x13 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && ~x7 && ~x8 && ~x9 && x14 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && ~x7 && ~x8 && ~x9 && ~x14 && x18 && x13 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && ~x7 && ~x8 && ~x9 && ~x14 && x18 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && ~x7 && ~x8 && ~x9 && ~x14 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && ~x16 && x7 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && ~x16 && ~x7 && x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && ~x16 && ~x7 && ~x8 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && ~x16 && ~x7 && ~x8 && ~x1 && x5 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && ~x16 && ~x7 && ~x8 && ~x1 && ~x5 && x9 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && ~x16 && ~x7 && ~x8 && ~x1 && ~x5 && ~x9 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && x9 && x10 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && x9 && ~x10 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && x9 && ~x10 && ~x8 && x18 && x14 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && x9 && ~x10 && ~x8 && x18 && ~x14 && x13 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && x9 && ~x10 && ~x8 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && x9 && ~x10 && ~x8 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && ~x9 && x8 && x12 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && ~x9 && x8 && ~x12 && x18 && x14 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && ~x9 && x8 && ~x12 && x18 && ~x14 && x13 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && ~x9 && x8 && ~x12 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && ~x9 && x8 && ~x12 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && ~x9 && ~x8 && x11 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && ~x9 && ~x8 && ~x11 && x18 && x14 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && ~x9 && ~x8 && ~x11 && x18 && ~x14 && x13 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && ~x9 && ~x8 && ~x11 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && ~x9 && ~x8 && ~x11 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && ~x16 && x5 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && ~x16 && ~x5 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s495;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && ~x22 && x4 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && ~x22 && x4 && ~x18 && x19 )
						nx_state = s160;
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && ~x22 && x4 && ~x18 && ~x19 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							nx_state = s165;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && ~x22 && ~x4 && x3 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && x65 && ~x67 && ~x68 && ~x21 && ~x22 && ~x4 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x68 && x21 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && x68 && ~x21 && x16 && x10 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x68 && ~x21 && x16 && ~x10 )
						begin
							y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s233;
						end
					else if( x69 && ~x70 && ~x65 && x66 && x68 && ~x21 && ~x16 )
						begin
							y5 = 1'b1;	y17 = 1'b1;	
							nx_state = s721;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && x63 && x64 && x6 && x15 && x8 )
						begin
							y21 = 1'b1;	
							nx_state = s822;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && x63 && x64 && x6 && x15 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && x63 && x64 && x6 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s822;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && x63 && x64 && x6 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s468;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && x63 && x64 && ~x6 )
						begin
							y21 = 1'b1;	
							nx_state = s822;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && x63 && ~x64 && x5 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s102;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && x63 && ~x64 && ~x5 && x18 && x15 && x8 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && x63 && ~x64 && ~x5 && x18 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && x63 && ~x64 && ~x5 && x18 && ~x15 && x16 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && x63 && ~x64 && ~x5 && x18 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s299;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && x63 && ~x64 && ~x5 && ~x18 )
						begin
							y31 = 1'b1;	
							nx_state = s164;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && ~x63 && x64 && x19 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && ~x63 && x64 && x19 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && ~x63 && x64 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && ~x63 && x64 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && ~x63 && ~x64 && x4 )
						begin
							y31 = 1'b1;	
							nx_state = s164;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && ~x63 && ~x64 && ~x4 && x17 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && ~x63 && ~x64 && ~x4 && x17 && x15 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && ~x63 && ~x64 && ~x4 && x17 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && ~x63 && ~x64 && ~x4 && x17 && ~x15 && ~x16 && x14 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s299;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && ~x63 && ~x64 && ~x4 && x17 && ~x15 && ~x16 && ~x14 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s295;
						end
					else if( x69 && ~x70 && ~x65 && x66 && ~x68 && ~x63 && ~x64 && ~x4 && ~x17 )
						begin
							y14 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s100;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && x68 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && x68 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && x68 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && x68 && x20 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && x68 && ~x20 && x21 && x3 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s890;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && x68 && ~x20 && x21 && ~x3 && x17 && x15 && x8 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s242;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && x68 && ~x20 && x21 && ~x3 && x17 && x15 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s556;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && x68 && ~x20 && x21 && ~x3 && x17 && ~x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && x68 && ~x20 && x21 && ~x3 && x17 && ~x15 && ~x16 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s76;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && x68 && ~x20 && x21 && ~x3 && ~x17 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && x68 && ~x20 && ~x21 && x15 && x8 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && x68 && ~x20 && ~x21 && x15 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s556;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && x68 && ~x20 && ~x21 && ~x15 && x16 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s131;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && x68 && ~x20 && ~x21 && ~x15 && ~x16 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s76;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && ~x68 && x24 && x26 && x16 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && ~x68 && x24 && x26 && x16 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && ~x68 && x24 && x26 && x16 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && ~x68 && x24 && x26 && x16 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && ~x68 && x24 && x26 && ~x16 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s304;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && ~x68 && x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && ~x68 && x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && ~x68 && x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && ~x68 && x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && ~x68 && ~x24 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && ~x68 && ~x24 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && ~x68 && ~x24 && x25 && x19 && ~x14 && ~x13 && x26 )
						nx_state = s160;
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && ~x68 && ~x24 && x25 && x19 && ~x14 && ~x13 && ~x26 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && ~x68 && ~x24 && x25 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && ~x68 && ~x24 && ~x25 && x26 )
						begin
							y17 = 1'b1;	
							nx_state = s98;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && ~x68 && ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && ~x68 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && ~x68 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && x67 && ~x68 && ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && x68 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && x68 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && x68 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && x68 && ~x3 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && ~x68 && x21 && x9 && x3 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && ~x68 && x21 && x9 && ~x3 && x4 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && ~x68 && x21 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && ~x68 && x21 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x5 && ~x4 && x22 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x5 && ~x4 && x22 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x5 && ~x4 && ~x22 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x5 && x22 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x5 && ~x22 && x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x5 && ~x22 && x4 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x5 && ~x22 && ~x4 )
						nx_state = s1;
					else if( ~x69 && x70 && x55 && x48 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s456;
						end
					else if( ~x69 && x70 && x55 && ~x48 && x57 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && x70 && x55 && ~x48 && ~x57 )
						nx_state = s160;
					else if( ~x69 && x70 && ~x55 && x37 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s456;
						end
					else if( ~x69 && x70 && ~x55 && ~x37 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x69 && ~x70 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x69 && ~x70 && ~x4 )
						nx_state = s160;
					else nx_state = s160;
				s161 : if( x22 && x20 && x19 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s161;
						end
					else if( x22 && x20 && ~x19 && x23 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x22 && x20 && ~x19 && ~x23 )
						nx_state = s161;
					else if( x22 && ~x20 && x23 && x19 )
						nx_state = s161;
					else if( x22 && ~x20 && x23 && ~x19 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x22 && ~x20 && ~x23 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x22 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else nx_state = s161;
				s162 : if( x70 && x64 && x62 && x66 && x32 )
						begin
							y29 = 1'b1;	
							nx_state = s771;
						end
					else if( x70 && x64 && x62 && x66 && ~x32 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s340;
						end
					else if( x70 && x64 && x62 && ~x66 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x70 && x64 && x62 && ~x66 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x70 && x64 && x62 && ~x66 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x70 && x64 && x62 && ~x66 && ~x19 )
						nx_state = s1;
					else if( x70 && x64 && ~x62 && x63 && x9 )
						begin
							y15 = 1'b1;	
							nx_state = s22;
						end
					else if( x70 && x64 && ~x62 && x63 && ~x9 && x20 )
						begin
							y54 = 1'b1;	
							nx_state = s525;
						end
					else if( x70 && x64 && ~x62 && x63 && ~x9 && ~x20 && x21 )
						begin
							y22 = 1'b1;	
							nx_state = s39;
						end
					else if( x70 && x64 && ~x62 && x63 && ~x9 && ~x20 && ~x21 )
						begin
							y15 = 1'b1;	
							nx_state = s22;
						end
					else if( x70 && x64 && ~x62 && ~x63 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x70 && x64 && ~x62 && ~x63 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x70 && x64 && ~x62 && ~x63 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && x64 && ~x62 && ~x63 && ~x14 )
						nx_state = s1;
					else if( x70 && ~x64 && x62 && x60 )
						begin
							y7 = 1'b1;	
							nx_state = s891;
						end
					else if( x70 && ~x64 && x62 && ~x60 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x70 && ~x64 && x62 && ~x60 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x70 && ~x64 && x62 && ~x60 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( x70 && ~x64 && x62 && ~x60 && ~x27 )
						nx_state = s1;
					else if( x70 && ~x64 && ~x62 && x65 && x63 && x66 && x30 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s892;
						end
					else if( x70 && ~x64 && ~x62 && x65 && x63 && x66 && x30 && ~x4 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x70 && ~x64 && ~x62 && x65 && x63 && x66 && ~x30 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x70 && ~x64 && ~x62 && x65 && x63 && x66 && ~x30 && ~x15 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x64 && ~x62 && x65 && x63 && ~x66 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x70 && ~x64 && ~x62 && x65 && x63 && ~x66 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x70 && ~x64 && ~x62 && x65 && x63 && ~x66 && x19 && ~x14 && ~x13 && x11 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( x70 && ~x64 && ~x62 && x65 && x63 && ~x66 && x19 && ~x14 && ~x13 && x11 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( x70 && ~x64 && ~x62 && x65 && x63 && ~x66 && x19 && ~x14 && ~x13 && ~x11 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( x70 && ~x64 && ~x62 && x65 && x63 && ~x66 && ~x19 )
						nx_state = s1;
					else if( x70 && ~x64 && ~x62 && x65 && ~x63 && x67 && x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x64 && ~x62 && x65 && ~x63 && x67 && x11 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x64 && ~x62 && x65 && ~x63 && x67 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x70 && ~x64 && ~x62 && x65 && ~x63 && x67 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x64 && ~x62 && x65 && ~x63 && ~x67 && x17 )
						begin
							y29 = 1'b1;	
							nx_state = s771;
						end
					else if( x70 && ~x64 && ~x62 && x65 && ~x63 && ~x67 && ~x17 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x64 && ~x62 && x65 && ~x63 && ~x67 && ~x17 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x64 && ~x62 && x65 && ~x63 && ~x67 && ~x17 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x70 && ~x64 && ~x62 && x65 && ~x63 && ~x67 && ~x17 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x64 && ~x62 && ~x65 && x63 && x16 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x64 && ~x62 && ~x65 && x63 && x16 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x64 && ~x62 && ~x65 && x63 && x16 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x70 && ~x64 && ~x62 && ~x65 && x63 && ~x16 )
						nx_state = s1;
					else if( x70 && ~x64 && ~x62 && ~x65 && ~x63 && x66 && x21 && x22 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( x70 && ~x64 && ~x62 && ~x65 && ~x63 && x66 && x21 && ~x22 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( x70 && ~x64 && ~x62 && ~x65 && ~x63 && x66 && x21 && ~x22 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x64 && ~x62 && ~x65 && ~x63 && x66 && ~x21 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( x70 && ~x64 && ~x62 && ~x65 && ~x63 && x66 && ~x21 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x64 && ~x62 && ~x65 && ~x63 && ~x66 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x64 && ~x62 && ~x65 && ~x63 && ~x66 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x64 && ~x62 && ~x65 && ~x63 && ~x66 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x64 && ~x62 && ~x65 && ~x63 && ~x66 && ~x17 )
						nx_state = s1;
					else if( ~x70 && x22 && x4 && x19 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s161;
						end
					else if( ~x70 && x22 && x4 && ~x19 && x20 )
						nx_state = s162;
					else if( ~x70 && x22 && x4 && ~x19 && ~x20 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x70 && x22 && ~x4 && x3 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x70 && x22 && ~x4 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x70 && ~x22 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	y29 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s162;
				s163 : if( x21 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && x18 && x15 && x9 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x21 && x22 && x23 && x18 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x21 && x22 && x23 && x18 && ~x15 && x16 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && x22 && x23 && x18 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s495;
						end
					else if( ~x21 && x22 && x23 && ~x18 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							nx_state = s165;
						end
					else if( ~x21 && x22 && ~x23 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							nx_state = s165;
						end
					else if( ~x21 && ~x22 && x23 && x15 && x9 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x21 && ~x22 && x23 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x21 && ~x22 && x23 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x22 && x23 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s495;
						end
					else if( ~x21 && ~x22 && ~x23 )
						nx_state = s1;
					else nx_state = s163;
				s164 : if( x70 && x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x70 && ~x64 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x70 && ~x64 && ~x8 && x10 && x9 )
						begin
							y27 = 1'b1;	
							nx_state = s893;
						end
					else if( x70 && ~x64 && ~x8 && x10 && ~x9 )
						begin
							y25 = 1'b1;	
							nx_state = s53;
						end
					else if( x70 && ~x64 && ~x8 && ~x10 && x9 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( x70 && ~x64 && ~x8 && ~x10 && ~x9 )
						begin
							y23 = 1'b1;	
							nx_state = s588;
						end
					else if( ~x70 && x65 && x21 && x17 && x15 && x9 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x70 && x65 && x21 && x17 && x15 && ~x9 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && x65 && x21 && x17 && ~x15 && x16 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x70 && x65 && x21 && x17 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s333;
						end
					else if( ~x70 && x65 && x21 && ~x17 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s494;
						end
					else if( ~x70 && x65 && ~x21 && x23 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s494;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && x22 && x5 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s494;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && x22 && ~x5 && x17 && x15 && x9 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && x22 && ~x5 && x17 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && x22 && ~x5 && x17 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && x22 && ~x5 && x17 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s495;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && x22 && ~x5 && ~x17 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && ~x22 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s406;
						end
					else if( ~x70 && ~x65 && x63 )
						begin
							y14 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x70 && ~x65 && ~x63 && x64 && x18 && x16 && x8 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x65 && ~x63 && x64 && x18 && x16 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && ~x65 && ~x63 && x64 && x18 && ~x16 && x4 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x70 && ~x65 && ~x63 && x64 && x18 && ~x16 && ~x4 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s299;
						end
					else if( ~x70 && ~x65 && ~x63 && x64 && ~x18 )
						begin
							y14 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x70 && ~x65 && ~x63 && ~x64 && x17 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x70 && ~x65 && ~x63 && ~x64 && x17 && x15 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && ~x65 && ~x63 && ~x64 && x17 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( ~x70 && ~x65 && ~x63 && ~x64 && x17 && ~x15 && ~x16 && x14 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s299;
						end
					else if( ~x70 && ~x65 && ~x63 && ~x64 && x17 && ~x15 && ~x16 && ~x14 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s295;
						end
					else if( ~x70 && ~x65 && ~x63 && ~x64 && ~x17 )
						begin
							y14 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s100;
						end
					else nx_state = s164;
				s165 : if( x23 && x22 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s166;
						end
					else if( x23 && ~x22 )
						nx_state = s1;
					else if( ~x23 && x22 )
						begin
							y21 = 1'b1;	
							nx_state = s822;
						end
					else if( ~x23 && ~x22 && x4 && x20 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x23 && ~x22 && x4 && ~x20 && x19 )
						nx_state = s165;
					else if( ~x23 && ~x22 && x4 && ~x20 && ~x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( ~x23 && ~x22 && ~x4 && x3 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s161;
						end
					else if( ~x23 && ~x22 && ~x4 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else nx_state = s165;
				s166 : if( x22 && x15 && x9 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x22 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x22 && ~x15 && x16 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x22 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s495;
						end
					else if( ~x22 && x19 && x20 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x22 && x19 && ~x20 )
						nx_state = s166;
					else if( ~x22 && ~x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else nx_state = s166;
				s167 : if( x23 && x22 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x23 && x22 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x23 && x22 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x23 && x22 && ~x17 )
						nx_state = s1;
					else if( x23 && ~x22 )
						nx_state = s1;
					else if( ~x23 )
						nx_state = s1;
					else nx_state = s167;
				s168 : if( x65 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x5 )
						nx_state = s1;
					else if( ~x65 && x21 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x16 && x12 && x19 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x16 && x12 && ~x19 && x18 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x65 && ~x21 && x22 && x16 && x12 && ~x19 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x16 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x16 )
						nx_state = s1;
					else if( ~x65 && ~x21 && ~x22 && x18 && x15 )
						begin
							y8 = 1'b1;	y18 = 1'b1;	
							nx_state = s152;
						end
					else if( ~x65 && ~x21 && ~x22 && x18 && ~x15 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s6;
						end
					else if( ~x65 && ~x21 && ~x22 && ~x18 && x19 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s835;
						end
					else if( ~x65 && ~x21 && ~x22 && ~x18 && x19 && ~x15 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && ~x21 && ~x22 && ~x18 && ~x19 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else nx_state = s168;
				s169 : if( x21 && x12 && x11 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x21 && x12 && ~x11 && x10 )
						nx_state = s169;
					else if( x21 && x12 && ~x11 && ~x10 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s170;
						end
					else if( x21 && ~x12 && x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x21 && ~x12 && ~x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x21 && x22 && x19 && x15 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y17 = 1'b1;	
							nx_state = s314;
						end
					else if( ~x21 && x22 && x19 && ~x15 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							nx_state = s315;
						end
					else if( ~x21 && x22 && ~x19 && x20 && x14 && x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s316;
						end
					else if( ~x21 && x22 && ~x19 && x20 && x14 && ~x18 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && ~x19 && x20 && x14 && ~x18 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && ~x19 && x20 && x14 && ~x18 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x20 && x14 && ~x18 && ~x5 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x20 && ~x14 && x15 && x16 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s316;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x14 && x15 && ~x16 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x14 && x15 && ~x16 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x14 && x15 && ~x16 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x20 && ~x14 && x15 && ~x16 && ~x5 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x20 && ~x14 && ~x15 && x17 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s316;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x14 && ~x15 && ~x17 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x14 && ~x15 && ~x17 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x14 && ~x15 && ~x17 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x20 && ~x14 && ~x15 && ~x17 && ~x5 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && ~x20 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( ~x21 && ~x22 && x7 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( ~x21 && ~x22 && ~x7 && x10 && x19 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && ~x22 && ~x7 && x10 && x19 && ~x15 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	
							nx_state = s315;
						end
					else if( ~x21 && ~x22 && ~x7 && x10 && ~x19 && x20 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( ~x21 && ~x22 && ~x7 && x10 && ~x19 && ~x20 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( ~x21 && ~x22 && ~x7 && ~x10 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s170;
						end
					else nx_state = s169;
				s170 : if( x21 )
						nx_state = s1;
					else if( ~x21 && x22 && x19 && x15 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y17 = 1'b1;	
							nx_state = s314;
						end
					else if( ~x21 && x22 && x19 && ~x15 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							nx_state = s315;
						end
					else if( ~x21 && x22 && ~x19 && x20 && x15 && x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s316;
						end
					else if( ~x21 && x22 && ~x19 && x20 && x15 && ~x14 && x16 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s316;
						end
					else if( ~x21 && x22 && ~x19 && x20 && x15 && ~x14 && ~x16 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && ~x19 && x20 && x15 && ~x14 && ~x16 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && ~x19 && x20 && x15 && ~x14 && ~x16 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x20 && x15 && ~x14 && ~x16 && ~x5 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x20 && ~x15 && x14 && x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s316;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x15 && x14 && ~x18 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x15 && x14 && ~x18 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x15 && x14 && ~x18 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x20 && ~x15 && x14 && ~x18 && ~x5 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x20 && ~x15 && ~x14 && x17 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s316;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && ~x5 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && ~x20 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( ~x21 && ~x22 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s313;
						end
					else nx_state = s170;
				s171 : if( x21 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x21 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x21 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x21 && ~x3 )
						nx_state = s1;
					else if( ~x21 && x22 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s894;
						end
					else if( ~x21 && ~x22 && x18 && x15 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s894;
						end
					else if( ~x21 && ~x22 && x18 && ~x15 && x4 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s377;
						end
					else if( ~x21 && ~x22 && x18 && ~x15 && ~x4 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s894;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && x15 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s894;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && x17 && x13 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s894;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && x17 && ~x13 && x16 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s894;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && x17 && ~x13 && ~x16 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && x17 && ~x13 && ~x16 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && x17 && ~x13 && ~x16 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && x17 && ~x13 && ~x16 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && ~x17 && x16 && x14 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s894;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && ~x17 && x16 && ~x14 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && ~x17 && x16 && ~x14 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && ~x17 && x16 && ~x14 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && ~x17 && x16 && ~x14 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && x12 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s894;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && ~x12 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && ~x12 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && ~x12 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && ~x12 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x18 && ~x19 && x4 )
						begin
							y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s378;
						end
					else if( ~x21 && ~x22 && ~x18 && ~x19 && ~x4 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s894;
						end
					else nx_state = s171;
				s172 : if( x21 && x8 && x19 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x21 && x8 && ~x19 && x20 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s313;
						end
					else if( x21 && x8 && ~x19 && ~x20 )
						begin
							y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s386;
						end
					else if( x21 && ~x8 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	
							nx_state = s895;
						end
					else if( ~x21 && x22 && x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y9 = 1'b1;	
							nx_state = s173;
						end
					else if( ~x21 && x22 && x11 && ~x2 )
						nx_state = s47;
					else if( ~x21 && x22 && ~x11 && x9 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x21 && x22 && ~x11 && ~x9 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x21 && ~x22 )
						nx_state = s1;
					else nx_state = s172;
				s173 : if( x21 && x19 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x21 && ~x19 )
						begin
							y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s386;
						end
					else if( ~x21 && x22 && x3 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y9 = 1'b1;	
							nx_state = s173;
						end
					else if( ~x21 && x22 && x3 && ~x2 )
						nx_state = s47;
					else if( ~x21 && x22 && ~x3 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( ~x21 && ~x22 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s438;
						end
					else nx_state = s173;
				s174 : if( x21 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s896;
						end
					else if( ~x21 && x22 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x22 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y9 = 1'b1;	
							nx_state = s173;
						end
					else nx_state = s174;
				s175 : if( x21 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( ~x21 && x22 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x21 && x22 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x21 && x22 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 )
						nx_state = s1;
					else nx_state = s175;
				s176 : if( x70 )
						begin
							y13 = 1'b1;	
							nx_state = s897;
						end
					else if( ~x70 && x45 && x12 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && x45 && ~x12 && x6 && x2 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s578;
						end
					else if( ~x70 && x45 && ~x12 && x6 && ~x2 )
						nx_state = s176;
					else if( ~x70 && x45 && ~x12 && ~x6 && x2 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && x45 && ~x12 && ~x6 && ~x2 )
						nx_state = s176;
					else if( ~x70 && ~x45 && x46 && x6 && x2 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s578;
						end
					else if( ~x70 && ~x45 && x46 && x6 && ~x2 )
						nx_state = s176;
					else if( ~x70 && ~x45 && x46 && ~x6 && x2 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && ~x45 && x46 && ~x6 && ~x2 )
						nx_state = s176;
					else if( ~x70 && ~x45 && ~x46 && x10 && x6 && x2 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s578;
						end
					else if( ~x70 && ~x45 && ~x46 && x10 && x6 && ~x2 )
						nx_state = s176;
					else if( ~x70 && ~x45 && ~x46 && x10 && ~x6 && x2 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && ~x45 && ~x46 && x10 && ~x6 && ~x2 )
						nx_state = s176;
					else if( ~x70 && ~x45 && ~x46 && ~x10 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else nx_state = s176;
				s177 : if( x70 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x70 && ~x1 && x2 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( x70 && ~x1 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && x45 && x12 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x70 && x45 && x12 && ~x1 && x2 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x45 && x12 && ~x1 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && x45 && ~x12 && x6 && x2 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s578;
						end
					else if( ~x70 && x45 && ~x12 && x6 && ~x2 )
						nx_state = s177;
					else if( ~x70 && x45 && ~x12 && ~x6 && x2 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && x45 && ~x12 && ~x6 && ~x2 )
						nx_state = s177;
					else if( ~x70 && ~x45 && x46 && x6 && x2 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s578;
						end
					else if( ~x70 && ~x45 && x46 && x6 && ~x2 )
						nx_state = s177;
					else if( ~x70 && ~x45 && x46 && ~x6 && x2 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && ~x45 && x46 && ~x6 && ~x2 )
						nx_state = s177;
					else if( ~x70 && ~x45 && ~x46 && x10 && x6 && x2 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s578;
						end
					else if( ~x70 && ~x45 && ~x46 && x10 && x6 && ~x2 )
						nx_state = s177;
					else if( ~x70 && ~x45 && ~x46 && x10 && ~x6 && x2 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && ~x45 && ~x46 && x10 && ~x6 && ~x2 )
						nx_state = s177;
					else if( ~x70 && ~x45 && ~x46 && ~x10 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x70 && ~x45 && ~x46 && ~x10 && ~x1 && x2 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x45 && ~x46 && ~x10 && ~x1 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else nx_state = s177;
				s178 : if( x69 && x65 && x66 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && x66 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && x66 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && x65 && x66 && x20 && ~x17 )
						nx_state = s1;
					else if( x69 && x65 && x66 && ~x20 && x15 && x10 && x11 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s600;
						end
					else if( x69 && x65 && x66 && ~x20 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s601;
						end
					else if( x69 && x65 && x66 && ~x20 && x15 && x10 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y13 = 1'b1;	
							nx_state = s600;
						end
					else if( x69 && x65 && x66 && ~x20 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( x69 && x65 && x66 && ~x20 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s602;
						end
					else if( x69 && x65 && x66 && ~x20 && ~x15 && x16 && x10 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s825;
						end
					else if( x69 && x65 && x66 && ~x20 && ~x15 && x16 && ~x10 && x12 && x11 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( x69 && x65 && x66 && ~x20 && ~x15 && x16 && ~x10 && x12 && ~x11 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s825;
						end
					else if( x69 && x65 && x66 && ~x20 && ~x15 && x16 && ~x10 && ~x12 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s825;
						end
					else if( x69 && x65 && x66 && ~x20 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s604;
						end
					else if( x69 && x65 && ~x66 && x21 && x68 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x69 && x65 && ~x66 && x21 && ~x68 && x7 && x16 && x13 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && x21 && ~x68 && x7 && x16 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s252;
						end
					else if( x69 && x65 && ~x66 && x21 && ~x68 && x7 && ~x16 && x17 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && x21 && ~x68 && x7 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s252;
						end
					else if( x69 && x65 && ~x66 && x21 && ~x68 && ~x7 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && x68 && x8 && x23 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && x68 && x8 && x23 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && x68 && x8 && x23 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && x22 && x68 && x8 && ~x23 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && x68 && x8 && ~x23 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && x68 && x8 && ~x23 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && x22 && x68 && ~x8 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && x16 && x18 && x19 && x10 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && x16 && x18 && x19 && ~x10 && x7 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && x16 && x18 && x19 && ~x10 && ~x7 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && x16 && x18 && ~x19 && x7 && x13 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && x16 && x18 && ~x19 && x7 && ~x13 )
						begin
							y26 = 1'b1;	
							nx_state = s262;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && x16 && x18 && ~x19 && ~x7 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && x16 && ~x18 && x13 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && x16 && ~x18 && ~x13 && x7 && x19 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s264;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && x16 && ~x18 && ~x13 && x7 && ~x19 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s252;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && x16 && ~x18 && ~x13 && ~x7 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && x10 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && x15 && x12 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && x15 && ~x12 && x14 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && x15 && ~x12 && ~x14 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && x15 && ~x12 && ~x14 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && x15 && ~x12 && ~x14 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && x15 && ~x12 && ~x14 && ~x4 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && ~x15 && x14 && x13 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && ~x15 && x14 && ~x13 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && ~x15 && x14 && ~x13 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && ~x15 && x14 && ~x13 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && ~x15 && x14 && ~x13 && ~x4 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && ~x15 && ~x14 && x11 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && ~x15 && ~x14 && ~x11 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && ~x15 && ~x14 && ~x11 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && ~x15 && ~x14 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && ~x15 && ~x14 && ~x11 && ~x4 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && ~x19 && x7 && x13 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && ~x19 && x7 && ~x13 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && ~x19 && ~x7 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && x13 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && x15 && x11 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && x15 && ~x11 && x14 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && x15 && ~x11 && ~x14 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && x15 && ~x11 && ~x14 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && x15 && ~x11 && ~x14 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && x15 && ~x11 && ~x14 && ~x4 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && x14 && x12 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && x14 && ~x12 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && x14 && ~x12 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && x14 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && x14 && ~x12 && ~x4 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && ~x14 && x10 && x19 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && ~x14 && x10 && ~x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && ~x14 && x10 && ~x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && ~x14 && x10 && ~x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && ~x14 && x10 && ~x19 && ~x4 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && ~x14 && ~x10 && x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && ~x14 && ~x10 && x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && ~x14 && ~x10 && x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && ~x14 && ~x10 && x19 && ~x4 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && ~x14 && ~x10 && ~x19 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && ~x17 && x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s252;
						end
					else if( x69 && x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && ~x17 && ~x7 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && x68 && x23 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && x68 && x23 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && x68 && x23 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && x68 && x23 && ~x9 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && x68 && ~x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && x68 && ~x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && x68 && ~x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && x68 && ~x23 && ~x8 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && x17 && x13 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && x17 && ~x13 && x7 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s264;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && x17 && ~x13 && ~x7 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && x13 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && x15 && x11 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && x15 && ~x11 && x14 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && x15 && ~x11 && ~x14 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && x15 && ~x11 && ~x14 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && x15 && ~x11 && ~x14 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && x15 && ~x11 && ~x14 && ~x4 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && ~x15 && x14 && x12 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && ~x15 && x14 && ~x12 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && ~x15 && x14 && ~x12 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && ~x15 && x14 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && ~x15 && x14 && ~x12 && ~x4 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && ~x15 && ~x14 && x10 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && ~x15 && ~x14 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && ~x15 && ~x14 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && ~x15 && ~x14 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && ~x15 && ~x14 && ~x10 && ~x4 )
						nx_state = s1;
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && ~x18 && x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s252;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && ~x18 && ~x7 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && ~x19 && x16 && x13 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && ~x19 && x16 && ~x13 && x7 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s252;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && ~x19 && x16 && ~x13 && ~x7 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && ~x19 && ~x16 && x17 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && ~x19 && ~x16 && ~x17 && x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s252;
						end
					else if( x69 && x65 && ~x66 && ~x21 && ~x22 && ~x68 && ~x19 && ~x16 && ~x17 && ~x7 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s898;
						end
					else if( x69 && ~x65 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x65 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x65 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x65 && x20 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x20 && x21 && x15 && x16 && x14 && x8 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s358;
						end
					else if( x69 && ~x65 && ~x20 && x21 && x15 && x16 && x14 && ~x8 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	y20 = 1'b1;	
							nx_state = s781;
						end
					else if( x69 && ~x65 && ~x20 && x21 && x15 && x16 && ~x14 && x7 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else if( x69 && ~x65 && ~x20 && x21 && x15 && x16 && ~x14 && x7 && ~x8 )
						begin
							y7 = 1'b1;	y12 = 1'b1;	
							nx_state = s610;
						end
					else if( x69 && ~x65 && ~x20 && x21 && x15 && x16 && ~x14 && ~x7 && x8 && x12 )
						begin
							y17 = 1'b1;	
							nx_state = s3;
						end
					else if( x69 && ~x65 && ~x20 && x21 && x15 && x16 && ~x14 && ~x7 && x8 && ~x12 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && ~x65 && ~x20 && x21 && x15 && x16 && ~x14 && ~x7 && x8 && ~x12 && x18 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x20 && x21 && x15 && x16 && ~x14 && ~x7 && x8 && ~x12 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x20 && x21 && x15 && x16 && ~x14 && ~x7 && ~x8 && x13 )
						begin
							y17 = 1'b1;	
							nx_state = s3;
						end
					else if( x69 && ~x65 && ~x20 && x21 && x15 && x16 && ~x14 && ~x7 && ~x8 && ~x13 && x18 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && ~x65 && ~x20 && x21 && x15 && x16 && ~x14 && ~x7 && ~x8 && ~x13 && x18 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x20 && x21 && x15 && x16 && ~x14 && ~x7 && ~x8 && ~x13 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x20 && x21 && x15 && ~x16 && x7 && x8 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( x69 && ~x65 && ~x20 && x21 && x15 && ~x16 && x7 && ~x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x65 && ~x20 && x21 && x15 && ~x16 && ~x7 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s899;
						end
					else if( x69 && ~x65 && ~x20 && x21 && x15 && ~x16 && ~x7 && ~x2 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x69 && ~x65 && ~x20 && x21 && x15 && ~x16 && ~x7 && ~x2 && ~x3 && x8 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x65 && ~x20 && x21 && x15 && ~x16 && ~x7 && ~x2 && ~x3 && ~x8 )
						begin
							y2 = 1'b1;	y13 = 1'b1;	
							nx_state = s780;
						end
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s899;
						end
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && x7 && x11 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && x7 && x11 && ~x3 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && x7 && ~x11 && x8 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && x7 && ~x11 && x8 && ~x3 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && x7 && ~x11 && ~x8 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && x7 && ~x11 && ~x8 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && x7 && ~x11 && ~x8 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && x7 && ~x11 && ~x8 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && x8 && x9 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && x8 && x9 && ~x3 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && x8 && ~x9 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && x8 && ~x9 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && x8 && ~x9 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && x8 && ~x9 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && x10 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && x10 && ~x3 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && ~x10 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && ~x10 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && ~x10 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && ~x10 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && ~x16 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x69 && ~x65 && ~x20 && x21 && ~x15 && ~x2 && ~x16 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s668;
						end
					else if( x69 && ~x65 && ~x20 && ~x21 && x6 && x15 && x8 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s890;
						end
					else if( x69 && ~x65 && ~x20 && ~x21 && x6 && x15 && ~x8 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s781;
						end
					else if( x69 && ~x65 && ~x20 && ~x21 && x6 && ~x15 && x16 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s890;
						end
					else if( x69 && ~x65 && ~x20 && ~x21 && x6 && ~x15 && ~x16 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s668;
						end
					else if( x69 && ~x65 && ~x20 && ~x21 && ~x6 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s890;
						end
					else if( ~x69 && x70 && x10 && x8 && x1 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x69 && x70 && x10 && x8 && ~x1 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s209;
						end
					else if( ~x69 && x70 && x10 && ~x8 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x69 && x70 && ~x10 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( ~x69 && x70 && ~x10 && ~x1 && x3 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x10 && ~x1 && ~x3 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s209;
						end
					else if( ~x69 && ~x70 && x3 && x5 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x70 && x3 && ~x5 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s209;
						end
					else if( ~x69 && ~x70 && ~x3 && x1 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x70 && ~x3 && ~x1 && x8 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s209;
						end
					else if( ~x69 && ~x70 && ~x3 && ~x1 && ~x8 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else nx_state = s178;
				s179 : if( x42 && x43 && x10 && x34 && x44 && x4 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( x42 && x43 && x10 && x34 && x44 && ~x4 )
						nx_state = s179;
					else if( x42 && x43 && x10 && x34 && ~x44 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x42 && x43 && x10 && x34 && ~x44 && ~x4 )
						nx_state = s179;
					else if( x42 && x43 && x10 && ~x34 && x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x42 && x43 && x10 && ~x34 && ~x4 )
						nx_state = s179;
					else if( x42 && x43 && ~x10 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s99;
						end
					else if( x42 && ~x43 && x13 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s99;
						end
					else if( x42 && ~x43 && ~x13 && x41 && x14 && x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x42 && ~x43 && ~x13 && x41 && x14 && ~x4 )
						nx_state = s179;
					else if( x42 && ~x43 && ~x13 && x41 && ~x14 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( x42 && ~x43 && ~x13 && x41 && ~x14 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( x42 && ~x43 && ~x13 && x41 && ~x14 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( x42 && ~x43 && ~x13 && x41 && ~x14 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x42 && ~x43 && ~x13 && x41 && ~x14 && x15 && ~x47 && ~x1 )
						nx_state = s179;
					else if( x42 && ~x43 && ~x13 && x41 && ~x14 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x42 && ~x43 && ~x13 && x41 && ~x14 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x42 && ~x43 && ~x13 && x41 && ~x14 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x42 && ~x43 && ~x13 && ~x41 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s99;
						end
					else if( ~x42 && x10 && x12 && x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x42 && x10 && x12 && ~x4 )
						nx_state = s179;
					else if( ~x42 && x10 && ~x12 && x44 && x45 && x35 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x42 && x10 && ~x12 && x44 && x45 && x35 && ~x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x42 && x10 && ~x12 && x44 && x45 && ~x35 )
						nx_state = s179;
					else if( ~x42 && x10 && ~x12 && x44 && ~x45 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x42 && x10 && ~x12 && x44 && ~x45 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x42 && x10 && ~x12 && x44 && ~x45 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x42 && x10 && ~x12 && x44 && ~x45 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && x10 && ~x12 && x44 && ~x45 && x15 && ~x47 && ~x1 )
						nx_state = s179;
					else if( ~x42 && x10 && ~x12 && x44 && ~x45 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && x10 && ~x12 && x44 && ~x45 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x42 && x10 && ~x12 && x44 && ~x45 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && x10 && ~x12 && ~x44 && x14 && x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x42 && x10 && ~x12 && ~x44 && x14 && ~x4 )
						nx_state = s179;
					else if( ~x42 && x10 && ~x12 && ~x44 && ~x14 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x42 && x10 && ~x12 && ~x44 && ~x14 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x42 && x10 && ~x12 && ~x44 && ~x14 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x42 && x10 && ~x12 && ~x44 && ~x14 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && x10 && ~x12 && ~x44 && ~x14 && x15 && ~x47 && ~x1 )
						nx_state = s179;
					else if( ~x42 && x10 && ~x12 && ~x44 && ~x14 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && x10 && ~x12 && ~x44 && ~x14 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x42 && x10 && ~x12 && ~x44 && ~x14 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && ~x10 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s99;
						end
					else nx_state = s179;
				s180 : if( x62 && x16 && x15 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x62 && x16 && ~x15 && x4 && x5 && x1 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s900;
						end
					else if( x62 && x16 && ~x15 && x4 && x5 && ~x1 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s194;
						end
					else if( x62 && x16 && ~x15 && x4 && ~x5 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s901;
						end
					else if( x62 && x16 && ~x15 && x4 && ~x5 && ~x1 )
						begin
							y10 = 1'b1;	
							nx_state = s193;
						end
					else if( x62 && x16 && ~x15 && ~x4 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x62 && ~x16 && x15 && x3 && x2 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s451;
						end
					else if( x62 && ~x16 && x15 && x3 && ~x2 )
						nx_state = s180;
					else if( x62 && ~x16 && x15 && ~x3 && x4 && x2 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s194;
						end
					else if( x62 && ~x16 && x15 && ~x3 && x4 && ~x2 )
						nx_state = s180;
					else if( x62 && ~x16 && x15 && ~x3 && ~x4 && x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x62 && ~x16 && x15 && ~x3 && ~x4 && ~x2 )
						nx_state = s180;
					else if( x62 && ~x16 && ~x15 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s900;
						end
					else if( ~x62 && x42 && x43 && x44 && x10 && x33 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x62 && x42 && x43 && x44 && x10 && ~x33 )
						nx_state = s180;
					else if( ~x62 && x42 && x43 && x44 && ~x10 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x62 && x42 && x43 && ~x44 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x62 && x42 && ~x43 && x13 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x62 && x42 && ~x43 && ~x13 && x41 && x2 && x45 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x62 && x42 && ~x43 && ~x13 && x41 && x2 && ~x45 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x62 && x42 && ~x43 && ~x13 && x41 && ~x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x62 && x42 && ~x43 && ~x13 && ~x41 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x62 && ~x42 && x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x62 && ~x42 && ~x12 && x44 && x14 && x10 && x33 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x62 && ~x42 && ~x12 && x44 && x14 && x10 && ~x33 )
						nx_state = s180;
					else if( ~x62 && ~x42 && ~x12 && x44 && x14 && ~x10 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x62 && ~x42 && ~x12 && x44 && ~x14 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x62 && ~x42 && ~x12 && ~x44 && x41 && x2 && x45 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x62 && ~x42 && ~x12 && ~x44 && x41 && x2 && ~x45 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x62 && ~x42 && ~x12 && ~x44 && x41 && ~x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x62 && ~x42 && ~x12 && ~x44 && ~x41 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else nx_state = s180;
				s181 : if( x69 && x21 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x69 && ~x21 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s827;
						end
					else if( ~x69 && x11 && x12 && x33 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s801;
						end
					else if( ~x69 && x11 && x12 && ~x33 )
						nx_state = s181;
					else if( ~x69 && x11 && ~x12 && x3 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x11 && ~x12 && x3 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x69 && x11 && ~x12 && x3 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x69 && x11 && ~x12 && x3 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x11 && ~x12 && x3 && x15 && ~x47 && ~x1 )
						nx_state = s181;
					else if( ~x69 && x11 && ~x12 && x3 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x11 && ~x12 && x3 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x69 && x11 && ~x12 && x3 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x11 && ~x12 && ~x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && ~x11 && x3 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && ~x11 && x3 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x69 && ~x11 && x3 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x69 && ~x11 && x3 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && ~x11 && x3 && x15 && ~x47 && ~x1 )
						nx_state = s181;
					else if( ~x69 && ~x11 && x3 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && ~x11 && x3 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x69 && ~x11 && x3 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && ~x11 && ~x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else nx_state = s181;
				s182 : if( x69 && x62 && x13 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s45;
						end
					else if( x69 && x62 && ~x13 && x10 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s551;
						end
					else if( x69 && x62 && ~x13 && x10 && ~x5 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s542;
						end
					else if( x69 && x62 && ~x13 && ~x10 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && ~x62 && x17 && x11 && x8 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && ~x62 && x17 && x11 && ~x8 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && x17 && ~x11 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && ~x17 && x18 && x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s551;
						end
					else if( x69 && ~x62 && ~x17 && x18 && ~x8 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s542;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x69 && x63 && x11 && x43 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s902;
						end
					else if( ~x69 && x63 && x11 && ~x43 && x13 && x7 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x63 && x11 && ~x43 && x13 && x7 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x69 && x63 && x11 && ~x43 && x13 && x7 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x69 && x63 && x11 && ~x43 && x13 && x7 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x63 && x11 && ~x43 && x13 && x7 && x15 && ~x47 && ~x1 )
						nx_state = s182;
					else if( ~x69 && x63 && x11 && ~x43 && x13 && x7 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x63 && x11 && ~x43 && x13 && x7 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x69 && x63 && x11 && ~x43 && x13 && x7 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x63 && x11 && ~x43 && x13 && ~x7 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s902;
						end
					else if( ~x69 && x63 && x11 && ~x43 && ~x13 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s902;
						end
					else if( ~x69 && x63 && ~x11 && x12 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s902;
						end
					else if( ~x69 && x63 && ~x11 && ~x12 && x45 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s902;
						end
					else if( ~x69 && x63 && ~x11 && ~x12 && ~x45 && x7 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x63 && ~x11 && ~x12 && ~x45 && x7 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x69 && x63 && ~x11 && ~x12 && ~x45 && x7 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x69 && x63 && ~x11 && ~x12 && ~x45 && x7 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x63 && ~x11 && ~x12 && ~x45 && x7 && x15 && ~x47 && ~x1 )
						nx_state = s182;
					else if( ~x69 && x63 && ~x11 && ~x12 && ~x45 && x7 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x63 && ~x11 && ~x12 && ~x45 && x7 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x69 && x63 && ~x11 && ~x12 && ~x45 && x7 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x63 && ~x11 && ~x12 && ~x45 && ~x7 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s902;
						end
					else if( ~x69 && ~x63 && x17 && x8 && x11 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( ~x69 && ~x63 && x17 && x8 && ~x11 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && ~x63 && x17 && ~x8 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && ~x63 && ~x17 && x18 && x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s551;
						end
					else if( ~x69 && ~x63 && ~x17 && x18 && ~x8 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s542;
						end
					else if( ~x69 && ~x63 && ~x17 && ~x18 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s543;
						end
					else nx_state = s182;
				s183 : if( x42 && x43 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x42 && x43 && ~x3 && x2 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( x42 && x43 && ~x3 && x2 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( x42 && x43 && ~x3 && x2 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( x42 && x43 && ~x3 && x2 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x42 && x43 && ~x3 && x2 && x15 && ~x47 && ~x1 )
						nx_state = s183;
					else if( x42 && x43 && ~x3 && x2 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x42 && x43 && ~x3 && x2 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x42 && x43 && ~x3 && x2 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x42 && x43 && ~x3 && ~x2 )
						nx_state = s183;
					else if( x42 && ~x43 && x13 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x42 && ~x43 && x13 && ~x3 && x2 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( x42 && ~x43 && x13 && ~x3 && x2 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( x42 && ~x43 && x13 && ~x3 && x2 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( x42 && ~x43 && x13 && ~x3 && x2 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x42 && ~x43 && x13 && ~x3 && x2 && x15 && ~x47 && ~x1 )
						nx_state = s183;
					else if( x42 && ~x43 && x13 && ~x3 && x2 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x42 && ~x43 && x13 && ~x3 && x2 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x42 && ~x43 && x13 && ~x3 && x2 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x42 && ~x43 && x13 && ~x3 && ~x2 )
						nx_state = s183;
					else if( x42 && ~x43 && ~x13 && x45 && x41 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s902;
						end
					else if( x42 && ~x43 && ~x13 && x45 && ~x41 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x42 && ~x43 && ~x13 && x45 && ~x41 && ~x3 && x2 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( x42 && ~x43 && ~x13 && x45 && ~x41 && ~x3 && x2 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( x42 && ~x43 && ~x13 && x45 && ~x41 && ~x3 && x2 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( x42 && ~x43 && ~x13 && x45 && ~x41 && ~x3 && x2 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x42 && ~x43 && ~x13 && x45 && ~x41 && ~x3 && x2 && x15 && ~x47 && ~x1 )
						nx_state = s183;
					else if( x42 && ~x43 && ~x13 && x45 && ~x41 && ~x3 && x2 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x42 && ~x43 && ~x13 && x45 && ~x41 && ~x3 && x2 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x42 && ~x43 && ~x13 && x45 && ~x41 && ~x3 && x2 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x42 && ~x43 && ~x13 && x45 && ~x41 && ~x3 && ~x2 )
						nx_state = s183;
					else if( x42 && ~x43 && ~x13 && ~x45 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x42 && ~x43 && ~x13 && ~x45 && ~x3 && x2 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( x42 && ~x43 && ~x13 && ~x45 && ~x3 && x2 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( x42 && ~x43 && ~x13 && ~x45 && ~x3 && x2 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( x42 && ~x43 && ~x13 && ~x45 && ~x3 && x2 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x42 && ~x43 && ~x13 && ~x45 && ~x3 && x2 && x15 && ~x47 && ~x1 )
						nx_state = s183;
					else if( x42 && ~x43 && ~x13 && ~x45 && ~x3 && x2 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x42 && ~x43 && ~x13 && ~x45 && ~x3 && x2 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x42 && ~x43 && ~x13 && ~x45 && ~x3 && x2 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x42 && ~x43 && ~x13 && ~x45 && ~x3 && ~x2 )
						nx_state = s183;
					else if( ~x42 && x12 && x41 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s902;
						end
					else if( ~x42 && x12 && ~x41 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x42 && x12 && ~x41 && ~x3 && x2 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x42 && x12 && ~x41 && ~x3 && x2 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x42 && x12 && ~x41 && ~x3 && x2 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x42 && x12 && ~x41 && ~x3 && x2 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && x12 && ~x41 && ~x3 && x2 && x15 && ~x47 && ~x1 )
						nx_state = s183;
					else if( ~x42 && x12 && ~x41 && ~x3 && x2 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && x12 && ~x41 && ~x3 && x2 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x42 && x12 && ~x41 && ~x3 && x2 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && x12 && ~x41 && ~x3 && ~x2 )
						nx_state = s183;
					else if( ~x42 && ~x12 && x44 && x14 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x42 && ~x12 && x44 && x14 && ~x3 && x2 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x42 && ~x12 && x44 && x14 && ~x3 && x2 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x42 && ~x12 && x44 && x14 && ~x3 && x2 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x42 && ~x12 && x44 && x14 && ~x3 && x2 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && ~x12 && x44 && x14 && ~x3 && x2 && x15 && ~x47 && ~x1 )
						nx_state = s183;
					else if( ~x42 && ~x12 && x44 && x14 && ~x3 && x2 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && ~x12 && x44 && x14 && ~x3 && x2 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x42 && ~x12 && x44 && x14 && ~x3 && x2 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && ~x12 && x44 && x14 && ~x3 && ~x2 )
						nx_state = s183;
					else if( ~x42 && ~x12 && x44 && ~x14 && x10 && x5 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s801;
						end
					else if( ~x42 && ~x12 && x44 && ~x14 && x10 && ~x5 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x42 && ~x12 && x44 && ~x14 && x10 && ~x5 && ~x32 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x42 && ~x12 && x44 && ~x14 && ~x10 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x42 && ~x12 && x44 && ~x14 && ~x10 && ~x3 && x2 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x42 && ~x12 && x44 && ~x14 && ~x10 && ~x3 && x2 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x42 && ~x12 && x44 && ~x14 && ~x10 && ~x3 && x2 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x42 && ~x12 && x44 && ~x14 && ~x10 && ~x3 && x2 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && ~x12 && x44 && ~x14 && ~x10 && ~x3 && x2 && x15 && ~x47 && ~x1 )
						nx_state = s183;
					else if( ~x42 && ~x12 && x44 && ~x14 && ~x10 && ~x3 && x2 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && ~x12 && x44 && ~x14 && ~x10 && ~x3 && x2 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x42 && ~x12 && x44 && ~x14 && ~x10 && ~x3 && x2 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && ~x12 && x44 && ~x14 && ~x10 && ~x3 && ~x2 )
						nx_state = s183;
					else if( ~x42 && ~x12 && ~x44 && x45 && x41 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s902;
						end
					else if( ~x42 && ~x12 && ~x44 && x45 && ~x41 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x42 && ~x12 && ~x44 && x45 && ~x41 && ~x3 && x2 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x42 && ~x12 && ~x44 && x45 && ~x41 && ~x3 && x2 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x42 && ~x12 && ~x44 && x45 && ~x41 && ~x3 && x2 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x42 && ~x12 && ~x44 && x45 && ~x41 && ~x3 && x2 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && ~x12 && ~x44 && x45 && ~x41 && ~x3 && x2 && x15 && ~x47 && ~x1 )
						nx_state = s183;
					else if( ~x42 && ~x12 && ~x44 && x45 && ~x41 && ~x3 && x2 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && ~x12 && ~x44 && x45 && ~x41 && ~x3 && x2 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x42 && ~x12 && ~x44 && x45 && ~x41 && ~x3 && x2 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && ~x12 && ~x44 && x45 && ~x41 && ~x3 && ~x2 )
						nx_state = s183;
					else if( ~x42 && ~x12 && ~x44 && ~x45 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x42 && ~x12 && ~x44 && ~x45 && ~x3 && x2 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x42 && ~x12 && ~x44 && ~x45 && ~x3 && x2 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x42 && ~x12 && ~x44 && ~x45 && ~x3 && x2 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x42 && ~x12 && ~x44 && ~x45 && ~x3 && x2 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && ~x12 && ~x44 && ~x45 && ~x3 && x2 && x15 && ~x47 && ~x1 )
						nx_state = s183;
					else if( ~x42 && ~x12 && ~x44 && ~x45 && ~x3 && x2 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && ~x12 && ~x44 && ~x45 && ~x3 && x2 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x42 && ~x12 && ~x44 && ~x45 && ~x3 && x2 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && ~x12 && ~x44 && ~x45 && ~x3 && ~x2 )
						nx_state = s183;
					else nx_state = s183;
				s184 : if( x69 && x65 )
						begin
							y15 = 1'b1;	y21 = 1'b1;	y28 = 1'b1;	
							nx_state = s832;
						end
					else if( x69 && ~x65 && x66 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && ~x65 && ~x66 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x69 && x62 && x64 && x61 && x17 && x19 && x10 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( ~x69 && x62 && x64 && x61 && x17 && x19 && ~x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x69 && x62 && x64 && x61 && x17 && ~x19 )
						nx_state = s184;
					else if( ~x69 && x62 && x64 && x61 && ~x17 && x20 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x69 && x62 && x64 && x61 && ~x17 && ~x20 && x2 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x62 && x64 && x61 && ~x17 && ~x20 && ~x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x62 && x64 && ~x61 && x11 && x10 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( ~x69 && x62 && x64 && ~x61 && x11 && ~x10 )
						begin
							y13 = 1'b1;	
							nx_state = s800;
						end
					else if( ~x69 && x62 && x64 && ~x61 && ~x11 && x10 && x12 && x4 && x1 )
						nx_state = s184;
					else if( ~x69 && x62 && x64 && ~x61 && ~x11 && x10 && x12 && x4 && ~x1 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x69 && x62 && x64 && ~x61 && ~x11 && x10 && x12 && ~x4 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x62 && x64 && ~x61 && ~x11 && x10 && ~x12 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && x62 && x64 && ~x61 && ~x11 && ~x10 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && x62 && ~x64 && x14 && x17 && x19 && x10 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( ~x69 && x62 && ~x64 && x14 && x17 && x19 && ~x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x69 && x62 && ~x64 && x14 && x17 && ~x19 )
						nx_state = s184;
					else if( ~x69 && x62 && ~x64 && x14 && ~x17 && x20 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x62 && ~x64 && x14 && ~x17 && ~x20 && x2 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x62 && ~x64 && x14 && ~x17 && ~x20 && ~x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x62 && ~x64 && ~x14 && x11 && x10 )
						nx_state = s1;
					else if( ~x69 && x62 && ~x64 && ~x14 && x11 && ~x10 )
						begin
							y13 = 1'b1;	
							nx_state = s800;
						end
					else if( ~x69 && x62 && ~x64 && ~x14 && ~x11 && x12 && x10 && x4 && x1 )
						nx_state = s184;
					else if( ~x69 && x62 && ~x64 && ~x14 && ~x11 && x12 && x10 && x4 && ~x1 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x69 && x62 && ~x64 && ~x14 && ~x11 && x12 && x10 && ~x4 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x62 && ~x64 && ~x14 && ~x11 && x12 && ~x10 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && x62 && ~x64 && ~x14 && ~x11 && ~x12 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && ~x62 && x11 && x43 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( ~x69 && ~x62 && x11 && ~x43 && x44 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( ~x69 && ~x62 && x11 && ~x43 && ~x44 && x45 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( ~x69 && ~x62 && x11 && ~x43 && ~x44 && ~x45 && x10 && x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( ~x69 && ~x62 && x11 && ~x43 && ~x44 && ~x45 && x10 && ~x32 && x33 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && ~x62 && x11 && ~x43 && ~x44 && ~x45 && x10 && ~x32 && ~x33 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && ~x62 && x11 && ~x43 && ~x44 && ~x45 && ~x10 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( ~x69 && ~x62 && ~x11 && x12 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( ~x69 && ~x62 && ~x11 && ~x12 && x13 && x14 && x41 && x37 && x2 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && ~x62 && ~x11 && ~x12 && x13 && x14 && x41 && x37 && ~x2 )
						nx_state = s184;
					else if( ~x69 && ~x62 && ~x11 && ~x12 && x13 && x14 && x41 && ~x37 && x2 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x69 && ~x62 && ~x11 && ~x12 && x13 && x14 && x41 && ~x37 && ~x2 )
						nx_state = s184;
					else if( ~x69 && ~x62 && ~x11 && ~x12 && x13 && x14 && ~x41 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( ~x69 && ~x62 && ~x11 && ~x12 && x13 && ~x14 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( ~x69 && ~x62 && ~x11 && ~x12 && ~x13 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else nx_state = s184;
				s185 : if( x70 && x63 && x64 && x11 && x43 && x41 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( x70 && x63 && x64 && x11 && x43 && x41 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( x70 && x63 && x64 && x11 && x43 && x41 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( x70 && x63 && x64 && x11 && x43 && x41 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x70 && x63 && x64 && x11 && x43 && x41 && x15 && ~x47 && ~x1 )
						nx_state = s185;
					else if( x70 && x63 && x64 && x11 && x43 && x41 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x70 && x63 && x64 && x11 && x43 && x41 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x70 && x63 && x64 && x11 && x43 && x41 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x70 && x63 && x64 && x11 && x43 && ~x41 && x4 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( x70 && x63 && x64 && x11 && x43 && ~x41 && x4 && ~x2 )
						nx_state = s185;
					else if( x70 && x63 && x64 && x11 && x43 && ~x41 && ~x4 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x70 && x63 && x64 && x11 && x43 && ~x41 && ~x4 && ~x2 )
						nx_state = s185;
					else if( x70 && x63 && x64 && x11 && ~x43 && x13 && x4 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( x70 && x63 && x64 && x11 && ~x43 && x13 && x4 && ~x2 )
						nx_state = s185;
					else if( x70 && x63 && x64 && x11 && ~x43 && x13 && ~x4 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x70 && x63 && x64 && x11 && ~x43 && x13 && ~x4 && ~x2 )
						nx_state = s185;
					else if( x70 && x63 && x64 && x11 && ~x43 && ~x13 && x45 && x41 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( x70 && x63 && x64 && x11 && ~x43 && ~x13 && x45 && x41 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( x70 && x63 && x64 && x11 && ~x43 && ~x13 && x45 && x41 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( x70 && x63 && x64 && x11 && ~x43 && ~x13 && x45 && x41 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x70 && x63 && x64 && x11 && ~x43 && ~x13 && x45 && x41 && x15 && ~x47 && ~x1 )
						nx_state = s185;
					else if( x70 && x63 && x64 && x11 && ~x43 && ~x13 && x45 && x41 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x70 && x63 && x64 && x11 && ~x43 && ~x13 && x45 && x41 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x70 && x63 && x64 && x11 && ~x43 && ~x13 && x45 && x41 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x70 && x63 && x64 && x11 && ~x43 && ~x13 && x45 && ~x41 && x4 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( x70 && x63 && x64 && x11 && ~x43 && ~x13 && x45 && ~x41 && x4 && ~x2 )
						nx_state = s185;
					else if( x70 && x63 && x64 && x11 && ~x43 && ~x13 && x45 && ~x41 && ~x4 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x70 && x63 && x64 && x11 && ~x43 && ~x13 && x45 && ~x41 && ~x4 && ~x2 )
						nx_state = s185;
					else if( x70 && x63 && x64 && x11 && ~x43 && ~x13 && ~x45 && x4 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( x70 && x63 && x64 && x11 && ~x43 && ~x13 && ~x45 && x4 && ~x2 )
						nx_state = s185;
					else if( x70 && x63 && x64 && x11 && ~x43 && ~x13 && ~x45 && ~x4 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x70 && x63 && x64 && x11 && ~x43 && ~x13 && ~x45 && ~x4 && ~x2 )
						nx_state = s185;
					else if( x70 && x63 && x64 && ~x11 && x12 && x41 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( x70 && x63 && x64 && ~x11 && x12 && x41 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( x70 && x63 && x64 && ~x11 && x12 && x41 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( x70 && x63 && x64 && ~x11 && x12 && x41 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x70 && x63 && x64 && ~x11 && x12 && x41 && x15 && ~x47 && ~x1 )
						nx_state = s185;
					else if( x70 && x63 && x64 && ~x11 && x12 && x41 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x70 && x63 && x64 && ~x11 && x12 && x41 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x70 && x63 && x64 && ~x11 && x12 && x41 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x70 && x63 && x64 && ~x11 && x12 && ~x41 && x4 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( x70 && x63 && x64 && ~x11 && x12 && ~x41 && x4 && ~x2 )
						nx_state = s185;
					else if( x70 && x63 && x64 && ~x11 && x12 && ~x41 && ~x4 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x70 && x63 && x64 && ~x11 && x12 && ~x41 && ~x4 && ~x2 )
						nx_state = s185;
					else if( x70 && x63 && x64 && ~x11 && ~x12 && x44 && x10 && x14 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && x44 && x10 && x14 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && x44 && x10 && x14 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && x44 && x10 && x14 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && x44 && x10 && x14 && x15 && ~x47 && ~x1 )
						nx_state = s185;
					else if( x70 && x63 && x64 && ~x11 && ~x12 && x44 && x10 && x14 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && x44 && x10 && x14 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && x44 && x10 && x14 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && x44 && x10 && ~x14 && x1 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s99;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && x44 && x10 && ~x14 && ~x1 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && x44 && ~x10 && x4 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && x44 && ~x10 && x4 && ~x2 )
						nx_state = s185;
					else if( x70 && x63 && x64 && ~x11 && ~x12 && x44 && ~x10 && ~x4 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && x44 && ~x10 && ~x4 && ~x2 )
						nx_state = s185;
					else if( x70 && x63 && x64 && ~x11 && ~x12 && ~x44 && x45 && x41 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && ~x44 && x45 && x41 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && ~x44 && x45 && x41 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && ~x44 && x45 && x41 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && ~x44 && x45 && x41 && x15 && ~x47 && ~x1 )
						nx_state = s185;
					else if( x70 && x63 && x64 && ~x11 && ~x12 && ~x44 && x45 && x41 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && ~x44 && x45 && x41 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && ~x44 && x45 && x41 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && ~x44 && x45 && ~x41 && x4 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && ~x44 && x45 && ~x41 && x4 && ~x2 )
						nx_state = s185;
					else if( x70 && x63 && x64 && ~x11 && ~x12 && ~x44 && x45 && ~x41 && ~x4 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && ~x44 && x45 && ~x41 && ~x4 && ~x2 )
						nx_state = s185;
					else if( x70 && x63 && x64 && ~x11 && ~x12 && ~x44 && ~x45 && x4 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && ~x44 && ~x45 && x4 && ~x2 )
						nx_state = s185;
					else if( x70 && x63 && x64 && ~x11 && ~x12 && ~x44 && ~x45 && ~x4 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x70 && x63 && x64 && ~x11 && ~x12 && ~x44 && ~x45 && ~x4 && ~x2 )
						nx_state = s185;
					else if( x70 && x63 && ~x64 && x15 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( x70 && x63 && ~x64 && x15 && ~x5 && x34 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x70 && x63 && ~x64 && x15 && ~x5 && ~x34 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x70 && x63 && ~x64 && ~x15 && x35 )
						nx_state = s1;
					else if( x70 && x63 && ~x64 && ~x15 && ~x35 && x13 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( x70 && x63 && ~x64 && ~x15 && ~x35 && ~x13 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( x70 && ~x63 && x40 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && x40 && ~x5 && x34 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s736;
						end
					else if( x70 && ~x63 && x40 && ~x5 && ~x34 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( x70 && ~x63 && ~x40 && x35 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x70 && ~x63 && ~x40 && ~x35 && x13 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( x70 && ~x63 && ~x40 && ~x35 && ~x13 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( ~x70 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x70 && ~x5 && x17 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x70 && ~x5 && ~x17 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else nx_state = s185;
				s186 : if( x70 && x63 && x64 && x55 && x30 && x16 && x37 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	y34 = 1'b1;	
							nx_state = s904;
						end
					else if( x70 && x63 && x64 && x55 && x30 && x16 && ~x37 && x39 && x19 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( x70 && x63 && x64 && x55 && x30 && x16 && ~x37 && x39 && ~x19 && x26 && x5 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s734;
						end
					else if( x70 && x63 && x64 && x55 && x30 && x16 && ~x37 && x39 && ~x19 && x26 && ~x5 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s735;
						end
					else if( x70 && x63 && x64 && x55 && x30 && x16 && ~x37 && x39 && ~x19 && ~x26 )
						begin
							y11 = 1'b1;	y36 = 1'b1;	
							nx_state = s739;
						end
					else if( x70 && x63 && x64 && x55 && x30 && x16 && ~x37 && ~x39 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( x70 && x63 && x64 && x55 && x30 && ~x16 && x41 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && x63 && x64 && x55 && x30 && ~x16 && ~x41 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( x70 && x63 && x64 && x55 && ~x30 && x36 && x9 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( x70 && x63 && x64 && x55 && ~x30 && x36 && ~x9 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s443;
						end
					else if( x70 && x63 && x64 && x55 && ~x30 && ~x36 && x3 && x42 )
						nx_state = s186;
					else if( x70 && x63 && x64 && x55 && ~x30 && ~x36 && x3 && ~x42 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( x70 && x63 && x64 && x55 && ~x30 && ~x36 && ~x3 && x11 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( x70 && x63 && x64 && x55 && ~x30 && ~x36 && ~x3 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( x70 && x63 && x64 && ~x55 && x51 && x24 && x5 && x36 )
						nx_state = s186;
					else if( x70 && x63 && x64 && ~x55 && x51 && x24 && x5 && ~x36 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s906;
						end
					else if( x70 && x63 && x64 && ~x55 && x51 && x24 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( x70 && x63 && x64 && ~x55 && x51 && ~x24 && x31 && x29 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s906;
						end
					else if( x70 && x63 && x64 && ~x55 && x51 && ~x24 && x31 && ~x29 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( x70 && x63 && x64 && ~x55 && x51 && ~x24 && ~x31 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s906;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x51 && x42 && x35 && x36 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s906;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x51 && x42 && x35 && ~x36 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x51 && x42 && ~x35 && x58 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x51 && x42 && ~x35 && ~x58 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x51 && ~x42 && x52 && x35 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s443;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x51 && ~x42 && x52 && ~x35 && x58 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x51 && ~x42 && x52 && ~x35 && ~x58 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x51 && ~x42 && ~x52 && x34 && x37 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x51 && ~x42 && ~x52 && x34 && ~x37 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x51 && ~x42 && ~x52 && ~x34 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( x70 && x63 && ~x64 && x15 && x30 && x16 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( x70 && x63 && ~x64 && x15 && x30 && x16 && ~x6 && x8 && x19 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( x70 && x63 && ~x64 && x15 && x30 && x16 && ~x6 && x8 && ~x19 && x26 && x5 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x70 && x63 && ~x64 && x15 && x30 && x16 && ~x6 && x8 && ~x19 && x26 && ~x5 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s192;
						end
					else if( x70 && x63 && ~x64 && x15 && x30 && x16 && ~x6 && x8 && ~x19 && ~x26 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s738;
						end
					else if( x70 && x63 && ~x64 && x15 && x30 && x16 && ~x6 && ~x8 )
						nx_state = s1;
					else if( x70 && x63 && ~x64 && x15 && x30 && ~x16 && x10 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && x63 && ~x64 && x15 && x30 && ~x16 && ~x10 )
						nx_state = s1;
					else if( x70 && x63 && ~x64 && x15 && ~x30 && x5 && x9 )
						nx_state = s1;
					else if( x70 && x63 && ~x64 && x15 && ~x30 && x5 && ~x9 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s443;
						end
					else if( x70 && x63 && ~x64 && x15 && ~x30 && ~x5 && x11 && x3 )
						nx_state = s186;
					else if( x70 && x63 && ~x64 && x15 && ~x30 && ~x5 && x11 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x70 && x63 && ~x64 && x15 && ~x30 && ~x5 && ~x11 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( x70 && x63 && ~x64 && x15 && ~x30 && ~x5 && ~x11 && ~x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x70 && x63 && ~x64 && ~x15 && x48 && x24 && x5 && x36 )
						nx_state = s186;
					else if( x70 && x63 && ~x64 && ~x15 && x48 && x24 && x5 && ~x36 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( x70 && x63 && ~x64 && ~x15 && x48 && x24 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( x70 && x63 && ~x64 && ~x15 && x48 && ~x24 && x31 && x29 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( x70 && x63 && ~x64 && ~x15 && x48 && ~x24 && x31 && ~x29 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( x70 && x63 && ~x64 && ~x15 && x48 && ~x24 && ~x31 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( x70 && x63 && ~x64 && ~x15 && ~x48 && x11 && x35 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( x70 && x63 && ~x64 && ~x15 && ~x48 && x11 && x35 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( x70 && x63 && ~x64 && ~x15 && ~x48 && x11 && ~x35 && x21 )
						nx_state = s1;
					else if( x70 && x63 && ~x64 && ~x15 && ~x48 && x11 && ~x35 && ~x21 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( x70 && x63 && ~x64 && ~x15 && ~x48 && ~x11 && x45 && x35 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s443;
						end
					else if( x70 && x63 && ~x64 && ~x15 && ~x48 && ~x11 && x45 && ~x35 && x21 )
						nx_state = s1;
					else if( x70 && x63 && ~x64 && ~x15 && ~x48 && ~x11 && x45 && ~x35 && ~x21 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( x70 && x63 && ~x64 && ~x15 && ~x48 && ~x11 && ~x45 && x3 && x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( x70 && x63 && ~x64 && ~x15 && ~x48 && ~x11 && ~x45 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( x70 && x63 && ~x64 && ~x15 && ~x48 && ~x11 && ~x45 && ~x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( x70 && ~x63 && x64 && x40 && x30 && x16 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( x70 && ~x63 && x64 && x40 && x30 && x16 && ~x6 && x8 && x19 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( x70 && ~x63 && x64 && x40 && x30 && x16 && ~x6 && x8 && ~x19 && x26 && x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s736;
						end
					else if( x70 && ~x63 && x64 && x40 && x30 && x16 && ~x6 && x8 && ~x19 && x26 && ~x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( x70 && ~x63 && x64 && x40 && x30 && x16 && ~x6 && x8 && ~x19 && ~x26 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s738;
						end
					else if( x70 && ~x63 && x64 && x40 && x30 && x16 && ~x6 && ~x8 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x70 && ~x63 && x64 && x40 && x30 && ~x16 && x10 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && ~x63 && x64 && x40 && x30 && ~x16 && ~x10 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x70 && ~x63 && x64 && x40 && ~x30 && x5 && x9 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x70 && ~x63 && x64 && x40 && ~x30 && x5 && ~x9 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s443;
						end
					else if( x70 && ~x63 && x64 && x40 && ~x30 && ~x5 && x11 && x3 )
						nx_state = s186;
					else if( x70 && ~x63 && x64 && x40 && ~x30 && ~x5 && x11 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( x70 && ~x63 && x64 && x40 && ~x30 && ~x5 && ~x11 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && x64 && x40 && ~x30 && ~x5 && ~x11 && ~x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x70 && ~x63 && x64 && ~x40 && x51 && x24 && x5 && x36 )
						nx_state = s186;
					else if( x70 && ~x63 && x64 && ~x40 && x51 && x24 && x5 && ~x36 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( x70 && ~x63 && x64 && ~x40 && x51 && x24 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && x64 && ~x40 && x51 && ~x24 && x31 && x29 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( x70 && ~x63 && x64 && ~x40 && x51 && ~x24 && x31 && ~x29 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && x64 && ~x40 && x51 && ~x24 && ~x31 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( x70 && ~x63 && x64 && ~x40 && ~x51 && x11 && x35 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( x70 && ~x63 && x64 && ~x40 && ~x51 && x11 && x35 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && x64 && ~x40 && ~x51 && x11 && ~x35 && x41 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x70 && ~x63 && x64 && ~x40 && ~x51 && x11 && ~x35 && ~x41 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && x64 && ~x40 && ~x51 && ~x11 && x49 && x35 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s443;
						end
					else if( x70 && ~x63 && x64 && ~x40 && ~x51 && ~x11 && x49 && ~x35 && x41 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x70 && ~x63 && x64 && ~x40 && ~x51 && ~x11 && x49 && ~x35 && ~x41 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && x64 && ~x40 && ~x51 && ~x11 && ~x49 && x3 && x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( x70 && ~x63 && x64 && ~x40 && ~x51 && ~x11 && ~x49 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && x64 && ~x40 && ~x51 && ~x11 && ~x49 && ~x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x30 && x16 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x30 && x16 && ~x6 && x8 && x19 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x30 && x16 && ~x6 && x8 && ~x19 && x26 && x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s737;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x30 && x16 && ~x6 && x8 && ~x19 && x26 && ~x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x30 && x16 && ~x6 && x8 && ~x19 && ~x26 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s738;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x30 && x16 && ~x6 && ~x8 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x30 && ~x16 && x10 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x30 && ~x16 && ~x10 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x70 && ~x63 && ~x64 && x44 && ~x30 && x5 && x9 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x70 && ~x63 && ~x64 && x44 && ~x30 && x5 && ~x9 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s907;
						end
					else if( x70 && ~x63 && ~x64 && x44 && ~x30 && ~x5 && x43 && x11 )
						nx_state = s186;
					else if( x70 && ~x63 && ~x64 && x44 && ~x30 && ~x5 && x43 && ~x11 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && ~x64 && x44 && ~x30 && ~x5 && ~x43 && x11 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s870;
						end
					else if( x70 && ~x63 && ~x64 && x44 && ~x30 && ~x5 && ~x43 && ~x11 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s867;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && x51 && x24 && x5 && x36 )
						nx_state = s186;
					else if( x70 && ~x63 && ~x64 && ~x44 && x51 && x24 && x5 && ~x36 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && x51 && x24 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && x51 && ~x24 && x31 && x29 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && x51 && ~x24 && x31 && ~x29 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && x51 && ~x24 && ~x31 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && ~x51 && x11 && x35 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && ~x51 && x11 && x35 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && ~x51 && x11 && ~x35 && x45 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && ~x51 && x11 && ~x35 && ~x45 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && ~x51 && ~x11 && x52 && x35 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s907;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && ~x51 && ~x11 && x52 && ~x35 && x45 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && ~x51 && ~x11 && x52 && ~x35 && ~x45 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && ~x51 && ~x11 && ~x52 && x3 && x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s868;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && ~x51 && ~x11 && ~x52 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && ~x51 && ~x11 && ~x52 && ~x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( ~x70 && x30 && x16 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( ~x70 && x30 && x16 && ~x6 && x8 && x19 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( ~x70 && x30 && x16 && ~x6 && x8 && ~x19 && x26 && x5 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x70 && x30 && x16 && ~x6 && x8 && ~x19 && x26 && ~x5 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x70 && x30 && x16 && ~x6 && x8 && ~x19 && ~x26 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s738;
						end
					else if( ~x70 && x30 && x16 && ~x6 && ~x8 )
						nx_state = s1;
					else if( ~x70 && x30 && ~x16 && x10 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x70 && x30 && ~x16 && ~x10 )
						nx_state = s1;
					else if( ~x70 && ~x30 && x5 && x9 )
						nx_state = s1;
					else if( ~x70 && ~x30 && x5 && ~x9 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s443;
						end
					else if( ~x70 && ~x30 && ~x5 && x11 && x3 )
						nx_state = s186;
					else if( ~x70 && ~x30 && ~x5 && x11 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x70 && ~x30 && ~x5 && ~x11 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x70 && ~x30 && ~x5 && ~x11 && ~x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else nx_state = s186;
				s187 : if( x70 && x63 && x64 && x55 && x43 && x27 && x33 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s908;
						end
					else if( x70 && x63 && x64 && x55 && x43 && x27 && ~x33 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && x63 && x64 && x55 && x43 && x27 && ~x33 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && x63 && x64 && x55 && x43 && ~x27 && x29 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s909;
						end
					else if( x70 && x63 && x64 && x55 && x43 && ~x27 && x29 && ~x1 )
						nx_state = s187;
					else if( x70 && x63 && x64 && x55 && x43 && ~x27 && ~x29 )
						nx_state = s187;
					else if( x70 && x63 && x64 && x55 && ~x43 && x29 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( x70 && x63 && x64 && x55 && ~x43 && ~x29 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s910;
						end
					else if( x70 && x63 && x64 && ~x55 && x48 )
						begin
							y13 = 1'b1;	y36 = 1'b1;	
							nx_state = s911;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x48 && x57 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s735;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x48 && ~x57 )
						nx_state = s187;
					else if( x70 && x63 && ~x64 && x15 && x12 && x27 && x33 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x70 && x63 && ~x64 && x15 && x12 && x27 && ~x33 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && x63 && ~x64 && x15 && x12 && x27 && ~x33 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && x63 && ~x64 && x15 && x12 && ~x27 && x29 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( x70 && x63 && ~x64 && x15 && x12 && ~x27 && x29 && ~x1 )
						nx_state = s187;
					else if( x70 && x63 && ~x64 && x15 && x12 && ~x27 && ~x29 )
						nx_state = s187;
					else if( x70 && x63 && ~x64 && x15 && ~x12 && x29 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( x70 && x63 && ~x64 && x15 && ~x12 && ~x29 )
						begin
							y12 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s912;
						end
					else if( x70 && x63 && ~x64 && ~x15 && x17 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s913;
						end
					else if( x70 && x63 && ~x64 && ~x15 && ~x17 && x41 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s192;
						end
					else if( x70 && x63 && ~x64 && ~x15 && ~x17 && ~x41 )
						nx_state = s187;
					else if( x70 && ~x63 && x40 && x12 && x27 && x33 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( x70 && ~x63 && x40 && x12 && x27 && ~x33 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && ~x63 && x40 && x12 && x27 && ~x33 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && ~x63 && x40 && x12 && ~x27 && x29 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( x70 && ~x63 && x40 && x12 && ~x27 && x29 && ~x1 )
						nx_state = s187;
					else if( x70 && ~x63 && x40 && x12 && ~x27 && ~x29 )
						nx_state = s187;
					else if( x70 && ~x63 && x40 && ~x12 && x29 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( x70 && ~x63 && x40 && ~x12 && ~x29 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s910;
						end
					else if( x70 && ~x63 && ~x40 && x17 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s913;
						end
					else if( x70 && ~x63 && ~x40 && ~x17 && x43 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( x70 && ~x63 && ~x40 && ~x17 && ~x43 )
						nx_state = s187;
					else if( ~x70 && x12 && x27 && x20 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x70 && x12 && x27 && ~x20 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x70 && x12 && x27 && ~x20 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x70 && x12 && ~x27 && x29 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x70 && x12 && ~x27 && x29 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x70 && x12 && ~x27 && ~x29 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( ~x70 && x12 && ~x27 && ~x29 && ~x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x70 && ~x12 && x29 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( ~x70 && ~x12 && ~x29 )
						begin
							y12 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s912;
						end
					else nx_state = s187;
				s188 : if( x70 && x63 && x15 && x7 && x35 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( x70 && x63 && x15 && x7 && x35 && ~x1 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && x63 && x15 && x7 && ~x35 && x1 )
						nx_state = s188;
					else if( x70 && x63 && x15 && x7 && ~x35 && ~x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x70 && x63 && x15 && ~x7 )
						nx_state = s188;
					else if( x70 && x63 && ~x15 && x3 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x70 && x63 && ~x15 && ~x3 && x2 )
						begin
							y12 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s912;
						end
					else if( x70 && x63 && ~x15 && ~x3 && ~x2 && x28 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x70 && x63 && ~x15 && ~x3 && ~x2 && ~x28 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && ~x63 && x64 && x40 && x7 && x35 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( x70 && ~x63 && x64 && x40 && x7 && x35 && ~x1 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && ~x63 && x64 && x40 && x7 && ~x35 && x1 )
						nx_state = s188;
					else if( x70 && ~x63 && x64 && x40 && x7 && ~x35 && ~x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x70 && ~x63 && x64 && x40 && ~x7 )
						nx_state = s188;
					else if( x70 && ~x63 && x64 && ~x40 && x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( x70 && ~x63 && x64 && ~x40 && ~x3 && x2 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s910;
						end
					else if( x70 && ~x63 && x64 && ~x40 && ~x3 && ~x2 && x28 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x70 && ~x63 && x64 && ~x40 && ~x3 && ~x2 && ~x28 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x35 && x36 && x7 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x35 && x36 && ~x7 )
						nx_state = s188;
					else if( x70 && ~x63 && ~x64 && x44 && x35 && ~x36 && x7 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x35 && ~x36 && ~x7 )
						nx_state = s188;
					else if( x70 && ~x63 && ~x64 && x44 && ~x35 && x37 )
						nx_state = s188;
					else if( x70 && ~x63 && ~x64 && x44 && ~x35 && ~x37 && x7 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s867;
						end
					else if( x70 && ~x63 && ~x64 && x44 && ~x35 && ~x37 && ~x7 )
						nx_state = s188;
					else if( x70 && ~x63 && ~x64 && ~x44 && x43 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && ~x43 && x2 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s910;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && ~x43 && ~x2 && x28 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s867;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && ~x43 && ~x2 && ~x28 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x70 && x7 && x15 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x70 && x7 && x15 && ~x1 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x70 && x7 && ~x15 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x70 && ~x7 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s913;
						end
					else nx_state = s188;
				s189 : if( x70 && x63 && x64 && x55 && x24 && x26 && x7 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s906;
						end
					else if( x70 && x63 && x64 && x55 && x24 && x26 && ~x7 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s280;
						end
					else if( x70 && x63 && x64 && x55 && x24 && ~x26 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s914;
						end
					else if( x70 && x63 && x64 && x55 && ~x24 && x28 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( x70 && x63 && x64 && x55 && ~x24 && ~x28 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( x70 && x63 && x64 && ~x55 && x31 && x50 && x10 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s734;
						end
					else if( x70 && x63 && x64 && ~x55 && x31 && x50 && ~x10 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s914;
						end
					else if( x70 && x63 && x64 && ~x55 && x31 && ~x50 )
						nx_state = s189;
					else if( x70 && x63 && x64 && ~x55 && ~x31 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s914;
						end
					else if( x70 && x63 && ~x64 && x15 && x24 && x26 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( x70 && x63 && ~x64 && x15 && x24 && x26 && ~x7 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s280;
						end
					else if( x70 && x63 && ~x64 && x15 && x24 && ~x26 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x70 && x63 && ~x64 && x15 && ~x24 && x28 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( x70 && x63 && ~x64 && x15 && ~x24 && ~x28 )
						nx_state = s1;
					else if( x70 && x63 && ~x64 && ~x15 && x31 && x19 && x10 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x70 && x63 && ~x64 && ~x15 && x31 && x19 && ~x10 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x70 && x63 && ~x64 && ~x15 && x31 && ~x19 )
						nx_state = s189;
					else if( x70 && x63 && ~x64 && ~x15 && ~x31 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x70 && ~x63 && x64 && x40 && x24 && x26 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( x70 && ~x63 && x64 && x40 && x24 && x26 && ~x7 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s280;
						end
					else if( x70 && ~x63 && x64 && x40 && x24 && ~x26 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s915;
						end
					else if( x70 && ~x63 && x64 && x40 && ~x24 && x28 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( x70 && ~x63 && x64 && x40 && ~x24 && ~x28 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x70 && ~x63 && x64 && ~x40 && x31 && x19 && x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s736;
						end
					else if( x70 && ~x63 && x64 && ~x40 && x31 && x19 && ~x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s915;
						end
					else if( x70 && ~x63 && x64 && ~x40 && x31 && ~x19 )
						nx_state = s189;
					else if( x70 && ~x63 && x64 && ~x40 && ~x31 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s915;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x24 && x26 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x24 && x26 && ~x7 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y30 = 1'b1;	
							nx_state = s916;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x24 && ~x26 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s915;
						end
					else if( x70 && ~x63 && ~x64 && x44 && ~x24 && x28 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s868;
						end
					else if( x70 && ~x63 && ~x64 && x44 && ~x24 && ~x28 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && x31 && x19 && x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s737;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && x31 && x19 && ~x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s915;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && x31 && ~x19 )
						nx_state = s189;
					else if( x70 && ~x63 && ~x64 && ~x44 && ~x31 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s915;
						end
					else if( ~x70 && x24 && x26 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x70 && x24 && x26 && ~x7 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s280;
						end
					else if( ~x70 && x24 && ~x26 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x70 && ~x24 && x28 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( ~x70 && ~x24 && ~x28 )
						nx_state = s1;
					else nx_state = s189;
				s190 : if( x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x2 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else nx_state = s190;
				s191 : if( x70 && x63 && x15 && x14 && x8 && x10 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && x63 && x15 && x14 && x8 && ~x10 )
						nx_state = s1;
					else if( x70 && x63 && x15 && x14 && ~x8 && x30 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( x70 && x63 && x15 && x14 && ~x8 && x30 && ~x1 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x70 && x63 && x15 && x14 && ~x8 && x30 && ~x1 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x70 && x63 && x15 && x14 && ~x8 && ~x30 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && x63 && x15 && ~x14 && x32 && x3 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s192;
						end
					else if( x70 && x63 && x15 && ~x14 && x32 && ~x3 )
						nx_state = s191;
					else if( x70 && x63 && x15 && ~x14 && ~x32 && x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && x63 && x15 && ~x14 && ~x32 && ~x3 )
						nx_state = s191;
					else if( x70 && x63 && ~x15 && x16 && x43 && x29 && x40 && x27 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( x70 && x63 && ~x15 && x16 && x43 && x29 && x40 && ~x27 )
						nx_state = s191;
					else if( x70 && x63 && ~x15 && x16 && x43 && x29 && ~x40 && x27 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && x63 && ~x15 && x16 && x43 && x29 && ~x40 && ~x27 )
						nx_state = s191;
					else if( x70 && x63 && ~x15 && x16 && x43 && ~x29 && x33 && x27 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && x63 && ~x15 && x16 && x43 && ~x29 && x33 && ~x27 )
						nx_state = s191;
					else if( x70 && x63 && ~x15 && x16 && x43 && ~x29 && ~x33 && x41 && x27 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x70 && x63 && ~x15 && x16 && x43 && ~x29 && ~x33 && x41 && ~x27 )
						nx_state = s191;
					else if( x70 && x63 && ~x15 && x16 && x43 && ~x29 && ~x33 && ~x41 && x27 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && x63 && ~x15 && x16 && x43 && ~x29 && ~x33 && ~x41 && ~x27 )
						nx_state = s191;
					else if( x70 && x63 && ~x15 && x16 && ~x43 )
						nx_state = s1;
					else if( x70 && x63 && ~x15 && ~x16 && x37 && x42 && x1 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && x63 && ~x15 && ~x16 && x37 && x42 && ~x1 )
						nx_state = s191;
					else if( x70 && x63 && ~x15 && ~x16 && x37 && ~x42 )
						nx_state = s1;
					else if( x70 && x63 && ~x15 && ~x16 && ~x37 && x25 )
						nx_state = s1;
					else if( x70 && x63 && ~x15 && ~x16 && ~x37 && ~x25 && x5 && x4 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( x70 && x63 && ~x15 && ~x16 && ~x37 && ~x25 && x5 && ~x4 )
						nx_state = s191;
					else if( x70 && x63 && ~x15 && ~x16 && ~x37 && ~x25 && ~x5 && x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && x63 && ~x15 && ~x16 && ~x37 && ~x25 && ~x5 && ~x4 )
						nx_state = s191;
					else if( x70 && ~x63 && x26 && x28 && x9 && x64 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( x70 && ~x63 && x26 && x28 && x9 && ~x64 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s917;
						end
					else if( x70 && ~x63 && x26 && x28 && ~x9 && x23 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( x70 && ~x63 && x26 && x28 && ~x9 && ~x23 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( x70 && ~x63 && x26 && ~x28 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else if( x70 && ~x63 && ~x26 && x27 && x4 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else if( x70 && ~x63 && ~x26 && x27 && ~x4 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x26 && ~x27 && x28 && x64 && x2 && x24 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s920;
						end
					else if( x70 && ~x63 && ~x26 && ~x27 && x28 && x64 && x2 && ~x24 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else if( x70 && ~x63 && ~x26 && ~x27 && x28 && x64 && ~x2 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else if( x70 && ~x63 && ~x26 && ~x27 && x28 && ~x64 && x32 && x24 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s920;
						end
					else if( x70 && ~x63 && ~x26 && ~x27 && x28 && ~x64 && x32 && ~x24 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else if( x70 && ~x63 && ~x26 && ~x27 && x28 && ~x64 && ~x32 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else if( x70 && ~x63 && ~x26 && ~x27 && ~x28 && x18 && x3 && x64 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s922;
						end
					else if( x70 && ~x63 && ~x26 && ~x27 && ~x28 && x18 && x3 && ~x64 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s923;
						end
					else if( x70 && ~x63 && ~x26 && ~x27 && ~x28 && x18 && ~x3 && x4 && x64 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( x70 && ~x63 && ~x26 && ~x27 && ~x28 && x18 && ~x3 && x4 && ~x64 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s924;
						end
					else if( x70 && ~x63 && ~x26 && ~x27 && ~x28 && x18 && ~x3 && ~x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else if( x70 && ~x63 && ~x26 && ~x27 && ~x28 && ~x18 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else if( ~x70 && x44 && x14 && x8 && x10 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x70 && x44 && x14 && x8 && ~x10 )
						nx_state = s1;
					else if( ~x70 && x44 && x14 && ~x8 && x30 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x70 && x44 && x14 && ~x8 && x30 && ~x1 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x70 && x44 && x14 && ~x8 && x30 && ~x1 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x70 && x44 && x14 && ~x8 && ~x30 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x70 && x44 && ~x14 && x3 && x21 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x70 && x44 && ~x14 && x3 && ~x21 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x70 && x44 && ~x14 && ~x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x70 && ~x44 && x2 && x4 )
						begin
							y5 = 1'b1;	y13 = 1'b1;	
							nx_state = s740;
						end
					else if( ~x70 && ~x44 && x2 && ~x4 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s738;
						end
					else if( ~x70 && ~x44 && ~x2 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else nx_state = s191;
				s192 : if( x70 && x15 && x10 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x70 && x15 && ~x10 && x25 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( x70 && x15 && ~x10 && ~x25 )
						begin
							y12 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s912;
						end
					else if( x70 && ~x15 && x8 && x44 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x70 && ~x15 && x8 && ~x44 && x37 )
						nx_state = s1;
					else if( x70 && ~x15 && x8 && ~x44 && ~x37 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x70 && ~x15 && ~x8 && x48 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x70 && ~x15 && ~x8 && ~x48 && x37 )
						nx_state = s1;
					else if( x70 && ~x15 && ~x8 && ~x48 && ~x37 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x70 && x10 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x70 && ~x10 && x25 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x70 && ~x10 && ~x25 )
						begin
							y12 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s912;
						end
					else nx_state = s192;
				s193 : if( x69 && x22 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	y38 = 1'b1;	
							nx_state = s925;
						end
					else if( x69 && ~x22 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	y26 = 1'b1;	
							nx_state = s926;
						end
					else if( ~x69 && x16 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s901;
						end
					else if( ~x69 && x16 && ~x15 && x4 && x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s901;
						end
					else if( ~x69 && x16 && ~x15 && x4 && ~x5 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s627;
						end
					else if( ~x69 && x16 && ~x15 && ~x4 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s927;
						end
					else if( ~x69 && ~x16 && x15 && x6 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s927;
						end
					else if( ~x69 && ~x16 && x15 && ~x6 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s195;
						end
					else if( ~x69 && ~x16 && ~x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s901;
						end
					else nx_state = s193;
				s194 : if( x15 && x16 && x5 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else if( x15 && x16 && ~x5 && x6 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( x15 && x16 && ~x5 && ~x6 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else if( x15 && ~x16 && x6 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x15 && ~x16 && ~x6 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s438;
						end
					else if( ~x15 && x16 && x4 && x5 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x15 && x16 && x4 && ~x5 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s436;
						end
					else if( ~x15 && x16 && ~x4 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s928;
						end
					else if( ~x15 && ~x16 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else nx_state = s194;
				s195 : if( x16 && x15 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s927;
						end
					else if( x16 && ~x15 && x4 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s627;
						end
					else if( x16 && ~x15 && ~x4 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s927;
						end
					else if( ~x16 && x15 && x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s901;
						end
					else if( ~x16 && x15 && ~x12 )
						nx_state = s195;
					else if( ~x16 && ~x15 && x14 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s927;
						end
					else if( ~x16 && ~x15 && ~x14 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s451;
						end
					else nx_state = s195;
				s196 : if( x63 && x46 && x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( x63 && x46 && ~x16 && x37 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s929;
						end
					else if( x63 && x46 && ~x16 && ~x37 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( x63 && ~x46 && x47 && x4 && x36 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( x63 && ~x46 && x47 && x4 && ~x36 )
						begin
							y21 = 1'b1;	y27 = 1'b1;	
							nx_state = s930;
						end
					else if( x63 && ~x46 && x47 && ~x4 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s929;
						end
					else if( x63 && ~x46 && ~x47 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( ~x63 && x16 && x15 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( ~x63 && x16 && ~x15 && x4 && x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( ~x63 && x16 && ~x15 && x4 && ~x5 )
						begin
							y21 = 1'b1;	y27 = 1'b1;	
							nx_state = s930;
						end
					else if( ~x63 && x16 && ~x15 && ~x4 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s929;
						end
					else if( ~x63 && ~x16 && x15 && x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s929;
						end
					else if( ~x63 && ~x16 && x15 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x63 && ~x16 && ~x15 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else nx_state = s196;
				s197 : if( x15 && x16 && x64 && x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s445;
						end
					else if( x15 && x16 && x64 && ~x5 && x6 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x15 && x16 && x64 && ~x5 && ~x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s445;
						end
					else if( x15 && x16 && ~x64 && x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s931;
						end
					else if( x15 && x16 && ~x64 && ~x5 && x6 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( x15 && x16 && ~x64 && ~x5 && ~x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s931;
						end
					else if( x15 && ~x16 && x6 && x64 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x15 && ~x16 && x6 && ~x64 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s540;
						end
					else if( x15 && ~x16 && ~x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s446;
						end
					else if( ~x15 && x16 && x4 && x5 && x64 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x15 && x16 && x4 && x5 && ~x64 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s540;
						end
					else if( ~x15 && x16 && x4 && ~x5 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x15 && x16 && ~x4 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s932;
						end
					else if( ~x15 && ~x16 && x64 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s445;
						end
					else if( ~x15 && ~x16 && ~x64 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s931;
						end
					else nx_state = s197;
				s198 : if( x63 && x46 && x16 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s929;
						end
					else if( x63 && x46 && ~x16 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( x63 && x46 && ~x16 && ~x12 )
						nx_state = s198;
					else if( x63 && ~x46 && x47 && x4 )
						begin
							y21 = 1'b1;	y27 = 1'b1;	
							nx_state = s930;
						end
					else if( x63 && ~x46 && x47 && ~x4 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s929;
						end
					else if( x63 && ~x46 && ~x47 && x14 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s929;
						end
					else if( x63 && ~x46 && ~x47 && ~x14 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s322;
						end
					else if( ~x63 && x16 && x15 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s929;
						end
					else if( ~x63 && x16 && ~x15 && x4 )
						begin
							y21 = 1'b1;	y27 = 1'b1;	
							nx_state = s930;
						end
					else if( ~x63 && x16 && ~x15 && ~x4 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s929;
						end
					else if( ~x63 && ~x16 && x15 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( ~x63 && ~x16 && x15 && ~x12 )
						nx_state = s198;
					else if( ~x63 && ~x16 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s929;
						end
					else if( ~x63 && ~x16 && ~x15 && ~x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s326;
						end
					else nx_state = s198;
				s199 : if( x62 && x15 && x16 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s900;
						end
					else if( x62 && x15 && ~x16 && x5 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else if( x62 && x15 && ~x16 && ~x5 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s900;
						end
					else if( x62 && ~x15 && x16 && x4 && x5 && x1 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s900;
						end
					else if( x62 && ~x15 && x16 && x4 && x5 && ~x1 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s194;
						end
					else if( x62 && ~x15 && x16 && x4 && ~x5 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s901;
						end
					else if( x62 && ~x15 && x16 && x4 && ~x5 && ~x1 )
						begin
							y10 = 1'b1;	
							nx_state = s193;
						end
					else if( x62 && ~x15 && x16 && ~x4 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s901;
						end
					else if( x62 && ~x15 && x16 && ~x4 && ~x1 )
						begin
							y10 = 1'b1;	
							nx_state = s193;
						end
					else if( x62 && ~x15 && ~x16 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s900;
						end
					else if( ~x62 && x15 && x63 && x47 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( ~x62 && x15 && x63 && ~x47 && x36 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s440;
						end
					else if( ~x62 && x15 && x63 && ~x47 && ~x36 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( ~x62 && x15 && ~x63 && x16 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( ~x62 && x15 && ~x63 && ~x16 && x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s445;
						end
					else if( ~x62 && x15 && ~x63 && ~x16 && ~x5 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( ~x62 && ~x15 && x16 && x63 && x35 && x5 && x1 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( ~x62 && ~x15 && x16 && x63 && x35 && x5 && ~x1 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x62 && ~x15 && x16 && x63 && x35 && ~x5 && x32 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( ~x62 && ~x15 && x16 && x63 && x35 && ~x5 && ~x32 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x62 && ~x15 && x16 && x63 && ~x35 && x32 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( ~x62 && ~x15 && x16 && x63 && ~x35 && ~x32 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x62 && ~x15 && x16 && ~x63 && x4 && x5 && x1 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( ~x62 && ~x15 && x16 && ~x63 && x4 && x5 && ~x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x62 && ~x15 && x16 && ~x63 && x4 && ~x5 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( ~x62 && ~x15 && x16 && ~x63 && x4 && ~x5 && ~x1 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x62 && ~x15 && x16 && ~x63 && ~x4 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( ~x62 && ~x15 && x16 && ~x63 && ~x4 && ~x1 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x62 && ~x15 && ~x16 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else nx_state = s199;
				s200 : if( x70 && x64 && x61 && x50 && x19 && x10 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( x70 && x64 && x61 && x50 && x19 && ~x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( x70 && x64 && x61 && x50 && ~x19 )
						nx_state = s200;
					else if( x70 && x64 && x61 && ~x50 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( x70 && x64 && ~x61 && x11 && x10 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( x70 && x64 && ~x61 && x11 && ~x10 && x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x70 && x64 && ~x61 && x11 && ~x10 && ~x7 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s933;
						end
					else if( x70 && x64 && ~x61 && ~x11 && x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( x70 && x64 && ~x61 && ~x11 && ~x10 && x12 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s205;
						end
					else if( x70 && x64 && ~x61 && ~x11 && ~x10 && ~x12 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s206;
						end
					else if( x70 && x64 && ~x61 && ~x11 && ~x10 && ~x12 && ~x1 && x4 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( x70 && x64 && ~x61 && ~x11 && ~x10 && ~x12 && ~x1 && ~x4 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( x70 && ~x64 && x14 && x42 && x19 && x10 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( x70 && ~x64 && x14 && x42 && x19 && ~x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( x70 && ~x64 && x14 && x42 && ~x19 )
						nx_state = s200;
					else if( x70 && ~x64 && x14 && ~x42 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( x70 && ~x64 && ~x14 && x11 && x10 )
						nx_state = s1;
					else if( x70 && ~x64 && ~x14 && x11 && ~x10 && x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x70 && ~x64 && ~x14 && x11 && ~x10 && ~x7 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s933;
						end
					else if( x70 && ~x64 && ~x14 && ~x11 && x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( x70 && ~x64 && ~x14 && ~x11 && ~x10 && x12 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s205;
						end
					else if( x70 && ~x64 && ~x14 && ~x11 && ~x10 && ~x12 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s206;
						end
					else if( x70 && ~x64 && ~x14 && ~x11 && ~x10 && ~x12 && ~x1 && x4 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( x70 && ~x64 && ~x14 && ~x11 && ~x10 && ~x12 && ~x1 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x11 && x10 )
						nx_state = s1;
					else if( ~x70 && x11 && ~x10 && x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x70 && x11 && ~x10 && ~x7 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s280;
						end
					else if( ~x70 && ~x11 && x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x70 && ~x11 && ~x10 && x12 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s215;
						end
					else if( ~x70 && ~x11 && ~x10 && ~x12 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s216;
						end
					else if( ~x70 && ~x11 && ~x10 && ~x12 && ~x1 && x4 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x70 && ~x11 && ~x10 && ~x12 && ~x1 && ~x4 )
						nx_state = s1;
					else nx_state = s200;
				s201 : if( x28 && x64 && x57 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( x28 && x64 && ~x57 )
						nx_state = s201;
					else if( x28 && ~x64 && x21 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( x28 && ~x64 && ~x21 )
						nx_state = s201;
					else if( ~x28 && x27 && x8 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( ~x28 && x27 && ~x8 && x37 && x64 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( ~x28 && x27 && ~x8 && x37 && ~x64 )
						nx_state = s1;
					else if( ~x28 && x27 && ~x8 && ~x37 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x28 && ~x27 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else nx_state = s201;
				s202 : if( x64 && x50 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x64 && ~x50 )
						nx_state = s202;
					else if( ~x64 && x42 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x64 && ~x42 )
						nx_state = s202;
					else nx_state = s202;
				s203 : if( x70 && x64 && x61 && x16 && x54 && x29 && x59 && x27 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else if( x70 && x64 && x61 && x16 && x54 && x29 && x59 && ~x27 )
						nx_state = s203;
					else if( x70 && x64 && x61 && x16 && x54 && x29 && ~x59 && x27 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( x70 && x64 && x61 && x16 && x54 && x29 && ~x59 && ~x27 )
						nx_state = s203;
					else if( x70 && x64 && x61 && x16 && x54 && ~x29 && x33 && x27 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( x70 && x64 && x61 && x16 && x54 && ~x29 && x33 && ~x27 )
						nx_state = s203;
					else if( x70 && x64 && x61 && x16 && x54 && ~x29 && ~x33 && x57 && x27 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x70 && x64 && x61 && x16 && x54 && ~x29 && ~x33 && x57 && ~x27 )
						nx_state = s203;
					else if( x70 && x64 && x61 && x16 && x54 && ~x29 && ~x33 && ~x57 && x27 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( x70 && x64 && x61 && x16 && x54 && ~x29 && ~x33 && ~x57 && ~x27 )
						nx_state = s203;
					else if( x70 && x64 && x61 && x16 && ~x54 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( x70 && x64 && x61 && ~x16 && x37 && x56 && x1 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( x70 && x64 && x61 && ~x16 && x37 && x56 && ~x1 )
						nx_state = s203;
					else if( x70 && x64 && x61 && ~x16 && x37 && ~x56 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( x70 && x64 && x61 && ~x16 && ~x37 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( x70 && x64 && x61 && ~x16 && ~x37 && ~x25 && x5 && x4 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s593;
						end
					else if( x70 && x64 && x61 && ~x16 && ~x37 && ~x25 && x5 && ~x4 )
						nx_state = s203;
					else if( x70 && x64 && x61 && ~x16 && ~x37 && ~x25 && ~x5 && x4 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( x70 && x64 && x61 && ~x16 && ~x37 && ~x25 && ~x5 && ~x4 )
						nx_state = s203;
					else if( x70 && x64 && ~x61 && x10 && x11 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( x70 && x64 && ~x61 && x10 && ~x11 && x12 && x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( x70 && x64 && ~x61 && x10 && ~x11 && x12 && ~x2 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( x70 && x64 && ~x61 && x10 && ~x11 && ~x12 && x1 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s201;
						end
					else if( x70 && x64 && ~x61 && x10 && ~x11 && ~x12 && x1 && ~x3 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( x70 && x64 && ~x61 && x10 && ~x11 && ~x12 && x1 && ~x3 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( x70 && x64 && ~x61 && x10 && ~x11 && ~x12 && ~x1 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( x70 && x64 && ~x61 && ~x10 && x12 && x2 && x4 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( x70 && x64 && ~x61 && ~x10 && x12 && x2 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( x70 && x64 && ~x61 && ~x10 && x12 && ~x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( x70 && x64 && ~x61 && ~x10 && ~x12 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s934;
						end
					else if( x70 && x64 && ~x61 && ~x10 && ~x12 && ~x9 && x5 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( x70 && x64 && ~x61 && ~x10 && ~x12 && ~x9 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x70 && ~x64 && x14 && x16 && x26 && x29 && x27 && x18 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else if( x70 && ~x64 && x14 && x16 && x26 && x29 && x27 && ~x18 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( x70 && ~x64 && x14 && x16 && x26 && x29 && ~x27 )
						nx_state = s203;
					else if( x70 && ~x64 && x14 && x16 && x26 && ~x29 && x27 && x33 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( x70 && ~x64 && x14 && x16 && x26 && ~x29 && x27 && ~x33 && x21 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x70 && ~x64 && x14 && x16 && x26 && ~x29 && x27 && ~x33 && ~x21 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( x70 && ~x64 && x14 && x16 && x26 && ~x29 && ~x27 )
						nx_state = s203;
					else if( x70 && ~x64 && x14 && x16 && ~x26 )
						nx_state = s1;
					else if( x70 && ~x64 && x14 && ~x16 && x37 && x22 && x1 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( x70 && ~x64 && x14 && ~x16 && x37 && x22 && ~x1 )
						nx_state = s203;
					else if( x70 && ~x64 && x14 && ~x16 && x37 && ~x22 )
						nx_state = s1;
					else if( x70 && ~x64 && x14 && ~x16 && ~x37 && x25 )
						nx_state = s1;
					else if( x70 && ~x64 && x14 && ~x16 && ~x37 && ~x25 && x5 && x4 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s593;
						end
					else if( x70 && ~x64 && x14 && ~x16 && ~x37 && ~x25 && x5 && ~x4 )
						nx_state = s203;
					else if( x70 && ~x64 && x14 && ~x16 && ~x37 && ~x25 && ~x5 && x4 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( x70 && ~x64 && x14 && ~x16 && ~x37 && ~x25 && ~x5 && ~x4 )
						nx_state = s203;
					else if( x70 && ~x64 && ~x14 && x10 && x11 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( x70 && ~x64 && ~x14 && x10 && ~x11 && x12 && x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( x70 && ~x64 && ~x14 && x10 && ~x11 && x12 && ~x2 )
						nx_state = s1;
					else if( x70 && ~x64 && ~x14 && x10 && ~x11 && ~x12 && x1 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s201;
						end
					else if( x70 && ~x64 && ~x14 && x10 && ~x11 && ~x12 && x1 && ~x3 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( x70 && ~x64 && ~x14 && x10 && ~x11 && ~x12 && x1 && ~x3 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( x70 && ~x64 && ~x14 && x10 && ~x11 && ~x12 && ~x1 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( x70 && ~x64 && ~x14 && ~x10 && x12 && x2 && x4 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( x70 && ~x64 && ~x14 && ~x10 && x12 && x2 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( x70 && ~x64 && ~x14 && ~x10 && x12 && ~x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( x70 && ~x64 && ~x14 && ~x10 && ~x12 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s934;
						end
					else if( x70 && ~x64 && ~x14 && ~x10 && ~x12 && ~x9 && x5 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( x70 && ~x64 && ~x14 && ~x10 && ~x12 && ~x9 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x70 && x44 && x10 && x11 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x70 && x44 && x10 && ~x11 && x12 && x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x70 && x44 && x10 && ~x11 && x12 && ~x2 )
						nx_state = s1;
					else if( ~x70 && x44 && x10 && ~x11 && ~x12 && x1 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( ~x70 && x44 && x10 && ~x11 && ~x12 && x1 && ~x3 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x70 && x44 && x10 && ~x11 && ~x12 && x1 && ~x3 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x70 && x44 && x10 && ~x11 && ~x12 && ~x1 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x70 && x44 && ~x10 && x12 && x2 && x4 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s733;
						end
					else if( ~x70 && x44 && ~x10 && x12 && x2 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x70 && x44 && ~x10 && x12 && ~x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x70 && x44 && ~x10 && ~x12 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s816;
						end
					else if( ~x70 && x44 && ~x10 && ~x12 && ~x9 && x5 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x70 && x44 && ~x10 && ~x12 && ~x9 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x70 && ~x44 && x45 && x7 && x11 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x70 && ~x44 && x45 && x7 && ~x11 && x2 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x44 && x45 && x7 && ~x11 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && ~x44 && x45 && ~x7 && x16 && x1 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s578;
						end
					else if( ~x70 && ~x44 && x45 && ~x7 && x16 && ~x1 )
						nx_state = s203;
					else if( ~x70 && ~x44 && x45 && ~x7 && ~x16 && x1 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && ~x44 && x45 && ~x7 && ~x16 && ~x1 )
						nx_state = s203;
					else if( ~x70 && ~x44 && ~x45 && x7 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x70 && ~x44 && ~x45 && x7 && ~x1 && x2 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x44 && ~x45 && x7 && ~x1 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && ~x44 && ~x45 && ~x7 && x6 && x2 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s578;
						end
					else if( ~x70 && ~x44 && ~x45 && ~x7 && x6 && ~x2 )
						nx_state = s203;
					else if( ~x70 && ~x44 && ~x45 && ~x7 && ~x6 && x2 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && ~x44 && ~x45 && ~x7 && ~x6 && ~x2 )
						nx_state = s203;
					else nx_state = s203;
				s204 : if( x70 && x64 && x61 && x51 && x24 && x5 && x36 )
						nx_state = s204;
					else if( x70 && x64 && x61 && x51 && x24 && x5 && ~x36 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x70 && x64 && x61 && x51 && x24 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x70 && x64 && x61 && x51 && ~x24 && x31 && x29 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x70 && x64 && x61 && x51 && ~x24 && x31 && ~x29 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x70 && x64 && x61 && x51 && ~x24 && ~x31 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x70 && x64 && x61 && ~x51 && x11 && x35 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x70 && x64 && x61 && ~x51 && x11 && x35 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x70 && x64 && x61 && ~x51 && x11 && ~x35 && x60 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( x70 && x64 && x61 && ~x51 && x11 && ~x35 && ~x60 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x70 && x64 && x61 && ~x51 && ~x11 && x52 && x35 )
						begin
							y13 = 1'b1;	
							nx_state = s800;
						end
					else if( x70 && x64 && x61 && ~x51 && ~x11 && x52 && ~x35 && x60 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( x70 && x64 && x61 && ~x51 && ~x11 && x52 && ~x35 && ~x60 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x70 && x64 && x61 && ~x51 && ~x11 && ~x52 && x3 && x6 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s205;
						end
					else if( x70 && x64 && x61 && ~x51 && ~x11 && ~x52 && x3 && ~x6 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x70 && x64 && x61 && ~x51 && ~x11 && ~x52 && ~x3 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x70 && x64 && ~x61 && x11 && x10 && x4 && x5 && x3 )
						nx_state = s204;
					else if( x70 && x64 && ~x61 && x11 && x10 && x4 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( x70 && x64 && ~x61 && x11 && x10 && x4 && ~x5 && x3 )
						nx_state = s204;
					else if( x70 && x64 && ~x61 && x11 && x10 && x4 && ~x5 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x70 && x64 && ~x61 && x11 && x10 && ~x4 && x3 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x70 && x64 && ~x61 && x11 && x10 && ~x4 && ~x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x70 && x64 && ~x61 && x11 && ~x10 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s201;
						end
					else if( x70 && x64 && ~x61 && x11 && ~x10 && ~x6 && x8 && x4 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s593;
						end
					else if( x70 && x64 && ~x61 && x11 && ~x10 && ~x6 && x8 && ~x4 && x1 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( x70 && x64 && ~x61 && x11 && ~x10 && ~x6 && x8 && ~x4 && x1 && ~x3 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( x70 && x64 && ~x61 && x11 && ~x10 && ~x6 && x8 && ~x4 && ~x1 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( x70 && x64 && ~x61 && x11 && ~x10 && ~x6 && ~x8 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( x70 && x64 && ~x61 && ~x11 && x10 && x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( x70 && x64 && ~x61 && ~x11 && x10 && ~x2 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( x70 && x64 && ~x61 && ~x11 && ~x10 && x12 && x9 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( x70 && x64 && ~x61 && ~x11 && ~x10 && x12 && ~x9 )
						begin
							y13 = 1'b1;	
							nx_state = s800;
						end
					else if( x70 && x64 && ~x61 && ~x11 && ~x10 && ~x12 && x6 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x70 && x64 && ~x61 && ~x11 && ~x10 && ~x12 && ~x6 && x9 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( x70 && x64 && ~x61 && ~x11 && ~x10 && ~x12 && ~x6 && ~x9 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x70 && ~x64 && x14 && x41 && x24 && x5 && x36 )
						nx_state = s204;
					else if( x70 && ~x64 && x14 && x41 && x24 && x5 && ~x36 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x70 && ~x64 && x14 && x41 && x24 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x70 && ~x64 && x14 && x41 && ~x24 && x31 && x29 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x70 && ~x64 && x14 && x41 && ~x24 && x31 && ~x29 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x70 && ~x64 && x14 && x41 && ~x24 && ~x31 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x70 && ~x64 && x14 && ~x41 && x11 && x35 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x70 && ~x64 && x14 && ~x41 && x11 && x35 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x70 && ~x64 && x14 && ~x41 && x11 && ~x35 && x15 )
						nx_state = s1;
					else if( x70 && ~x64 && x14 && ~x41 && x11 && ~x35 && ~x15 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x70 && ~x64 && x14 && ~x41 && ~x11 && x40 && x35 )
						begin
							y13 = 1'b1;	
							nx_state = s800;
						end
					else if( x70 && ~x64 && x14 && ~x41 && ~x11 && x40 && ~x35 && x15 )
						nx_state = s1;
					else if( x70 && ~x64 && x14 && ~x41 && ~x11 && x40 && ~x35 && ~x15 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x70 && ~x64 && x14 && ~x41 && ~x11 && ~x40 && x3 && x6 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s205;
						end
					else if( x70 && ~x64 && x14 && ~x41 && ~x11 && ~x40 && x3 && ~x6 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x70 && ~x64 && x14 && ~x41 && ~x11 && ~x40 && ~x3 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x70 && ~x64 && ~x14 && x11 && x10 && x4 && x5 && x3 )
						nx_state = s204;
					else if( x70 && ~x64 && ~x14 && x11 && x10 && x4 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( x70 && ~x64 && ~x14 && x11 && x10 && x4 && ~x5 && x3 )
						nx_state = s204;
					else if( x70 && ~x64 && ~x14 && x11 && x10 && x4 && ~x5 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x70 && ~x64 && ~x14 && x11 && x10 && ~x4 && x3 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x70 && ~x64 && ~x14 && x11 && x10 && ~x4 && ~x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x70 && ~x64 && ~x14 && x11 && ~x10 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s201;
						end
					else if( x70 && ~x64 && ~x14 && x11 && ~x10 && ~x6 && x8 && x4 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s593;
						end
					else if( x70 && ~x64 && ~x14 && x11 && ~x10 && ~x6 && x8 && ~x4 && x1 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( x70 && ~x64 && ~x14 && x11 && ~x10 && ~x6 && x8 && ~x4 && x1 && ~x3 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( x70 && ~x64 && ~x14 && x11 && ~x10 && ~x6 && x8 && ~x4 && ~x1 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( x70 && ~x64 && ~x14 && x11 && ~x10 && ~x6 && ~x8 )
						nx_state = s1;
					else if( x70 && ~x64 && ~x14 && ~x11 && x10 && x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( x70 && ~x64 && ~x14 && ~x11 && x10 && ~x2 )
						nx_state = s1;
					else if( x70 && ~x64 && ~x14 && ~x11 && ~x10 && x12 && x9 )
						nx_state = s1;
					else if( x70 && ~x64 && ~x14 && ~x11 && ~x10 && x12 && ~x9 )
						begin
							y13 = 1'b1;	
							nx_state = s800;
						end
					else if( x70 && ~x64 && ~x14 && ~x11 && ~x10 && ~x12 && x6 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x70 && ~x64 && ~x14 && ~x11 && ~x10 && ~x12 && ~x6 && x9 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( x70 && ~x64 && ~x14 && ~x11 && ~x10 && ~x12 && ~x6 && ~x9 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x70 && x11 && x10 && x4 && x5 && x3 )
						nx_state = s204;
					else if( ~x70 && x11 && x10 && x4 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x70 && x11 && x10 && x4 && ~x5 && x3 )
						nx_state = s204;
					else if( ~x70 && x11 && x10 && x4 && ~x5 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x70 && x11 && x10 && ~x4 && x3 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x70 && x11 && x10 && ~x4 && ~x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x70 && x11 && ~x10 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( ~x70 && x11 && ~x10 && ~x6 && x8 && x4 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s320;
						end
					else if( ~x70 && x11 && ~x10 && ~x6 && x8 && ~x4 && x1 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x70 && x11 && ~x10 && ~x6 && x8 && ~x4 && x1 && ~x3 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s733;
						end
					else if( ~x70 && x11 && ~x10 && ~x6 && x8 && ~x4 && ~x1 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x70 && x11 && ~x10 && ~x6 && ~x8 )
						nx_state = s1;
					else if( ~x70 && ~x11 && x10 && x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x70 && ~x11 && x10 && ~x2 )
						nx_state = s1;
					else if( ~x70 && ~x11 && ~x10 && x12 && x9 )
						nx_state = s1;
					else if( ~x70 && ~x11 && ~x10 && x12 && ~x9 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x70 && ~x11 && ~x10 && ~x12 && x6 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x70 && ~x11 && ~x10 && ~x12 && ~x6 && x9 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x70 && ~x11 && ~x10 && ~x12 && ~x6 && ~x9 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else nx_state = s204;
				s205 : if( x64 && x61 && x8 && x53 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x64 && x61 && x8 && ~x53 && x37 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( x64 && x61 && x8 && ~x53 && ~x37 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x64 && x61 && ~x8 && x51 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x64 && x61 && ~x8 && ~x51 && x37 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( x64 && x61 && ~x8 && ~x51 && ~x37 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x64 && ~x61 && x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( x64 && ~x61 && ~x10 && x11 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s205;
						end
					else if( x64 && ~x61 && ~x10 && ~x11 && x12 && x8 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x64 && ~x61 && ~x10 && ~x11 && x12 && ~x8 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s933;
						end
					else if( x64 && ~x61 && ~x10 && ~x11 && ~x12 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s935;
						end
					else if( ~x64 && x14 && x8 && x30 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x64 && x14 && x8 && ~x30 && x37 )
						nx_state = s1;
					else if( ~x64 && x14 && x8 && ~x30 && ~x37 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x64 && x14 && ~x8 && x41 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x64 && x14 && ~x8 && ~x41 && x37 )
						nx_state = s1;
					else if( ~x64 && x14 && ~x8 && ~x41 && ~x37 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x64 && ~x14 && x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x64 && ~x14 && ~x10 && x11 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x64 && ~x14 && ~x10 && ~x11 && x12 && x8 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x64 && ~x14 && ~x10 && ~x11 && x12 && ~x8 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s933;
						end
					else if( ~x64 && ~x14 && ~x10 && ~x11 && ~x12 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s935;
						end
					else nx_state = s205;
				s206 : if( x64 && x61 && x29 && x50 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s933;
						end
					else if( x64 && x61 && x29 && ~x50 )
						nx_state = s206;
					else if( x64 && x61 && ~x29 && x60 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( x64 && x61 && ~x29 && ~x60 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x64 && ~x61 && x11 && x6 && x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s201;
						end
					else if( x64 && ~x61 && x11 && x6 && ~x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s759;
						end
					else if( x64 && ~x61 && x11 && ~x6 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s205;
						end
					else if( x64 && ~x61 && ~x11 && x8 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x64 && ~x61 && ~x11 && ~x8 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s593;
						end
					else if( ~x64 && x14 && x29 && x42 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s933;
						end
					else if( ~x64 && x14 && x29 && ~x42 )
						nx_state = s206;
					else if( ~x64 && x14 && ~x29 && x15 )
						nx_state = s1;
					else if( ~x64 && x14 && ~x29 && ~x15 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x64 && ~x14 && x11 && x6 && x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s201;
						end
					else if( ~x64 && ~x14 && x11 && x6 && ~x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s759;
						end
					else if( ~x64 && ~x14 && x11 && ~x6 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x64 && ~x14 && ~x11 && x8 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x64 && ~x14 && ~x11 && ~x8 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s593;
						end
					else nx_state = s206;
				s207 : if( x44 && x3 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x44 && ~x3 && x2 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x44 && ~x3 && ~x2 && x28 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x44 && ~x3 && ~x2 && ~x28 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x44 && x11 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x44 && ~x11 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x44 && ~x11 && ~x5 && x1 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x44 && ~x11 && ~x5 && ~x1 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else nx_state = s207;
				s208 : if( x69 && x70 && x64 && x63 && x21 && x20 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s936;
						end
					else if( x69 && x70 && x64 && x63 && x21 && ~x20 )
						begin
							y22 = 1'b1;	
							nx_state = s39;
						end
					else if( x69 && x70 && x64 && x63 && ~x21 && x20 )
						begin
							y54 = 1'b1;	
							nx_state = s525;
						end
					else if( x69 && x70 && x64 && x63 && ~x21 && ~x20 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s936;
						end
					else if( x69 && x70 && x64 && ~x63 && x65 && x67 && x21 )
						begin
							y5 = 1'b1;	
							nx_state = s937;
						end
					else if( x69 && x70 && x64 && ~x63 && x65 && x67 && ~x21 && x20 )
						begin
							y5 = 1'b1;	
							nx_state = s937;
						end
					else if( x69 && x70 && x64 && ~x63 && x65 && x67 && ~x21 && ~x20 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x69 && x70 && x64 && ~x63 && x65 && ~x67 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x63 && ~x65 && x66 )
						nx_state = s1;
					else if( x69 && x70 && x64 && ~x63 && ~x65 && ~x66 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s938;
						end
					else if( x69 && x70 && ~x64 && x63 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && x23 && x10 && x11 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && x23 && x10 && ~x11 && x12 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && x23 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && x23 && ~x10 )
						nx_state = s1;
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && x9 && x10 && x11 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && x9 && x10 && ~x11 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && x9 && ~x10 && x13 && x14 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && x9 && ~x10 && x13 && ~x14 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && x9 && ~x10 && x13 && ~x14 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && x9 && ~x10 && x13 && ~x14 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && x9 && ~x10 && x13 && ~x14 && ~x20 )
						nx_state = s1;
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && x9 && ~x10 && ~x13 && x15 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && x9 && ~x10 && ~x13 && ~x15 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && x9 && ~x10 && ~x13 && ~x15 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && x9 && ~x10 && ~x13 && ~x15 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && x9 && ~x10 && ~x13 && ~x15 && ~x20 )
						nx_state = s1;
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && ~x9 && x16 && x17 && x18 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && ~x9 && x16 && x17 && ~x18 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && ~x9 && x16 && x17 && ~x18 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && ~x9 && x16 && x17 && ~x18 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && ~x9 && x16 && x17 && ~x18 && ~x20 )
						nx_state = s1;
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && ~x9 && x16 && ~x17 && x19 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && ~x9 && x16 && ~x17 && ~x19 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && ~x9 && x16 && ~x17 && ~x19 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && ~x9 && x16 && ~x17 && ~x19 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && ~x9 && x16 && ~x17 && ~x19 && ~x20 )
						nx_state = s1;
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && x7 && ~x9 && ~x16 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && x24 && ~x23 && ~x7 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && ~x24 && x7 && x23 )
						begin
							y31 = 1'b1;	
							nx_state = s164;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && ~x24 && x7 && ~x23 && x9 && x10 && x8 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && ~x24 && x7 && ~x23 && x9 && x10 && ~x8 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && ~x24 && x7 && ~x23 && x9 && ~x10 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && ~x24 && x7 && ~x23 && x9 && ~x10 && ~x8 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && ~x24 && x7 && ~x23 && ~x9 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && ~x24 && x7 && ~x23 && ~x9 && x8 && ~x10 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && ~x24 && x7 && ~x23 && ~x9 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s98;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && x67 && ~x24 && ~x7 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && ~x67 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && ~x67 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x64 && ~x63 && x66 && ~x67 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x69 && x70 && ~x64 && ~x63 && x66 && ~x67 && ~x23 )
						nx_state = s1;
					else if( x69 && x70 && ~x64 && ~x63 && ~x66 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x70 && ~x64 && ~x63 && ~x66 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x70 && ~x64 && ~x63 && ~x66 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x69 && x70 && ~x64 && ~x63 && ~x66 && ~x15 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && x61 && x60 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x66 && x65 && x61 && x60 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x70 && x66 && x65 && x61 && x60 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x66 && x65 && x61 && x60 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x69 && ~x70 && x66 && x65 && x61 && ~x60 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x66 && x65 && x61 && ~x60 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x70 && x66 && x65 && x61 && ~x60 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && x61 && ~x60 && x62 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && x65 && x61 && ~x60 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x66 && x65 && x61 && ~x60 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x66 && x65 && x61 && ~x60 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( x69 && ~x70 && x66 && x65 && x61 && ~x60 && ~x62 && ~x18 )
						nx_state = s118;
					else if( x69 && ~x70 && x66 && x65 && ~x61 && x60 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x61 && x60 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x61 && x60 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( x69 && ~x70 && x66 && x65 && ~x61 && x60 && ~x18 )
						nx_state = s118;
					else if( x69 && ~x70 && x66 && x65 && ~x61 && ~x60 && x62 && x11 && x10 && x15 )
						nx_state = s47;
					else if( x69 && ~x70 && x66 && x65 && ~x61 && ~x60 && x62 && x11 && x10 && ~x15 && x7 )
						nx_state = s47;
					else if( x69 && ~x70 && x66 && x65 && ~x61 && ~x60 && x62 && x11 && x10 && ~x15 && ~x7 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x61 && ~x60 && x62 && x11 && ~x10 )
						nx_state = s47;
					else if( x69 && ~x70 && x66 && x65 && ~x61 && ~x60 && x62 && ~x11 && x12 && x9 && x15 )
						nx_state = s47;
					else if( x69 && ~x70 && x66 && x65 && ~x61 && ~x60 && x62 && ~x11 && x12 && x9 && ~x15 && x7 )
						nx_state = s47;
					else if( x69 && ~x70 && x66 && x65 && ~x61 && ~x60 && x62 && ~x11 && x12 && x9 && ~x15 && ~x7 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x61 && ~x60 && x62 && ~x11 && x12 && ~x9 )
						nx_state = s47;
					else if( x69 && ~x70 && x66 && x65 && ~x61 && ~x60 && x62 && ~x11 && ~x12 && x8 && x15 )
						nx_state = s47;
					else if( x69 && ~x70 && x66 && x65 && ~x61 && ~x60 && x62 && ~x11 && ~x12 && x8 && ~x15 && x7 )
						nx_state = s47;
					else if( x69 && ~x70 && x66 && x65 && ~x61 && ~x60 && x62 && ~x11 && ~x12 && x8 && ~x15 && ~x7 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x69 && ~x70 && x66 && x65 && ~x61 && ~x60 && x62 && ~x11 && ~x12 && ~x8 )
						nx_state = s47;
					else if( x69 && ~x70 && x66 && x65 && ~x61 && ~x60 && ~x62 )
						nx_state = s47;
					else if( x69 && ~x70 && x66 && ~x65 && x67 && x62 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s298;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && x67 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && x21 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x23 && x22 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x23 && x22 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x23 && x22 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x23 && x22 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x23 && ~x22 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x23 && ~x22 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x23 && ~x22 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && x23 && ~x22 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x23 && x22 && x18 && x14 )
						nx_state = s47;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x23 && x22 && x18 && ~x14 && x13 )
						nx_state = s47;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x23 && x22 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x23 && x22 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && x66 && ~x65 && ~x67 && ~x21 && ~x23 && ~x22 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x70 && ~x66 && x65 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && x65 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && x26 && x11 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s300;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && x26 && ~x11 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && x26 && ~x11 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && x26 && ~x11 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && x26 && ~x11 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && ~x26 && x19 && x16 && x11 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s368;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && ~x26 && x19 && x16 && x11 && ~x12 && x13 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && ~x26 && x19 && x16 && x11 && ~x12 && ~x13 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && ~x26 && x19 && x16 && ~x11 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s300;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && ~x26 && x19 && ~x16 && x17 && x11 && x13 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && ~x26 && x19 && ~x16 && x17 && x11 && ~x13 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s122;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && ~x26 && x19 && ~x16 && x17 && ~x11 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && ~x26 && x19 && ~x16 && ~x17 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && x24 && ~x26 && ~x19 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && x25 && x19 && ~x14 && ~x13 && x26 )
						nx_state = s208;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && x25 && x19 && ~x14 && ~x13 && ~x26 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && x25 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && x10 && x12 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && x10 && x12 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && x10 && x12 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && x10 && x12 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && x10 && ~x12 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s304;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && ~x10 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && ~x10 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && ~x10 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && ~x10 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && x10 && x12 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && x10 && x12 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && x10 && x12 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && x10 && x12 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && x10 && ~x12 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && ~x10 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && ~x10 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && ~x10 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && ~x10 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && x21 && x9 && x3 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && x21 && x9 && ~x3 && x4 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && x21 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && x21 && ~x9 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x66 && ~x65 && ~x67 && ~x21 )
						nx_state = s1;
					else if( ~x69 && x44 && x35 )
						nx_state = s1;
					else if( ~x69 && x44 && ~x35 && x13 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && x44 && ~x35 && ~x13 )
						begin
							y8 = 1'b1;	y17 = 1'b1;	
							nx_state = s408;
						end
					else if( ~x69 && ~x44 && x11 )
						nx_state = s1;
					else if( ~x69 && ~x44 && ~x11 && x1 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && ~x44 && ~x11 && ~x1 )
						begin
							y8 = 1'b1;	y17 = 1'b1;	
							nx_state = s408;
						end
					else nx_state = s208;
				s209 : if( x69 && x21 && x20 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( x69 && x21 && ~x20 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x21 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && x70 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x3 && x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x69 && ~x70 && x3 && ~x4 )
						nx_state = s209;
					else if( ~x69 && ~x70 && ~x3 )
						nx_state = s1;
					else nx_state = s209;
				s210 : if( x69 && x62 && x17 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							nx_state = s939;
						end
					else if( x69 && x62 && ~x17 )
						begin
							y1 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s940;
						end
					else if( x69 && ~x62 && x63 && x64 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x69 && ~x62 && x63 && x64 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x69 && ~x62 && x63 && x64 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x62 && x63 && x64 && ~x22 )
						nx_state = s1;
					else if( x69 && ~x62 && x63 && ~x64 && x66 && x7 && x31 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && ~x62 && x63 && ~x64 && x66 && x7 && ~x31 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x69 && ~x62 && x63 && ~x64 && x66 && ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x62 && x63 && ~x64 && ~x66 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x69 && ~x62 && x63 && ~x64 && ~x66 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x69 && ~x62 && x63 && ~x64 && ~x66 && x19 && ~x14 && ~x13 && x11 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( x69 && ~x62 && x63 && ~x64 && ~x66 && x19 && ~x14 && ~x13 && x11 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( x69 && ~x62 && x63 && ~x64 && ~x66 && x19 && ~x14 && ~x13 && ~x11 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( x69 && ~x62 && x63 && ~x64 && ~x66 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x62 && ~x63 && x64 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x62 && ~x63 && x64 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x62 && ~x63 && x64 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x69 && ~x62 && ~x63 && x64 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x62 && ~x63 && ~x64 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x62 && ~x63 && ~x64 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x62 && ~x63 && ~x64 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x69 && ~x62 && ~x63 && ~x64 && ~x23 )
						nx_state = s1;
					else if( ~x69 && x70 && x15 && x62 && x16 )
						begin
							y13 = 1'b1;	
							nx_state = s450;
						end
					else if( ~x69 && x70 && x15 && x62 && ~x16 && x11 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s436;
						end
					else if( ~x69 && x70 && x15 && x62 && ~x16 && ~x11 && x10 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s448;
						end
					else if( ~x69 && x70 && x15 && x62 && ~x16 && ~x11 && ~x10 )
						nx_state = s210;
					else if( ~x69 && x70 && x15 && ~x62 && x63 && x64 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x69 && x70 && x15 && ~x62 && x63 && ~x64 && x33 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && x70 && x15 && ~x62 && x63 && ~x64 && ~x33 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && x70 && x15 && ~x62 && x63 && ~x64 && ~x33 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && x70 && x15 && ~x62 && ~x63 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x69 && x70 && ~x15 && x62 && x16 && x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s451;
						end
					else if( ~x69 && x70 && ~x15 && x62 && x16 && ~x3 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s927;
						end
					else if( ~x69 && x70 && ~x15 && x62 && ~x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && x47 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && x47 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && x64 && ~x47 )
						begin
							y21 = 1'b1;	y27 = 1'b1;	
							nx_state = s930;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && ~x64 && x49 )
						begin
							y12 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s912;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && x63 && ~x64 && ~x49 )
						nx_state = s210;
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && x16 && x64 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && x16 && x64 && ~x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && x16 && ~x64 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && x16 && ~x64 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && x70 && ~x15 && ~x62 && ~x63 && ~x16 )
						begin
							y21 = 1'b1;	y27 = 1'b1;	
							nx_state = s930;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x46 && x8 && x26 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x46 && x8 && ~x26 && x37 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x44 && x45 && x46 && x8 && ~x26 && ~x37 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x46 && ~x8 && x40 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x46 && ~x8 && ~x40 && x37 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x44 && x45 && x46 && ~x8 && ~x40 && ~x37 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x46 && x11 && x6 && x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x46 && x11 && x6 && ~x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x46 && x11 && ~x6 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s215;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x46 && ~x11 && x8 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x46 && ~x11 && ~x8 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s320;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x20 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x20 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x20 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && ~x70 && ~x44 && x46 && x10 && x11 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x69 && ~x70 && ~x44 && x46 && x10 && ~x11 && x7 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x44 && x46 && x10 && ~x11 && ~x7 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x69 && ~x70 && ~x44 && x46 && ~x10 && x13 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x69 && ~x70 && ~x44 && x46 && ~x10 && ~x13 && x7 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x44 && x46 && ~x10 && ~x13 && ~x7 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x46 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x46 && ~x5 && x6 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x46 && ~x5 && ~x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else nx_state = s210;
				s211 : if( x46 && x45 && x12 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x46 && x45 && ~x12 )
						nx_state = s211;
					else if( x46 && ~x45 && x4 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x46 && ~x45 && ~x4 )
						nx_state = s211;
					else if( ~x46 && x45 && x12 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x46 && x45 && ~x12 && x4 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x46 && x45 && ~x12 && ~x4 )
						nx_state = s211;
					else if( ~x46 && ~x45 && x10 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x46 && ~x45 && ~x10 && x4 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x46 && ~x45 && ~x10 && ~x4 )
						nx_state = s211;
					else nx_state = s211;
				s212 : if( x46 && x45 && x13 && x6 && x16 && x10 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x46 && x45 && x13 && x6 && x16 && ~x10 )
						nx_state = s212;
					else if( x46 && x45 && x13 && x6 && ~x16 && x10 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x46 && x45 && x13 && x6 && ~x16 && ~x10 )
						nx_state = s212;
					else if( x46 && x45 && x13 && ~x6 )
						nx_state = s1;
					else if( x46 && x45 && ~x13 && x15 && x10 && x4 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x46 && x45 && ~x13 && x15 && x10 && ~x4 )
						nx_state = s212;
					else if( x46 && x45 && ~x13 && x15 && ~x10 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x46 && x45 && ~x13 && x15 && ~x10 && ~x4 )
						nx_state = s212;
					else if( x46 && x45 && ~x13 && ~x15 )
						nx_state = s1;
					else if( x46 && ~x45 && x47 && x8 && x4 && x3 && x7 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x46 && ~x45 && x47 && x8 && x4 && x3 && ~x7 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( x46 && ~x45 && x47 && x8 && x4 && ~x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x46 && ~x45 && x47 && x8 && ~x4 )
						nx_state = s212;
					else if( x46 && ~x45 && x47 && ~x8 )
						nx_state = s1;
					else if( x46 && ~x45 && ~x47 && x4 && x9 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x46 && ~x45 && ~x47 && x4 && ~x9 && x10 && x11 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x46 && ~x45 && ~x47 && x4 && ~x9 && x10 && ~x11 && x3 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( x46 && ~x45 && ~x47 && x4 && ~x9 && x10 && ~x11 && ~x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x46 && ~x45 && ~x47 && x4 && ~x9 && ~x10 && x3 && x11 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x46 && ~x45 && ~x47 && x4 && ~x9 && ~x10 && x3 && ~x11 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s177;
						end
					else if( x46 && ~x45 && ~x47 && x4 && ~x9 && ~x10 && ~x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x46 && ~x45 && ~x47 && ~x4 )
						nx_state = s212;
					else if( ~x46 && x45 && x12 )
						nx_state = s1;
					else if( ~x46 && x45 && ~x12 && x4 && x9 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x46 && x45 && ~x12 && x4 && ~x9 && x10 && x11 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x46 && x45 && ~x12 && x4 && ~x9 && x10 && ~x11 && x3 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( ~x46 && x45 && ~x12 && x4 && ~x9 && x10 && ~x11 && ~x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x46 && x45 && ~x12 && x4 && ~x9 && ~x10 && x3 && x11 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x46 && x45 && ~x12 && x4 && ~x9 && ~x10 && x3 && ~x11 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s177;
						end
					else if( ~x46 && x45 && ~x12 && x4 && ~x9 && ~x10 && ~x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x46 && x45 && ~x12 && ~x4 )
						nx_state = s212;
					else if( ~x46 && ~x45 && x10 && x11 && x4 && x13 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x46 && ~x45 && x10 && x11 && x4 && ~x13 && x3 && x12 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( ~x46 && ~x45 && x10 && x11 && x4 && ~x13 && x3 && ~x12 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s177;
						end
					else if( ~x46 && ~x45 && x10 && x11 && x4 && ~x13 && ~x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x46 && ~x45 && x10 && x11 && ~x4 )
						nx_state = s212;
					else if( ~x46 && ~x45 && x10 && ~x11 )
						nx_state = s1;
					else if( ~x46 && ~x45 && ~x10 && x12 && x4 && x11 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x46 && ~x45 && ~x10 && x12 && x4 && ~x11 && x3 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x46 && ~x45 && ~x10 && x12 && x4 && ~x11 && ~x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x46 && ~x45 && ~x10 && x12 && ~x4 )
						nx_state = s212;
					else if( ~x46 && ~x45 && ~x10 && ~x12 )
						nx_state = s1;
					else nx_state = s212;
				s213 : if( x45 && x16 && x1 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s578;
						end
					else if( x45 && x16 && ~x1 )
						nx_state = s213;
					else if( x45 && ~x16 && x1 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x45 && ~x16 && ~x1 )
						nx_state = s213;
					else if( ~x45 && x6 && x2 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s578;
						end
					else if( ~x45 && x6 && ~x2 )
						nx_state = s213;
					else if( ~x45 && ~x6 && x2 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x45 && ~x6 && ~x2 )
						nx_state = s213;
					else nx_state = s213;
				s214 : if( x46 && x2 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x46 && ~x2 )
						nx_state = s214;
					else if( ~x46 && x10 && x2 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x46 && x10 && ~x2 )
						nx_state = s214;
					else if( ~x46 && ~x10 && x45 && x2 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x46 && ~x10 && x45 && ~x2 )
						nx_state = s214;
					else if( ~x46 && ~x10 && ~x45 && x3 )
						nx_state = s1;
					else if( ~x46 && ~x10 && ~x45 && ~x3 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s212;
						end
					else nx_state = s214;
				s215 : if( x69 && x17 && x18 && x5 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && x17 && x18 && ~x5 && x6 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && x17 && x18 && ~x5 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && x17 && ~x18 && x14 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x69 && x17 && ~x18 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x17 && x6 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s320;
						end
					else if( x69 && ~x17 && ~x6 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s280;
						end
					else if( ~x69 && x70 && x61 && x12 && x27 && x33 )
						begin
							y10 = 1'b1;	
							nx_state = s841;
						end
					else if( ~x69 && x70 && x61 && x12 && x27 && ~x33 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( ~x69 && x70 && x61 && x12 && x27 && ~x33 && ~x13 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s840;
						end
					else if( ~x69 && x70 && x61 && x12 && ~x27 && x29 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s874;
						end
					else if( ~x69 && x70 && x61 && x12 && ~x27 && x29 && ~x1 && x9 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x69 && x70 && x61 && x12 && ~x27 && x29 && ~x1 && x9 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s875;
						end
					else if( ~x69 && x70 && x61 && x12 && ~x27 && x29 && ~x1 && ~x9 )
						nx_state = s215;
					else if( ~x69 && x70 && x61 && x12 && ~x27 && ~x29 )
						nx_state = s215;
					else if( ~x69 && x70 && x61 && ~x12 && x29 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s320;
						end
					else if( ~x69 && x70 && x61 && ~x12 && ~x29 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s842;
						end
					else if( ~x69 && x70 && ~x61 && x17 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s913;
						end
					else if( ~x69 && x70 && ~x61 && ~x17 && x57 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s733;
						end
					else if( ~x69 && x70 && ~x61 && ~x17 && ~x57 )
						nx_state = s215;
					else if( ~x69 && ~x70 && x44 && x6 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s320;
						end
					else if( ~x69 && ~x70 && x44 && ~x6 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s280;
						end
					else if( ~x69 && ~x70 && ~x44 && x10 && x6 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s320;
						end
					else if( ~x69 && ~x70 && ~x44 && x10 && ~x6 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s280;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 )
						nx_state = s215;
					else nx_state = s215;
				s216 : if( x70 && x62 && x26 && x28 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( x70 && x62 && x26 && x28 && ~x1 && x2 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s941;
						end
					else if( x70 && x62 && x26 && x28 && ~x1 && ~x2 && x25 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s941;
						end
					else if( x70 && x62 && x26 && x28 && ~x1 && ~x2 && ~x25 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( x70 && x62 && x26 && ~x28 && x1 && x2 && x3 && x25 )
						nx_state = s216;
					else if( x70 && x62 && x26 && ~x28 && x1 && x2 && x3 && ~x25 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( x70 && x62 && x26 && ~x28 && x1 && x2 && ~x3 && x4 && x5 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s942;
						end
					else if( x70 && x62 && x26 && ~x28 && x1 && x2 && ~x3 && x4 && ~x5 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( x70 && x62 && x26 && ~x28 && x1 && x2 && ~x3 && ~x4 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( x70 && x62 && x26 && ~x28 && x1 && ~x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s943;
						end
					else if( x70 && x62 && x26 && ~x28 && ~x1 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s941;
						end
					else if( x70 && x62 && ~x26 && x27 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s943;
						end
					else if( x70 && x62 && ~x26 && ~x27 && x28 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( x70 && x62 && ~x26 && ~x27 && x28 && ~x1 && x4 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s941;
						end
					else if( x70 && x62 && ~x26 && ~x27 && x28 && ~x1 && ~x4 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( x70 && x62 && ~x26 && ~x27 && ~x28 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s943;
						end
					else if( x70 && ~x62 && x26 && x28 && x64 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( x70 && ~x62 && x26 && x28 && x64 && ~x1 && x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( x70 && ~x62 && x26 && x28 && x64 && ~x1 && ~x2 && x25 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( x70 && ~x62 && x26 && x28 && x64 && ~x1 && ~x2 && ~x25 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( x70 && ~x62 && x26 && x28 && ~x64 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s944;
						end
					else if( x70 && ~x62 && x26 && x28 && ~x64 && ~x37 && x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( x70 && ~x62 && x26 && x28 && ~x64 && ~x37 && ~x2 && x25 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( x70 && ~x62 && x26 && x28 && ~x64 && ~x37 && ~x2 && ~x25 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( x70 && ~x62 && x26 && ~x28 && x64 && x1 && x2 && x3 && x25 )
						nx_state = s216;
					else if( x70 && ~x62 && x26 && ~x28 && x64 && x1 && x2 && x3 && ~x25 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( x70 && ~x62 && x26 && ~x28 && x64 && x1 && x2 && ~x3 && x4 && x5 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else if( x70 && ~x62 && x26 && ~x28 && x64 && x1 && x2 && ~x3 && x4 && ~x5 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( x70 && ~x62 && x26 && ~x28 && x64 && x1 && x2 && ~x3 && ~x4 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( x70 && ~x62 && x26 && ~x28 && x64 && x1 && ~x2 )
						begin
							y11 = 1'b1;	
							nx_state = s247;
						end
					else if( x70 && ~x62 && x26 && ~x28 && x64 && ~x1 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( x70 && ~x62 && x26 && ~x28 && ~x64 && x37 && x32 && x3 && x25 )
						nx_state = s216;
					else if( x70 && ~x62 && x26 && ~x28 && ~x64 && x37 && x32 && x3 && ~x25 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( x70 && ~x62 && x26 && ~x28 && ~x64 && x37 && x32 && ~x3 && x4 && x5 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else if( x70 && ~x62 && x26 && ~x28 && ~x64 && x37 && x32 && ~x3 && x4 && ~x5 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s917;
						end
					else if( x70 && ~x62 && x26 && ~x28 && ~x64 && x37 && x32 && ~x3 && ~x4 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s944;
						end
					else if( x70 && ~x62 && x26 && ~x28 && ~x64 && x37 && ~x32 )
						begin
							y11 = 1'b1;	
							nx_state = s247;
						end
					else if( x70 && ~x62 && x26 && ~x28 && ~x64 && ~x37 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( x70 && ~x62 && ~x26 && x27 )
						begin
							y11 = 1'b1;	
							nx_state = s247;
						end
					else if( x70 && ~x62 && ~x26 && ~x27 && x28 && x1 && x64 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( x70 && ~x62 && ~x26 && ~x27 && x28 && x1 && ~x64 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s944;
						end
					else if( x70 && ~x62 && ~x26 && ~x27 && x28 && ~x1 && x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( x70 && ~x62 && ~x26 && ~x27 && x28 && ~x1 && ~x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( x70 && ~x62 && ~x26 && ~x27 && ~x28 )
						begin
							y11 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x70 && x3 && x5 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s733;
						end
					else if( ~x70 && x3 && ~x5 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x70 && ~x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else nx_state = s216;
				s217 : if( x69 && x65 && x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x65 && x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && x65 && x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x69 && x65 && x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && x65 && x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && x65 && x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && x65 && x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( x69 && x65 && ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x65 && ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x65 && ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && x65 && ~x21 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x65 && x66 && x21 )
						nx_state = s1;
					else if( x69 && ~x65 && x66 && ~x21 && x22 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( x69 && ~x65 && x66 && ~x21 && x22 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( x69 && ~x65 && x66 && ~x21 && x22 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x65 && x66 && ~x21 && x22 && x23 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x65 && x66 && ~x21 && x22 && ~x23 && x19 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s608;
						end
					else if( x69 && ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && x20 && x15 && x10 && x11 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s4;
						end
					else if( x69 && ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && x20 && x15 && x10 && ~x11 && x12 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s4;
						end
					else if( x69 && ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && x20 && x15 && x10 && ~x11 && ~x12 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && x20 && x15 && ~x10 && x12 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( x69 && ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && x20 && x15 && ~x10 && x12 && ~x11 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && x20 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( x69 && ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && x20 && ~x15 && x16 && x10 && x12 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && x20 && ~x15 && x16 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s365;
						end
					else if( x69 && ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && x20 && ~x15 && x16 && ~x10 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && x20 && ~x15 && ~x16 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s151;
						end
					else if( x69 && ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && ~x20 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && x23 && x3 )
						begin
							y3 = 1'b1;	
							nx_state = s835;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && x23 && ~x3 && x18 && x15 && x7 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s151;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && x23 && ~x3 && x18 && x15 && ~x7 && x9 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && x23 && ~x3 && x18 && x15 && ~x7 && ~x9 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && x23 && ~x3 && x18 && ~x15 && x7 && x9 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s274;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && x23 && ~x3 && x18 && ~x15 && x7 && ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && x23 && ~x3 && x18 && ~x15 && ~x7 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s274;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && x23 && ~x3 && ~x18 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && ~x23 && x15 && x7 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s151;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && ~x23 && x15 && ~x7 && x9 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s361;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && ~x23 && x15 && ~x7 && ~x9 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && ~x23 && ~x15 && x7 && x9 )
						begin
							y3 = 1'b1;	
							nx_state = s835;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && ~x23 && ~x15 && x7 && ~x9 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s275;
						end
					else if( x69 && ~x65 && x66 && ~x21 && ~x22 && ~x23 && ~x15 && ~x7 )
						begin
							y3 = 1'b1;	
							nx_state = s835;
						end
					else if( x69 && ~x65 && ~x66 && x24 && x26 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x69 && ~x65 && ~x66 && x24 && x26 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x69 && ~x65 && ~x66 && x24 && x26 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x66 && x24 && x26 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x66 && x24 && ~x26 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( x69 && ~x65 && ~x66 && ~x24 && x25 && x26 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x65 && ~x66 && ~x24 && x25 && x26 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x65 && ~x66 && ~x24 && x25 && x26 && x19 && ~x14 && ~x13 )
						nx_state = s217;
					else if( x69 && ~x65 && ~x66 && ~x24 && x25 && x26 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x66 && ~x24 && x25 && ~x26 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x65 && ~x66 && ~x24 && ~x25 && x26 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x65 && ~x66 && ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x65 && ~x66 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x69 && ~x65 && ~x66 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x65 && ~x66 && ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else if( ~x69 && x10 && x9 )
						nx_state = s1;
					else if( ~x69 && x10 && ~x9 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x69 && ~x10 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( ~x69 && ~x10 && ~x6 && x8 && x4 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s320;
						end
					else if( ~x69 && ~x10 && ~x6 && x8 && ~x4 && x1 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x69 && ~x10 && ~x6 && x8 && ~x4 && x1 && ~x3 )
						begin
							y5 = 1'b1;	y13 = 1'b1;	
							nx_state = s740;
						end
					else if( ~x69 && ~x10 && ~x6 && x8 && ~x4 && ~x1 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s738;
						end
					else if( ~x69 && ~x10 && ~x6 && ~x8 )
						nx_state = s1;
					else nx_state = s217;
				s218 : if( 1'b1 )
						begin
							y5 = 1'b1;	
							nx_state = s945;
						end
					else nx_state = s218;
				s219 : if( 1'b1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y9 = 1'b1;	
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s946;
						end
					else nx_state = s219;
				s220 : if( x70 && x63 && x13 )
						begin
							y7 = 1'b1;	
							nx_state = s891;
						end
					else if( x70 && x63 && ~x13 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x70 && x63 && ~x13 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x70 && x63 && ~x13 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && x63 && ~x13 && ~x14 )
						nx_state = s1;
					else if( x70 && ~x63 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x70 && ~x63 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x70 && ~x63 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x8 )
						nx_state = s1;
					else if( ~x70 && x21 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x21 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x21 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x9 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x22 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x70 && ~x21 && x22 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x70 && ~x21 && x22 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x22 && ~x7 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x70 && ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x70 && ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s220;
				s221 : if( x70 && x62 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							y8 = 1'b1;	
							nx_state = s219;
						end
					else if( x70 && ~x62 && x63 && x31 && x30 && x8 )
						begin
							y42 = 1'b1;	
							nx_state = s754;
						end
					else if( x70 && ~x62 && x63 && x31 && x30 && ~x8 )
						begin
							y40 = 1'b1;	
							nx_state = s947;
						end
					else if( x70 && ~x62 && x63 && x31 && ~x30 && x7 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x70 && ~x62 && x63 && x31 && ~x30 && ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && x63 && ~x31 && x7 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x70 && ~x62 && x63 && ~x31 && ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && x65 && x28 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x65 && x28 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x65 && x28 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && x65 && x28 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && x65 && ~x28 )
						begin
							y8 = 1'b1;	
							nx_state = s783;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x65 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x65 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x65 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x65 && ~x8 )
						nx_state = s1;
					else if( ~x70 && x65 && x21 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( ~x70 && x65 && x21 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( ~x70 && x65 && x21 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x70 && x65 && x21 && ~x8 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && x23 && x22 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && x23 && x22 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && x23 && x22 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && x23 && x22 && ~x8 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && x23 && ~x22 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && x23 && ~x22 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && x23 && ~x22 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && x23 && ~x22 && ~x9 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && ~x23 && x8 && x22 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && x8 && x22 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && x8 && x22 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && ~x23 && x8 && ~x22 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && x8 && ~x22 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && x8 && ~x22 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && ~x23 && ~x8 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && ~x65 && x66 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && ~x65 && x66 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && x62 && ~x61 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x65 && x66 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && ~x65 && x66 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x65 && x66 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && ~x65 && x66 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && x66 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x65 && x66 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && x66 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x65 && x66 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && x21 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x21 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else nx_state = s221;
				s222 : if( x65 && x70 && x62 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x65 && x70 && x62 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x65 && x70 && x62 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( x65 && x70 && x62 && ~x27 )
						nx_state = s1;
					else if( x65 && x70 && ~x62 && x63 && x66 && x7 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x65 && x70 && ~x62 && x63 && x66 && ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && x70 && ~x62 && x63 && ~x66 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s656;
						end
					else if( x65 && x70 && ~x62 && ~x63 && x66 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x65 && x70 && ~x62 && ~x63 && x66 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x65 && x70 && ~x62 && ~x63 && x66 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && x70 && ~x62 && ~x63 && x66 && ~x14 )
						nx_state = s1;
					else if( x65 && x70 && ~x62 && ~x63 && ~x66 )
						begin
							y8 = 1'b1;	
							nx_state = s783;
						end
					else if( x65 && ~x70 && x66 && x68 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( x65 && ~x70 && x66 && ~x68 && x60 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x65 && ~x70 && x66 && ~x68 && ~x60 && x61 && x62 && x20 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	
							nx_state = s330;
						end
					else if( x65 && ~x70 && x66 && ~x68 && ~x60 && x61 && x62 && ~x20 && x16 && x11 && x12 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s278;
						end
					else if( x65 && ~x70 && x66 && ~x68 && ~x60 && x61 && x62 && ~x20 && x16 && x11 && ~x12 && x13 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s278;
						end
					else if( x65 && ~x70 && x66 && ~x68 && ~x60 && x61 && x62 && ~x20 && x16 && x11 && ~x12 && ~x13 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( x65 && ~x70 && x66 && ~x68 && ~x60 && x61 && x62 && ~x20 && x16 && ~x11 && x13 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s135;
						end
					else if( x65 && ~x70 && x66 && ~x68 && ~x60 && x61 && x62 && ~x20 && x16 && ~x11 && ~x13 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x65 && ~x70 && x66 && ~x68 && ~x60 && x61 && x62 && ~x20 && ~x16 && x17 && x11 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x65 && ~x70 && x66 && ~x68 && ~x60 && x61 && x62 && ~x20 && ~x16 && x17 && x11 && ~x13 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x65 && ~x70 && x66 && ~x68 && ~x60 && x61 && x62 && ~x20 && ~x16 && x17 && ~x11 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x65 && ~x70 && x66 && ~x68 && ~x60 && x61 && x62 && ~x20 && ~x16 && ~x17 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x65 && ~x70 && x66 && ~x68 && ~x60 && x61 && ~x62 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x65 && ~x70 && x66 && ~x68 && ~x60 && ~x61 )
						begin
							y2 = 1'b1;	y19 = 1'b1;	y24 = 1'b1;	
							nx_state = s837;
						end
					else if( x65 && ~x70 && ~x66 && x67 && x21 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x65 && ~x70 && ~x66 && x67 && x21 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x65 && ~x70 && ~x66 && x67 && x21 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x65 && ~x70 && ~x66 && x67 && x21 && ~x8 )
						nx_state = s1;
					else if( x65 && ~x70 && ~x66 && x67 && ~x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s111;
						end
					else if( x65 && ~x70 && ~x66 && ~x67 && x20 && x19 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && ~x70 && ~x66 && ~x67 && x20 && x19 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && ~x70 && ~x66 && ~x67 && x20 && x19 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x70 && ~x66 && ~x67 && x20 && x19 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x70 && ~x66 && ~x67 && x20 && ~x19 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	y25 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && ~x70 && ~x66 && ~x67 && ~x20 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	y25 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x65 && x70 && x62 && x17 && x18 && x5 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x65 && x70 && x62 && x17 && x18 && ~x5 && x6 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x65 && x70 && x62 && x17 && x18 && ~x5 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && x70 && x62 && x17 && ~x18 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( ~x65 && x70 && x62 && x17 && ~x18 && ~x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x65 && x70 && x62 && ~x17 && x18 && x1 )
						nx_state = s1;
					else if( ~x65 && x70 && x62 && ~x17 && x18 && ~x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x65 && x70 && x62 && ~x17 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && x63 && x9 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( ~x65 && x70 && ~x62 && x63 && ~x9 )
						nx_state = s222;
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && x5 && x18 && x19 && x12 )
						begin
							y54 = 1'b1;	
							nx_state = s525;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && x5 && x18 && x19 && ~x12 )
						begin
							y55 = 1'b1;	
							nx_state = s526;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && x5 && x18 && ~x19 && x12 && x6 )
						begin
							y16 = 1'b1;	y50 = 1'b1;	
							nx_state = s527;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && x5 && x18 && ~x19 && x12 && ~x6 && x16 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && x5 && x18 && ~x19 && x12 && ~x6 && ~x16 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && x5 && x18 && ~x19 && x12 && ~x6 && ~x16 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && x5 && x18 && ~x19 && x12 && ~x6 && ~x16 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && x5 && x18 && ~x19 && x12 && ~x6 && ~x16 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && x5 && x18 && ~x19 && ~x12 && x6 )
						begin
							y12 = 1'b1;	y48 = 1'b1;	
							nx_state = s529;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && x5 && x18 && ~x19 && ~x12 && ~x6 && x15 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && x5 && x18 && ~x19 && ~x12 && ~x6 && ~x15 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && x5 && x18 && ~x19 && ~x12 && ~x6 && ~x15 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && x5 && x18 && ~x19 && ~x12 && ~x6 && ~x15 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && x5 && x18 && ~x19 && ~x12 && ~x6 && ~x15 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && x5 && ~x18 && x19 )
						begin
							y27 = 1'b1;	y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s284;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && x5 && ~x18 && ~x19 && x6 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && x5 && ~x18 && ~x19 && ~x6 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && x19 && x6 && x12 && x11 )
						begin
							y46 = 1'b1;	
							nx_state = s531;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && x19 && x6 && x12 && ~x11 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && x19 && x6 && x12 && ~x11 && x9 && ~x10 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && x19 && x6 && x12 && ~x11 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && x19 && x6 && ~x12 && x10 )
						begin
							y46 = 1'b1;	
							nx_state = s531;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && x19 && x6 && ~x12 && ~x10 && x9 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && x19 && x6 && ~x12 && ~x10 && x9 && ~x11 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && x19 && x6 && ~x12 && ~x10 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && x19 && ~x6 && x12 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && x19 && ~x6 && ~x12 )
						begin
							y56 = 1'b1;	y57 = 1'b1;	
							nx_state = s284;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && ~x19 && x6 && x12 && x14 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && ~x19 && x6 && x12 && ~x14 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && ~x19 && x6 && x12 && ~x14 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && ~x19 && x6 && x12 && ~x14 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && ~x19 && x6 && x12 && ~x14 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && ~x19 && x6 && ~x12 && x13 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && ~x19 && x6 && ~x12 && ~x13 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && ~x19 && x6 && ~x12 && ~x13 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && ~x19 && x6 && ~x12 && ~x13 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && ~x19 && x6 && ~x12 && ~x13 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && x18 && ~x19 && ~x6 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && ~x18 && x19 && x12 && x6 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && ~x18 && x19 && x12 && ~x6 )
						begin
							y38 = 1'b1;	
							nx_state = s532;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && ~x18 && x19 && ~x12 && x6 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && ~x18 && x19 && ~x12 && ~x6 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && x8 && ~x5 && ~x18 && ~x19 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && x66 && ~x8 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x65 && x70 && ~x62 && ~x63 && ~x66 )
						begin
							y7 = 1'b1;	
							nx_state = s82;
						end
					else if( ~x65 && ~x70 && x67 && x68 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x65 && ~x70 && x67 && x68 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x65 && ~x70 && x67 && x68 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x67 && x68 && x21 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x67 && x68 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x70 && x67 && x68 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x70 && x67 && x68 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x67 && x68 && ~x21 && ~x20 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x67 && ~x68 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x65 && ~x70 && x67 && ~x68 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x65 && ~x70 && x67 && ~x68 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x67 && ~x68 && x62 && ~x61 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x67 && ~x68 && ~x62 && x63 && x17 && x13 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && ~x70 && x67 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && ~x70 && x67 && ~x68 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x67 && ~x68 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x67 && ~x68 && ~x62 && ~x63 && x64 && x4 )
						begin
							y31 = 1'b1;	
							nx_state = s164;
						end
					else if( ~x65 && ~x70 && x67 && ~x68 && ~x62 && ~x63 && x64 && ~x4 && x18 && x16 && x8 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x65 && ~x70 && x67 && ~x68 && ~x62 && ~x63 && x64 && ~x4 && x18 && x16 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x65 && ~x70 && x67 && ~x68 && ~x62 && ~x63 && x64 && ~x4 && x18 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s299;
						end
					else if( ~x65 && ~x70 && x67 && ~x68 && ~x62 && ~x63 && x64 && ~x4 && ~x18 )
						begin
							y14 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && ~x70 && x67 && ~x68 && ~x62 && ~x63 && ~x64 && x19 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x65 && ~x70 && x67 && ~x68 && ~x62 && ~x63 && ~x64 && x19 && ~x13 && x12 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x65 && ~x70 && x67 && ~x68 && ~x62 && ~x63 && ~x64 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x70 && x67 && ~x68 && ~x62 && ~x63 && ~x64 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x67 && x21 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( ~x65 && ~x70 && ~x67 && ~x21 && x23 && x22 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x65 && ~x70 && ~x67 && ~x21 && x23 && ~x22 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x65 && ~x70 && ~x67 && ~x21 && x23 && ~x22 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x65 && ~x70 && ~x67 && ~x21 && x23 && ~x22 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x67 && ~x21 && x23 && ~x22 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x70 && ~x67 && ~x21 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else nx_state = s222;
				s223 : if( x63 && x12 )
						begin
							y17 = 1'b1;	
							nx_state = s98;
						end
					else if( x63 && ~x12 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x63 && ~x12 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x63 && ~x12 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x63 && ~x12 && ~x1 )
						nx_state = s1;
					else if( ~x63 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s948;
						end
					else nx_state = s223;
				s224 : if( x21 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x21 && ~x20 )
						nx_state = s1;
					else nx_state = s224;
				s225 : if( x25 && x24 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x25 && ~x24 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x25 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else nx_state = s225;
				s226 : if( x21 && x20 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y22 = 1'b1;	
							y32 = 1'b1;	y33 = 1'b1;	
							nx_state = s949;
						end
					else if( x21 && ~x20 )
						begin
							y28 = 1'b1;	
							nx_state = s469;
						end
					else if( ~x21 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x21 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x21 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x21 && ~x10 )
						nx_state = s1;
					else nx_state = s226;
				s227 : if( x69 && x70 && x62 )
						begin
							y22 = 1'b1;	
							nx_state = s39;
						end
					else if( x69 && x70 && ~x62 && x63 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x21 && x20 )
						begin
							y16 = 1'b1;	
							nx_state = s293;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x21 && ~x20 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x21 && ~x20 && ~x12 && x17 && x16 && x19 && x11 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x21 && ~x20 && ~x12 && x17 && x16 && x19 && ~x11 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x21 && ~x20 && ~x12 && x17 && x16 && ~x19 && x18 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x21 && ~x20 && ~x12 && x17 && x16 && ~x19 && ~x18 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x21 && ~x20 && ~x12 && x17 && ~x16 && x11 )
						begin
							y3 = 1'b1;	
							nx_state = s788;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x21 && ~x20 && ~x12 && x17 && ~x16 && ~x11 )
						begin
							y32 = 1'b1;	
							nx_state = s854;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x21 && ~x20 && ~x12 && ~x17 && x16 && x19 && x14 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x21 && ~x20 && ~x12 && ~x17 && x16 && x19 && ~x14 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x21 && ~x20 && ~x12 && ~x17 && x16 && ~x19 && x13 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x21 && ~x20 && ~x12 && ~x17 && x16 && ~x19 && ~x13 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && x21 && ~x20 && ~x12 && ~x17 && ~x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x70 && ~x62 && ~x63 && x64 && ~x21 )
						begin
							y16 = 1'b1;	
							nx_state = s293;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && x23 && x10 && x11 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && x23 && x10 && ~x11 && x12 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && x23 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && x23 && ~x10 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && x9 && x10 && x11 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && x9 && x10 && ~x11 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && x9 && ~x10 && x13 && x14 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && x9 && ~x10 && x13 && ~x14 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && x9 && ~x10 && x13 && ~x14 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && x9 && ~x10 && x13 && ~x14 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && x9 && ~x10 && x13 && ~x14 && ~x20 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && x9 && ~x10 && ~x13 && x15 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && x9 && ~x10 && ~x13 && ~x15 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && x9 && ~x10 && ~x13 && ~x15 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && x9 && ~x10 && ~x13 && ~x15 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && x9 && ~x10 && ~x13 && ~x15 && ~x20 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && ~x9 && x16 && x17 && x18 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && ~x9 && x16 && x17 && ~x18 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && ~x9 && x16 && x17 && ~x18 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && ~x9 && x16 && x17 && ~x18 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && ~x9 && x16 && x17 && ~x18 && ~x20 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && ~x9 && x16 && ~x17 && x19 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && ~x9 && x16 && ~x17 && ~x19 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && ~x9 && x16 && ~x17 && ~x19 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && ~x9 && x16 && ~x17 && ~x19 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && ~x9 && x16 && ~x17 && ~x19 && ~x20 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && x7 && ~x9 && ~x16 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && x24 && ~x23 && ~x6 && ~x7 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && ~x24 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && ~x24 && ~x6 && x7 && x23 )
						begin
							y31 = 1'b1;	
							nx_state = s164;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && ~x24 && ~x6 && x7 && ~x23 && x9 && x10 && x8 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && ~x24 && ~x6 && x7 && ~x23 && x9 && x10 && ~x8 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && ~x24 && ~x6 && x7 && ~x23 && x9 && ~x10 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && ~x24 && ~x6 && x7 && ~x23 && x9 && ~x10 && ~x8 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && ~x24 && ~x6 && x7 && ~x23 && ~x9 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && ~x24 && ~x6 && x7 && ~x23 && ~x9 && x8 && ~x10 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && ~x24 && ~x6 && x7 && ~x23 && ~x9 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s98;
						end
					else if( x69 && x70 && ~x62 && ~x63 && ~x64 && ~x24 && ~x6 && ~x7 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && ~x70 && x65 && x60 && x61 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s707;
						end
					else if( x69 && ~x70 && x65 && x60 && ~x61 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x60 && ~x61 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && x60 && ~x61 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( x69 && ~x70 && x65 && x60 && ~x61 && ~x18 )
						nx_state = s118;
					else if( x69 && ~x70 && x65 && ~x60 && x62 && x61 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x70 && x65 && ~x60 && x62 && ~x61 )
						nx_state = s331;
					else if( x69 && ~x70 && x65 && ~x60 && ~x62 && x61 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && ~x60 && ~x62 && x61 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && ~x70 && x65 && ~x60 && ~x62 && x61 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( x69 && ~x70 && x65 && ~x60 && ~x62 && x61 && ~x18 )
						nx_state = s118;
					else if( x69 && ~x70 && x65 && ~x60 && ~x62 && ~x61 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x69 && ~x70 && ~x65 && x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x69 && ~x70 && ~x65 && x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && x21 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x21 && x22 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( x69 && ~x70 && ~x65 && ~x21 && x22 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( x69 && ~x70 && ~x65 && ~x21 && x22 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x21 && x22 && x23 && ~x17 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x21 && x22 && ~x23 && x18 && x14 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && ~x21 && x22 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s47;
					else if( x69 && ~x70 && ~x65 && ~x21 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x21 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x70 && ~x65 && ~x21 && ~x22 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s362;
						end
					else if( ~x69 && x44 && x43 && x3 && x23 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x69 && x44 && x43 && x3 && ~x23 )
						nx_state = s227;
					else if( ~x69 && x44 && x43 && ~x3 )
						nx_state = s1;
					else if( ~x69 && x44 && ~x43 && x2 && x23 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x69 && x44 && ~x43 && x2 && ~x23 )
						nx_state = s227;
					else if( ~x69 && x44 && ~x43 && ~x2 )
						nx_state = s1;
					else if( ~x69 && ~x44 && x10 && x11 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x69 && ~x44 && x10 && x11 && ~x4 )
						nx_state = s227;
					else if( ~x69 && ~x44 && x10 && ~x11 )
						nx_state = s1;
					else if( ~x69 && ~x44 && ~x10 && x13 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x69 && ~x44 && ~x10 && x13 && ~x4 )
						nx_state = s227;
					else if( ~x69 && ~x44 && ~x10 && ~x13 )
						nx_state = s1;
					else nx_state = s227;
				s228 : if( x70 && x62 )
						begin
							y5 = 1'b1;	
							nx_state = s950;
						end
					else if( x70 && ~x62 && x63 && x31 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x70 && ~x62 && x63 && x31 && ~x15 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && x63 && ~x31 && x7 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x70 && ~x62 && x63 && ~x31 && ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x66 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x66 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x66 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && x66 && ~x14 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && x21 && x9 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && x21 && ~x9 && x6 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && x21 && ~x9 && x6 && ~x7 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && x21 && ~x9 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && x21 && ~x9 && ~x6 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x21 && x5 )
						begin
							y30 = 1'b1;	
							nx_state = s416;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x21 && ~x5 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x23 )
						nx_state = s1;
					else if( ~x70 && x65 && x60 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s592;
						end
					else if( ~x70 && x65 && ~x60 )
						begin
							y11 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x70 && ~x65 && x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && ~x65 && x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && ~x65 && x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && x22 && x23 && x10 && x12 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x70 && ~x65 && ~x21 && x22 && x23 && x10 && x12 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x70 && ~x65 && ~x21 && x22 && x23 && x10 && x12 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && x22 && x23 && x10 && x12 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && x22 && x23 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s365;
						end
					else if( ~x70 && ~x65 && ~x21 && x22 && x23 && ~x10 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x70 && ~x65 && ~x21 && x22 && x23 && ~x10 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x70 && ~x65 && ~x21 && x22 && x23 && ~x10 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && x22 && x23 && ~x10 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && x22 && ~x23 && x18 && x14 )
						nx_state = s47;
					else if( ~x70 && ~x65 && ~x21 && x22 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s47;
					else if( ~x70 && ~x65 && ~x21 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && ~x22 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s362;
						end
					else nx_state = s228;
				s229 : if( x21 && x15 && x10 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s274;
						end
					else if( x21 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x21 && x15 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s124;
						end
					else if( x21 && ~x15 && x16 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x21 && ~x15 && ~x16 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s357;
						end
					else if( ~x21 && x22 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( ~x21 && ~x22 )
						nx_state = s1;
					else nx_state = s229;
				s230 : if( x62 && x12 )
						begin
							y16 = 1'b1;	
							nx_state = s293;
						end
					else if( x62 && ~x12 )
						nx_state = s230;
					else if( ~x62 && x15 && x13 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else if( ~x62 && x15 && ~x13 )
						begin
							y16 = 1'b1;	
							nx_state = s293;
						end
					else if( ~x62 && ~x15 && x12 )
						begin
							y16 = 1'b1;	
							nx_state = s293;
						end
					else if( ~x62 && ~x15 && ~x12 )
						nx_state = s230;
					else nx_state = s230;
				s231 : if( x62 && x6 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x62 && ~x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x62 && x15 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	
							nx_state = s276;
						end
					else if( ~x62 && ~x15 && x6 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x62 && ~x15 && ~x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else nx_state = s231;
				s232 : if( 1'b1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s951;
						end
					else nx_state = s232;
				s233 : if( x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x21 && ~x19 )
						nx_state = s1;
					else if( ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x21 && ~x20 )
						nx_state = s1;
					else nx_state = s233;
				s234 : if( x70 && x11 )
						begin
							y2 = 1'b1;	y22 = 1'b1;	
							nx_state = s952;
						end
					else if( x70 && ~x11 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && x65 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x5 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x65 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x65 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x21 && ~x19 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x70 && ~x65 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x70 && ~x65 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && ~x20 )
						nx_state = s1;
					else nx_state = s234;
				s235 : if( x65 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x5 )
						nx_state = s1;
					else if( ~x65 && x21 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x65 && ~x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s224;
						end
					else nx_state = s235;
				s236 : if( x70 && x69 && x64 && x62 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s953;
						end
					else if( x70 && x69 && x64 && x62 && ~x17 )
						begin
							y1 = 1'b1;	y12 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s382;
						end
					else if( x70 && x69 && x64 && ~x62 && x66 && x21 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && x69 && x64 && ~x62 && x66 && x21 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && x69 && x64 && ~x62 && x66 && x21 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && x69 && x64 && ~x62 && x66 && x21 && ~x10 )
						nx_state = s1;
					else if( x70 && x69 && x64 && ~x62 && x66 && ~x21 )
						begin
							y29 = 1'b1;	
							nx_state = s771;
						end
					else if( x70 && x69 && x64 && ~x62 && ~x66 && x67 && x11 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x70 && x69 && x64 && ~x62 && ~x66 && x67 && x11 && ~x4 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s577;
						end
					else if( x70 && x69 && x64 && ~x62 && ~x66 && x67 && ~x11 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && x69 && x64 && ~x62 && ~x66 && ~x67 && x10 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && x69 && x64 && ~x62 && ~x66 && ~x67 && ~x10 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x70 && x69 && x64 && ~x62 && ~x66 && ~x67 && ~x10 && ~x4 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s577;
						end
					else if( x70 && x69 && ~x64 && x62 && x17 && x18 && x5 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x70 && x69 && ~x64 && x62 && x17 && x18 && ~x5 && x6 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x70 && x69 && ~x64 && x62 && x17 && x18 && ~x5 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x70 && x69 && ~x64 && x62 && x17 && ~x18 && x2 )
						nx_state = s1;
					else if( x70 && x69 && ~x64 && x62 && x17 && ~x18 && ~x2 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s215;
						end
					else if( x70 && x69 && ~x64 && x62 && ~x17 && x9 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x70 && x69 && ~x64 && x62 && ~x17 && ~x9 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && x7 && x6 && x12 && x10 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && x7 && x6 && x12 && ~x10 && x11 && x13 )
						begin
							y13 = 1'b1;	
							nx_state = s240;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && x7 && x6 && x12 && ~x10 && x11 && ~x13 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && x7 && x6 && x12 && ~x10 && x11 && ~x13 && x19 && ~x14 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && x7 && x6 && x12 && ~x10 && x11 && ~x13 && ~x19 )
						nx_state = s1;
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && x7 && x6 && x12 && ~x10 && ~x11 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y32 = 1'b1;	
							y53 = 1'b1;	
							nx_state = s954;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && x7 && x6 && ~x12 && x10 )
						begin
							y25 = 1'b1;	
							nx_state = s955;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && x7 && x6 && ~x12 && ~x10 && x11 && x14 )
						begin
							y13 = 1'b1;	
							nx_state = s240;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && x7 && x6 && ~x12 && ~x10 && x11 && ~x14 && x19 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && x7 && x6 && ~x12 && ~x10 && x11 && ~x14 && x19 && ~x13 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && x7 && x6 && ~x12 && ~x10 && x11 && ~x14 && ~x19 )
						nx_state = s1;
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && x7 && x6 && ~x12 && ~x10 && ~x11 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y54 = 1'b1;	
							nx_state = s956;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && x7 && ~x6 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s957;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && x7 && ~x6 && ~x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s958;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && x5 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s957;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && x5 && ~x9 && x10 && x11 && x12 && x6 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && x5 && ~x9 && x10 && x11 && x12 && ~x6 )
						begin
							y4 = 1'b1;	y33 = 1'b1;	y34 = 1'b1;	
							y38 = 1'b1;	y42 = 1'b1;	
							nx_state = s720;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && x5 && ~x9 && x10 && x11 && ~x12 && x6 )
						begin
							y29 = 1'b1;	
							nx_state = s771;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && x5 && ~x9 && x10 && x11 && ~x12 && ~x6 )
						begin
							y4 = 1'b1;	y33 = 1'b1;	y34 = 1'b1;	
							y38 = 1'b1;	y41 = 1'b1;	
							nx_state = s720;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && x5 && ~x9 && x10 && ~x11 && x6 && x12 )
						begin
							y30 = 1'b1;	
							nx_state = s291;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && x5 && ~x9 && x10 && ~x11 && x6 && ~x12 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && x5 && ~x9 && x10 && ~x11 && ~x6 )
						begin
							y4 = 1'b1;	y33 = 1'b1;	y34 = 1'b1;	
							y38 = 1'b1;	y40 = 1'b1;	
							nx_state = s720;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && x5 && ~x9 && ~x10 && x11 && x12 && x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s959;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && x5 && ~x9 && ~x10 && x11 && x12 && ~x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y59 = 1'b1;	
							y60 = 1'b1;	
							nx_state = s960;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && x5 && ~x9 && ~x10 && x11 && ~x12 && x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y31 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s720;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && x5 && ~x9 && ~x10 && x11 && ~x12 && ~x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y63 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s961;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && x5 && ~x9 && ~x10 && ~x11 && x12 && x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && x5 && ~x9 && ~x10 && ~x11 && x12 && ~x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y61 = 1'b1;	
							y62 = 1'b1;	
							nx_state = s962;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && x5 && ~x9 && ~x10 && ~x11 && ~x12 && x6 )
						begin
							y36 = 1'b1;	
							nx_state = s963;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && x5 && ~x9 && ~x10 && ~x11 && ~x12 && ~x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y65 = 1'b1;	
							y66 = 1'b1;	
							nx_state = s646;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && ~x5 && x8 && x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && ~x5 && x8 && ~x6 && x11 && x12 )
						begin
							y4 = 1'b1;	y34 = 1'b1;	y38 = 1'b1;	
							y39 = 1'b1;	y42 = 1'b1;	
							nx_state = s720;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && ~x5 && x8 && ~x6 && x11 && ~x12 )
						begin
							y4 = 1'b1;	y34 = 1'b1;	y38 = 1'b1;	
							y39 = 1'b1;	y41 = 1'b1;	
							nx_state = s720;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && ~x5 && x8 && ~x6 && ~x11 )
						begin
							y4 = 1'b1;	y34 = 1'b1;	y38 = 1'b1;	
							y39 = 1'b1;	y40 = 1'b1;	
							nx_state = s720;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && x4 && ~x7 && ~x5 && ~x8 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s958;
						end
					else if( x70 && x69 && ~x64 && ~x62 && x3 && ~x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s964;
						end
					else if( x70 && x69 && ~x64 && ~x62 && ~x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x70 && ~x69 && x62 && x61 && x9 )
						begin
							y13 = 1'b1;	
							nx_state = s240;
						end
					else if( x70 && ~x69 && x62 && x61 && ~x9 && x3 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( x70 && ~x69 && x62 && x61 && ~x9 && ~x3 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( x70 && ~x69 && x62 && ~x61 && x29 && x50 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s842;
						end
					else if( x70 && ~x69 && x62 && ~x61 && x29 && ~x50 )
						nx_state = s236;
					else if( x70 && ~x69 && x62 && ~x61 && ~x29 && x60 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( x70 && ~x69 && x62 && ~x61 && ~x29 && ~x60 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( x70 && ~x69 && ~x62 && x33 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s801;
						end
					else if( x70 && ~x69 && ~x62 && ~x33 )
						nx_state = s236;
					else if( ~x70 && x69 && x21 )
						nx_state = s1;
					else if( ~x70 && x69 && ~x21 && x22 && x12 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s377;
						end
					else if( ~x70 && x69 && ~x21 && x22 && ~x12 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x70 && x69 && ~x21 && x22 && ~x12 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x70 && x69 && ~x21 && x22 && ~x12 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x70 && x69 && ~x21 && x22 && ~x12 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x69 && ~x21 && ~x22 && x7 && x18 && x15 )
						begin
							y8 = 1'b1;	y18 = 1'b1;	
							nx_state = s152;
						end
					else if( ~x70 && x69 && ~x21 && ~x22 && x7 && x18 && ~x15 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s6;
						end
					else if( ~x70 && x69 && ~x21 && ~x22 && x7 && ~x18 && x19 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s835;
						end
					else if( ~x70 && x69 && ~x21 && ~x22 && x7 && ~x18 && x19 && ~x15 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x69 && ~x21 && ~x22 && x7 && ~x18 && ~x19 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x70 && x69 && ~x21 && ~x22 && ~x7 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s376;
						end
					else if( ~x70 && ~x69 && x44 && x11 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && ~x69 && x44 && ~x11 && x9 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && ~x69 && x44 && ~x11 && ~x9 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x70 && ~x69 && ~x44 && x46 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && ~x69 && ~x44 && ~x46 && x45 && x47 && x10 && x9 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && ~x69 && ~x44 && ~x46 && x45 && x47 && x10 && ~x9 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x70 && ~x69 && ~x44 && ~x46 && x45 && x47 && ~x10 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x70 && ~x69 && ~x44 && ~x46 && x45 && ~x47 && x12 && x4 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && ~x69 && ~x44 && ~x46 && x45 && ~x47 && x12 && ~x4 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s578;
						end
					else if( ~x70 && ~x69 && ~x44 && ~x46 && x45 && ~x47 && ~x12 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && ~x69 && ~x44 && ~x46 && ~x45 && x10 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && ~x69 && ~x44 && ~x46 && ~x45 && ~x10 && x4 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && ~x69 && ~x44 && ~x46 && ~x45 && ~x10 && ~x4 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s578;
						end
					else nx_state = s236;
				s237 : if( x70 && x5 )
						begin
							y1 = 1'b1;	y46 = 1'b1;	
							nx_state = s966;
						end
					else if( x70 && ~x5 && x32 && x13 && x15 && x33 )
						begin
							y9 = 1'b1;	
							nx_state = s967;
						end
					else if( x70 && ~x5 && x32 && x13 && x15 && ~x33 && x14 )
						begin
							y6 = 1'b1;	y35 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s338;
						end
					else if( x70 && ~x5 && x32 && x13 && x15 && ~x33 && ~x14 && x16 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s347;
						end
					else if( x70 && ~x5 && x32 && x13 && x15 && ~x33 && ~x14 && ~x16 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s348;
						end
					else if( x70 && ~x5 && x32 && x13 && ~x15 && x33 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s968;
						end
					else if( x70 && ~x5 && x32 && x13 && ~x15 && ~x33 && x14 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s349;
						end
					else if( x70 && ~x5 && x32 && x13 && ~x15 && ~x33 && ~x14 && x7 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y35 = 1'b1;	y40 = 1'b1;	
							nx_state = s351;
						end
					else if( x70 && ~x5 && x32 && x13 && ~x15 && ~x33 && ~x14 && ~x7 )
						begin
							y8 = 1'b1;	y36 = 1'b1;	y42 = 1'b1;	
							nx_state = s969;
						end
					else if( x70 && ~x5 && x32 && ~x13 && x14 && x33 && x15 && x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s970;
						end
					else if( x70 && ~x5 && x32 && ~x13 && x14 && x33 && x15 && ~x12 && x10 && x11 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s470;
						end
					else if( x70 && ~x5 && x32 && ~x13 && x14 && x33 && x15 && ~x12 && x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x5 && x32 && ~x13 && x14 && x33 && x15 && ~x12 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x5 && x32 && ~x13 && x14 && x33 && ~x15 && x11 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s971;
						end
					else if( x70 && ~x5 && x32 && ~x13 && x14 && x33 && ~x15 && ~x11 && x10 && x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s470;
						end
					else if( x70 && ~x5 && x32 && ~x13 && x14 && x33 && ~x15 && ~x11 && x10 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x5 && x32 && ~x13 && x14 && x33 && ~x15 && ~x11 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x5 && x32 && ~x13 && x14 && ~x33 && x15 && x7 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s972;
						end
					else if( x70 && ~x5 && x32 && ~x13 && x14 && ~x33 && x15 && ~x7 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s973;
						end
					else if( x70 && ~x5 && x32 && ~x13 && x14 && ~x33 && ~x15 && x7 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s340;
						end
					else if( x70 && ~x5 && x32 && ~x13 && x14 && ~x33 && ~x15 && ~x7 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s974;
						end
					else if( x70 && ~x5 && x32 && ~x13 && ~x14 && x15 && x33 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x70 && ~x5 && x32 && ~x13 && ~x14 && x15 && ~x33 && x17 )
						nx_state = s1;
					else if( x70 && ~x5 && x32 && ~x13 && ~x14 && x15 && ~x33 && ~x17 && x7 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s975;
						end
					else if( x70 && ~x5 && x32 && ~x13 && ~x14 && x15 && ~x33 && ~x17 && ~x7 )
						begin
							y30 = 1'b1;	
							nx_state = s976;
						end
					else if( x70 && ~x5 && x32 && ~x13 && ~x14 && ~x15 && x33 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s311;
						end
					else if( x70 && ~x5 && x32 && ~x13 && ~x14 && ~x15 && ~x33 && x18 )
						nx_state = s1;
					else if( x70 && ~x5 && x32 && ~x13 && ~x14 && ~x15 && ~x33 && ~x18 && x7 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s977;
						end
					else if( x70 && ~x5 && x32 && ~x13 && ~x14 && ~x15 && ~x33 && ~x18 && ~x7 )
						begin
							y6 = 1'b1;	y47 = 1'b1;	
							nx_state = s978;
						end
					else if( x70 && ~x5 && ~x32 && x13 && x14 && x33 && x15 && x7 )
						begin
							y6 = 1'b1;	y35 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s338;
						end
					else if( x70 && ~x5 && ~x32 && x13 && x14 && x33 && x15 && ~x7 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y27 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s339;
						end
					else if( x70 && ~x5 && ~x32 && x13 && x14 && x33 && ~x15 )
						begin
							y53 = 1'b1;	
							nx_state = s344;
						end
					else if( x70 && ~x5 && ~x32 && x13 && x14 && ~x33 && x7 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y27 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s339;
						end
					else if( x70 && ~x5 && ~x32 && x13 && x14 && ~x33 && ~x7 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s350;
						end
					else if( x70 && ~x5 && ~x32 && x13 && ~x14 && x15 && x33 && x31 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( x70 && ~x5 && ~x32 && x13 && ~x14 && x15 && x33 && ~x31 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x70 && ~x5 && ~x32 && x13 && ~x14 && x15 && x33 && ~x31 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x70 && ~x5 && ~x32 && x13 && ~x14 && x15 && x33 && ~x31 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x5 && ~x32 && x13 && ~x14 && x15 && x33 && ~x31 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x5 && ~x32 && x13 && ~x14 && x15 && ~x33 && x7 )
						begin
							y8 = 1'b1;	y36 = 1'b1;	y42 = 1'b1;	
							nx_state = s969;
						end
					else if( x70 && ~x5 && ~x32 && x13 && ~x14 && x15 && ~x33 && ~x7 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s343;
						end
					else if( x70 && ~x5 && ~x32 && x13 && ~x14 && ~x15 && x33 && x16 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( x70 && ~x5 && ~x32 && x13 && ~x14 && ~x15 && x33 && ~x16 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x70 && ~x5 && ~x32 && x13 && ~x14 && ~x15 && x33 && ~x16 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x70 && ~x5 && ~x32 && x13 && ~x14 && ~x15 && x33 && ~x16 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x5 && ~x32 && x13 && ~x14 && ~x15 && x33 && ~x16 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x5 && ~x32 && x13 && ~x14 && ~x15 && ~x33 && x7 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s979;
						end
					else if( x70 && ~x5 && ~x32 && x13 && ~x14 && ~x15 && ~x33 && ~x7 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s980;
						end
					else if( x70 && ~x5 && ~x32 && ~x13 && x33 && x14 && x15 && x8 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( x70 && ~x5 && ~x32 && ~x13 && x33 && x14 && x15 && ~x8 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x70 && ~x5 && ~x32 && ~x13 && x33 && x14 && x15 && ~x8 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x70 && ~x5 && ~x32 && ~x13 && x33 && x14 && x15 && ~x8 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x5 && ~x32 && ~x13 && x33 && x14 && x15 && ~x8 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x5 && ~x32 && ~x13 && x33 && x14 && ~x15 && x30 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( x70 && ~x5 && ~x32 && ~x13 && x33 && x14 && ~x15 && ~x30 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x70 && ~x5 && ~x32 && ~x13 && x33 && x14 && ~x15 && ~x30 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x70 && ~x5 && ~x32 && ~x13 && x33 && x14 && ~x15 && ~x30 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x5 && ~x32 && ~x13 && x33 && x14 && ~x15 && ~x30 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x5 && ~x32 && ~x13 && x33 && ~x14 && x15 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( x70 && ~x5 && ~x32 && ~x13 && x33 && ~x14 && ~x15 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s345;
						end
					else if( x70 && ~x5 && ~x32 && ~x13 && ~x33 && x7 )
						begin
							y6 = 1'b1;	y35 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s338;
						end
					else if( x70 && ~x5 && ~x32 && ~x13 && ~x33 && ~x7 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s347;
						end
					else if( ~x70 && x21 && x19 && x20 && x17 && x5 )
						begin
							y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s572;
						end
					else if( ~x70 && x21 && x19 && x20 && x17 && ~x5 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && x21 && x19 && x20 && x17 && ~x5 && x3 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x21 && x19 && x20 && x17 && ~x5 && ~x3 )
						nx_state = s1;
					else if( ~x70 && x21 && x19 && x20 && ~x17 && x4 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s377;
						end
					else if( ~x70 && x21 && x19 && x20 && ~x17 && ~x4 && x3 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && x21 && x19 && x20 && ~x17 && ~x4 && x3 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x21 && x19 && x20 && ~x17 && ~x4 && ~x3 )
						nx_state = s1;
					else if( ~x70 && x21 && x19 && ~x20 && x12 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x70 && x21 && x19 && ~x20 && x12 && ~x2 && x17 && x8 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x70 && x21 && x19 && ~x20 && x12 && ~x2 && x17 && ~x8 )
						begin
							y18 = 1'b1;	
							nx_state = s574;
						end
					else if( ~x70 && x21 && x19 && ~x20 && x12 && ~x2 && ~x17 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( ~x70 && x21 && x19 && ~x20 && x12 && ~x2 && ~x17 && ~x8 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( ~x70 && x21 && x19 && ~x20 && ~x12 && x16 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && x21 && x19 && ~x20 && ~x12 && ~x16 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x70 && x21 && x19 && ~x20 && ~x12 && ~x16 && ~x2 && x8 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x70 && x21 && x19 && ~x20 && ~x12 && ~x16 && ~x2 && ~x8 && x17 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( ~x70 && x21 && x19 && ~x20 && ~x12 && ~x16 && ~x2 && ~x8 && ~x17 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s6;
						end
					else if( ~x70 && x21 && ~x19 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s384;
						end
					else if( ~x70 && x21 && ~x19 && ~x2 && x20 && x12 && x8 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x70 && x21 && ~x19 && ~x2 && x20 && x12 && ~x8 )
						begin
							y18 = 1'b1;	
							nx_state = s574;
						end
					else if( ~x70 && x21 && ~x19 && ~x2 && x20 && ~x12 && x17 && x16 && x8 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x70 && x21 && ~x19 && ~x2 && x20 && ~x12 && x17 && x16 && ~x8 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s377;
						end
					else if( ~x70 && x21 && ~x19 && ~x2 && x20 && ~x12 && x17 && ~x16 && x14 && x8 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x70 && x21 && ~x19 && ~x2 && x20 && ~x12 && x17 && ~x16 && x14 && ~x8 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s377;
						end
					else if( ~x70 && x21 && ~x19 && ~x2 && x20 && ~x12 && x17 && ~x16 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x19 && ~x2 && x20 && ~x12 && ~x17 && x16 && x15 && x8 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x70 && x21 && ~x19 && ~x2 && x20 && ~x12 && ~x17 && x16 && x15 && ~x8 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s377;
						end
					else if( ~x70 && x21 && ~x19 && ~x2 && x20 && ~x12 && ~x17 && x16 && ~x15 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x19 && ~x2 && x20 && ~x12 && ~x17 && ~x16 && x13 && x8 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x70 && x21 && ~x19 && ~x2 && x20 && ~x12 && ~x17 && ~x16 && x13 && ~x8 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s377;
						end
					else if( ~x70 && x21 && ~x19 && ~x2 && x20 && ~x12 && ~x17 && ~x16 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x19 && ~x2 && ~x20 && x8 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x70 && x21 && ~x19 && ~x2 && ~x20 && ~x8 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s981;
						end
					else if( ~x70 && x21 && ~x19 && ~x2 && ~x20 && ~x8 && ~x12 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( ~x70 && ~x21 && x22 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else nx_state = s237;
				s238 : if( x63 && x1 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x63 && x1 && ~x2 && x5 && x3 )
						nx_state = s238;
					else if( x63 && x1 && ~x2 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x63 && x1 && ~x2 && ~x5 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	
							nx_state = s7;
						end
					else if( x63 && ~x1 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( ~x63 && x64 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x64 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x64 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x63 && x64 && ~x9 )
						nx_state = s1;
					else if( ~x63 && ~x64 && x31 && x14 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && ~x64 && x31 && ~x14 )
						begin
							y47 = 1'b1;	y53 = 1'b1;	y61 = 1'b1;	
							y69 = 1'b1;	
							nx_state = s982;
						end
					else if( ~x63 && ~x64 && ~x31 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s568;
						end
					else if( ~x63 && ~x64 && ~x31 && ~x14 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else nx_state = s238;
				s239 : if( x63 && x11 )
						begin
							y18 = 1'b1;	y27 = 1'b1;	
							nx_state = s983;
						end
					else if( x63 && ~x11 )
						begin
							y10 = 1'b1;	y20 = 1'b1;	y26 = 1'b1;	
							nx_state = s984;
						end
					else if( ~x63 && x64 )
						begin
							y7 = 1'b1;	
							nx_state = s985;
						end
					else if( ~x63 && ~x64 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s986;
						end
					else nx_state = s239;
				s240 : if( x69 && x62 && x64 && x17 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							nx_state = s987;
						end
					else if( x69 && x62 && x64 && ~x17 )
						begin
							y1 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s988;
						end
					else if( x69 && x62 && ~x64 && x25 && x9 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && x62 && ~x64 && x25 && ~x9 )
						begin
							y13 = 1'b1;	
							nx_state = s240;
						end
					else if( x69 && x62 && ~x64 && ~x25 && x13 )
						begin
							y13 = 1'b1;	
							nx_state = s240;
						end
					else if( x69 && x62 && ~x64 && ~x25 && ~x13 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x69 && ~x62 )
						begin
							y13 = 1'b1;	
							nx_state = s769;
						end
					else if( ~x69 && x61 && x33 )
						begin
							y10 = 1'b1;	
							nx_state = s841;
						end
					else if( ~x69 && x61 && ~x33 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( ~x69 && x61 && ~x33 && ~x13 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s840;
						end
					else if( ~x69 && ~x61 && x50 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s842;
						end
					else if( ~x69 && ~x61 && ~x50 )
						nx_state = s240;
					else nx_state = s240;
				s241 : if( x70 && x62 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y37 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s989;
						end
					else if( x70 && ~x62 && x65 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x70 && ~x62 && ~x65 && x67 )
						begin
							y5 = 1'b1;	y13 = 1'b1;	y17 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s990;
						end
					else if( x70 && ~x62 && ~x65 && ~x67 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x65 && x22 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	
							nx_state = s486;
						end
					else if( ~x70 && x65 && ~x22 && x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x65 && ~x22 && ~x23 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x65 && x68 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x65 && x68 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x65 && x68 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x68 && ~x9 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x68 && x23 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x70 && ~x65 && ~x68 && ~x23 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else nx_state = s241;
				s242 : if( x65 && x60 && x61 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x65 && x60 && x61 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x65 && x60 && x61 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x65 && x60 && x61 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x65 && x60 && ~x61 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x65 && x60 && ~x61 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x65 && x60 && ~x61 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( x65 && x60 && ~x61 && ~x18 )
						nx_state = s118;
					else if( x65 && ~x60 && x61 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x65 && ~x60 && x61 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x65 && ~x60 && x61 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x65 && ~x60 && x61 && x62 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x60 && x61 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x65 && ~x60 && x61 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x65 && ~x60 && x61 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( x65 && ~x60 && x61 && ~x62 && ~x18 )
						nx_state = s118;
					else if( x65 && ~x60 && ~x61 )
						nx_state = s47;
					else if( ~x65 && x20 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x65 && ~x20 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x65 && ~x20 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x65 && ~x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x20 && ~x18 )
						nx_state = s1;
					else nx_state = s242;
				s243 : if( x70 && x63 && x20 )
						begin
							y28 = 1'b1;	
							nx_state = s991;
						end
					else if( x70 && x63 && ~x20 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( x70 && ~x63 )
						begin
							y6 = 1'b1;	
							nx_state = s368;
						end
					else if( ~x70 && x65 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x65 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s122;
						end
					else nx_state = s243;
				s244 : if( x65 && x60 )
						nx_state = s143;
					else if( x65 && ~x60 && x61 )
						nx_state = s143;
					else if( x65 && ~x60 && ~x61 )
						nx_state = s47;
					else if( ~x65 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else nx_state = s244;
				s245 : if( x65 && x66 )
						nx_state = s47;
					else if( x65 && ~x66 && x21 && x5 )
						begin
							y3 = 1'b1;	y12 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s113;
						end
					else if( x65 && ~x66 && x21 && ~x5 && x6 && x18 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x65 && ~x66 && x21 && ~x5 && x6 && x18 && x15 && ~x17 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	
							nx_state = s807;
						end
					else if( x65 && ~x66 && x21 && ~x5 && x6 && x18 && ~x15 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x65 && ~x66 && x21 && ~x5 && x6 && ~x18 && x19 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x65 && ~x66 && x21 && ~x5 && x6 && ~x18 && x19 && x15 && ~x17 )
						begin
							y8 = 1'b1;	
							nx_state = s568;
						end
					else if( x65 && ~x66 && x21 && ~x5 && x6 && ~x18 && x19 && ~x15 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s795;
						end
					else if( x65 && ~x66 && x21 && ~x5 && x6 && ~x18 && ~x19 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s110;
						end
					else if( x65 && ~x66 && x21 && ~x5 && ~x6 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s666;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x23 && x7 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x23 && x7 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x23 && x7 && ~x18 && x19 && x15 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s666;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x23 && x7 && ~x18 && x19 && ~x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x23 && x7 && ~x18 && ~x19 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s112;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x23 && ~x7 )
						begin
							y3 = 1'b1;	y12 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s113;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x23 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s301;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && x23 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s301;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x23 && x7 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x23 && x7 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x23 && x7 && ~x18 && x19 && x15 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s666;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x23 && x7 && ~x18 && x19 && ~x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x23 && x7 && ~x18 && ~x19 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s112;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x23 && ~x7 )
						begin
							y3 = 1'b1;	y12 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s113;
						end
					else if( ~x65 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else nx_state = s245;
				s246 : if( x70 && x62 && x66 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s992;
						end
					else if( x70 && x62 && ~x66 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x70 && x62 && ~x66 && ~x11 && x10 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( x70 && x62 && ~x66 && ~x11 && ~x10 )
						nx_state = s246;
					else if( x70 && ~x62 && x63 && x66 && x31 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x70 && ~x62 && x63 && x66 && x31 && ~x15 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && x63 && x66 && ~x31 && x7 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x70 && ~x62 && x63 && x66 && ~x31 && ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && x63 && ~x66 && x15 )
						nx_state = s1;
					else if( x70 && ~x62 && x63 && ~x66 && ~x15 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x70 && ~x62 && x63 && ~x66 && ~x15 && ~x11 && x10 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( x70 && ~x62 && x63 && ~x66 && ~x15 && ~x11 && ~x10 )
						nx_state = s246;
					else if( x70 && ~x62 && ~x63 && x64 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x23 )
						nx_state = s1;
					else if( ~x70 && x65 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x70 && ~x65 && x66 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x70 && ~x65 && x66 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x70 && ~x65 && x66 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && ~x4 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && x20 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s668;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else nx_state = s246;
				s247 : if( x69 && x65 && x60 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s135;
						end
					else if( x69 && x65 && ~x60 && x61 && x62 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y23 = 1'b1;	
							nx_state = s993;
						end
					else if( x69 && x65 && ~x60 && x61 && ~x62 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s135;
						end
					else if( x69 && x65 && ~x60 && ~x61 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x69 && ~x65 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x69 && x26 && x28 && x9 && x63 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( ~x69 && x26 && x28 && x9 && ~x63 && x64 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( ~x69 && x26 && x28 && x9 && ~x63 && ~x64 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s917;
						end
					else if( ~x69 && x26 && x28 && ~x9 && x23 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( ~x69 && x26 && x28 && ~x9 && ~x23 && x63 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x69 && x26 && x28 && ~x9 && ~x23 && ~x63 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && x26 && ~x28 && x63 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( ~x69 && x26 && ~x28 && ~x63 && x64 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( ~x69 && x26 && ~x28 && ~x63 && ~x64 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s944;
						end
					else if( ~x69 && ~x26 && x63 && x27 && x1 && x33 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( ~x69 && ~x26 && x63 && x27 && x1 && ~x33 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( ~x69 && ~x26 && x63 && x27 && x1 && ~x33 && ~x34 )
						nx_state = s247;
					else if( ~x69 && ~x26 && x63 && x27 && ~x1 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( ~x69 && ~x26 && x63 && ~x27 && x1 && x5 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s922;
						end
					else if( ~x69 && ~x26 && x63 && ~x27 && x1 && x5 && ~x3 && x4 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s994;
						end
					else if( ~x69 && ~x26 && x63 && ~x27 && x1 && x5 && ~x3 && ~x4 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s995;
						end
					else if( ~x69 && ~x26 && x63 && ~x27 && x1 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x69 && ~x26 && x63 && ~x27 && ~x1 && x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( ~x69 && ~x26 && x63 && ~x27 && ~x1 && ~x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( ~x69 && ~x26 && ~x63 && x27 && x64 && x1 && x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( ~x69 && ~x26 && ~x63 && x27 && x64 && x1 && ~x2 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( ~x69 && ~x26 && ~x63 && x27 && x64 && x1 && ~x2 && ~x3 )
						nx_state = s247;
					else if( ~x69 && ~x26 && ~x63 && x27 && x64 && ~x1 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( ~x69 && ~x26 && ~x63 && x27 && ~x64 && x36 && x32 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s944;
						end
					else if( ~x69 && ~x26 && ~x63 && x27 && ~x64 && x36 && ~x32 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( ~x69 && ~x26 && ~x63 && x27 && ~x64 && x36 && ~x32 && ~x3 )
						nx_state = s247;
					else if( ~x69 && ~x26 && ~x63 && x27 && ~x64 && ~x36 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s917;
						end
					else if( ~x69 && ~x26 && ~x63 && ~x27 && x64 && x1 && x5 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s922;
						end
					else if( ~x69 && ~x26 && ~x63 && ~x27 && x64 && x1 && x5 && ~x3 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( ~x69 && ~x26 && ~x63 && ~x27 && x64 && x1 && x5 && ~x3 && ~x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else if( ~x69 && ~x26 && ~x63 && ~x27 && x64 && x1 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && ~x26 && ~x63 && ~x27 && x64 && ~x1 && x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( ~x69 && ~x26 && ~x63 && ~x27 && x64 && ~x1 && ~x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( ~x69 && ~x26 && ~x63 && ~x27 && ~x64 && x36 && x5 && x3 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s923;
						end
					else if( ~x69 && ~x26 && ~x63 && ~x27 && ~x64 && x36 && x5 && ~x3 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s924;
						end
					else if( ~x69 && ~x26 && ~x63 && ~x27 && ~x64 && x36 && x5 && ~x3 && ~x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else if( ~x69 && ~x26 && ~x63 && ~x27 && ~x64 && x36 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && ~x26 && ~x63 && ~x27 && ~x64 && ~x36 && x2 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s944;
						end
					else if( ~x69 && ~x26 && ~x63 && ~x27 && ~x64 && ~x36 && ~x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else nx_state = s247;
				s248 : if( x69 && x65 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x69 && ~x65 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x69 && x63 && x46 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s996;
						end
					else if( ~x69 && x63 && ~x46 && x34 && x2 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s691;
						end
					else if( ~x69 && x63 && ~x46 && x34 && ~x2 )
						nx_state = s248;
					else if( ~x69 && x63 && ~x46 && ~x34 && x35 && x2 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s997;
						end
					else if( ~x69 && x63 && ~x46 && ~x34 && x35 && ~x2 )
						nx_state = s248;
					else if( ~x69 && x63 && ~x46 && ~x34 && ~x35 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s998;
						end
					else if( ~x69 && x63 && ~x46 && ~x34 && ~x35 && ~x2 )
						nx_state = s248;
					else if( ~x69 && ~x63 && x15 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s477;
						end
					else if( ~x69 && ~x63 && ~x15 && x3 && x64 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( ~x69 && ~x63 && ~x15 && x3 && x64 && ~x2 )
						nx_state = s248;
					else if( ~x69 && ~x63 && ~x15 && x3 && ~x64 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s700;
						end
					else if( ~x69 && ~x63 && ~x15 && x3 && ~x64 && ~x2 )
						nx_state = s248;
					else if( ~x69 && ~x63 && ~x15 && ~x3 && x4 && x64 && x2 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s997;
						end
					else if( ~x69 && ~x63 && ~x15 && ~x3 && x4 && x64 && ~x2 )
						nx_state = s248;
					else if( ~x69 && ~x63 && ~x15 && ~x3 && x4 && ~x64 && x2 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s999;
						end
					else if( ~x69 && ~x63 && ~x15 && ~x3 && x4 && ~x64 && ~x2 )
						nx_state = s248;
					else if( ~x69 && ~x63 && ~x15 && ~x3 && ~x4 && x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1000;
						end
					else if( ~x69 && ~x63 && ~x15 && ~x3 && ~x4 && ~x2 )
						nx_state = s248;
					else nx_state = s248;
				s249 : if( x65 && x61 && x60 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s384;
						end
					else if( x65 && x61 && ~x60 && x62 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( x65 && x61 && ~x60 && ~x62 && ~x2 && x19 && x15 )
						nx_state = s143;
					else if( x65 && x61 && ~x60 && ~x62 && ~x2 && x19 && ~x15 && x16 )
						begin
							y12 = 1'b1;	
							nx_state = s244;
						end
					else if( x65 && x61 && ~x60 && ~x62 && ~x2 && x19 && ~x15 && ~x16 )
						nx_state = s143;
					else if( x65 && x61 && ~x60 && ~x62 && ~x2 && ~x19 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y24 = 1'b1;	
							nx_state = s136;
						end
					else if( x65 && ~x61 && x60 && x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( x65 && ~x61 && x60 && ~x2 && x19 && x15 )
						nx_state = s143;
					else if( x65 && ~x61 && x60 && ~x2 && x19 && ~x15 && x16 )
						begin
							y12 = 1'b1;	
							nx_state = s244;
						end
					else if( x65 && ~x61 && x60 && ~x2 && x19 && ~x15 && ~x16 )
						nx_state = s143;
					else if( x65 && ~x61 && x60 && ~x2 && ~x19 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y24 = 1'b1;	
							nx_state = s136;
						end
					else if( x65 && ~x61 && ~x60 && x62 )
						nx_state = s47;
					else if( x65 && ~x61 && ~x60 && ~x62 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && x15 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && x15 && ~x7 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && x15 && ~x7 && ~x11 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s242;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && x4 )
						nx_state = s47;
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && ~x4 && x11 && x9 )
						nx_state = s47;
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && ~x4 && x11 && ~x9 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && ~x4 && x11 && ~x9 && ~x7 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s559;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && ~x4 && ~x11 && x9 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && ~x4 && ~x11 && x9 && ~x7 && x10 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && ~x4 && ~x11 && x9 && ~x7 && ~x10 )
						nx_state = s47;
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && x7 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && x7 && ~x8 )
						nx_state = s47;
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && ~x7 && x12 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && ~x7 && ~x12 )
						nx_state = s47;
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && ~x18 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y24 = 1'b1;	
							nx_state = s136;
						end
					else if( ~x65 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s6;
						end
					else nx_state = s249;
				s250 : if( x69 && x65 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x69 && ~x65 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x69 && x63 && x55 && x11 && x25 && x34 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x69 && x63 && x55 && x11 && x25 && ~x34 && x36 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && x63 && x55 && x11 && x25 && ~x34 && ~x36 )
						nx_state = s250;
					else if( ~x69 && x63 && x55 && x11 && ~x25 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( ~x69 && x63 && x55 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x69 && x63 && ~x55 && x53 && x47 )
						nx_state = s250;
					else if( ~x69 && x63 && ~x55 && x53 && ~x47 && x59 && x51 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x69 && x63 && ~x55 && x53 && ~x47 && x59 && ~x51 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && x63 && ~x55 && x53 && ~x47 && ~x59 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && x63 && ~x55 && x53 && ~x47 && ~x59 && ~x34 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x69 && x63 && ~x55 && ~x53 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x69 && ~x63 && x64 && x40 && x11 && x25 && x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && ~x63 && x64 && x40 && x11 && x25 && ~x3 && x5 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && ~x63 && x64 && x40 && x11 && x25 && ~x3 && ~x5 )
						nx_state = s250;
					else if( ~x69 && ~x63 && x64 && x40 && x11 && ~x25 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( ~x69 && ~x63 && x64 && x40 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && ~x63 && x64 && ~x40 && x48 && x42 && x51 && x47 )
						nx_state = s250;
					else if( ~x69 && ~x63 && x64 && ~x40 && x48 && x42 && x51 && ~x47 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && ~x63 && x64 && ~x40 && x48 && x42 && ~x51 && x47 )
						nx_state = s250;
					else if( ~x69 && ~x63 && x64 && ~x40 && x48 && x42 && ~x51 && ~x47 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && ~x63 && x64 && ~x40 && x48 && ~x42 && x47 )
						nx_state = s250;
					else if( ~x69 && ~x63 && x64 && ~x40 && x48 && ~x42 && ~x47 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && ~x63 && x64 && ~x40 && x48 && ~x42 && ~x47 && ~x34 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && ~x63 && x64 && ~x40 && ~x48 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && ~x63 && ~x64 && x44 && x11 && x25 && x42 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s867;
						end
					else if( ~x69 && ~x63 && ~x64 && x44 && x11 && x25 && ~x42 && x5 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && ~x63 && ~x64 && x44 && x11 && x25 && ~x42 && ~x5 )
						nx_state = s250;
					else if( ~x69 && ~x63 && ~x64 && x44 && x11 && ~x25 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s870;
						end
					else if( ~x69 && ~x63 && ~x64 && x44 && ~x11 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s867;
						end
					else if( ~x69 && ~x63 && ~x64 && ~x44 && x53 && x47 )
						nx_state = s250;
					else if( ~x69 && ~x63 && ~x64 && ~x44 && x53 && ~x47 && x48 && x51 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s867;
						end
					else if( ~x69 && ~x63 && ~x64 && ~x44 && x53 && ~x47 && x48 && ~x51 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && ~x63 && ~x64 && ~x44 && x53 && ~x47 && ~x48 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && ~x63 && ~x64 && ~x44 && x53 && ~x47 && ~x48 && ~x34 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s867;
						end
					else if( ~x69 && ~x63 && ~x64 && ~x44 && ~x53 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s867;
						end
					else nx_state = s250;
				s251 : if( x70 && x23 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							y18 = 1'b1;	y29 = 1'b1;	
							nx_state = s1001;
						end
					else if( x70 && x23 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1002;
						end
					else if( x70 && ~x23 && x22 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							y18 = 1'b1;	y29 = 1'b1;	
							nx_state = s1001;
						end
					else if( x70 && ~x23 && x22 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1002;
						end
					else if( x70 && ~x23 && ~x22 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1002;
						end
					else if( x70 && ~x23 && ~x22 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							y18 = 1'b1;	y29 = 1'b1;	
							nx_state = s1001;
						end
					else if( ~x70 && x60 && x61 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x60 && x61 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x60 && x61 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( ~x70 && x60 && x61 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( ~x70 && x60 && ~x61 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x60 && ~x61 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x60 && ~x61 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( ~x70 && x60 && ~x61 && ~x18 )
						nx_state = s118;
					else if( ~x70 && ~x60 && x61 && x62 )
						nx_state = s1;
					else if( ~x70 && ~x60 && x61 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x60 && x61 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x60 && x61 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( ~x70 && ~x60 && x61 && ~x62 && ~x18 )
						nx_state = s118;
					else if( ~x70 && ~x60 && ~x61 )
						nx_state = s47;
					else nx_state = s251;
				s252 : if( x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x4 )
						nx_state = s1;
					else nx_state = s252;
				s253 : if( x70 )
						nx_state = s1;
					else if( ~x70 && x65 && x22 && x21 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && x22 && x21 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && x22 && x21 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && x22 && x21 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && x22 && ~x21 && x18 && x19 )
						nx_state = s1;
					else if( ~x70 && x65 && x22 && ~x21 && x18 && ~x19 && x10 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x70 && x65 && x22 && ~x21 && x18 && ~x19 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && x22 && ~x21 && x18 && ~x19 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && x22 && ~x21 && x18 && ~x19 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && x22 && ~x21 && x18 && ~x19 && ~x10 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && x22 && ~x21 && ~x18 && x19 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && x22 && ~x21 && ~x18 && x19 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && x22 && ~x21 && ~x18 && x19 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && x22 && ~x21 && ~x18 && ~x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && x22 && ~x21 && ~x18 && ~x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && x22 && ~x21 && ~x18 && ~x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && x22 && ~x21 && ~x18 && ~x19 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x22 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x22 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x22 && ~x4 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x21 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x65 && x21 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x65 && x21 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x21 && ~x9 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && x22 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && ~x22 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x70 && ~x65 && ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x70 && ~x65 && ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s253;
				s254 : if( x21 && x18 && x10 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( x21 && x18 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x21 && x18 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x21 && x18 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x21 && x18 && ~x10 && ~x4 )
						nx_state = s1;
					else if( x21 && ~x18 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x21 && ~x18 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x21 && ~x18 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x21 && ~x18 && ~x4 )
						nx_state = s1;
					else if( ~x21 && x22 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && x22 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x4 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x20 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && ~x22 && x20 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && ~x22 && x20 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x20 && ~x4 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x20 && x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && ~x22 && ~x20 && x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && ~x22 && ~x20 && x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x20 && x19 && ~x4 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x20 && ~x19 && x10 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x21 && ~x22 && ~x20 && ~x19 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && ~x22 && ~x20 && ~x19 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && ~x22 && ~x20 && ~x19 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x20 && ~x19 && ~x10 && ~x4 )
						nx_state = s1;
					else nx_state = s254;
				s255 : if( x70 && x2 )
						begin
							y5 = 1'b1;	
							nx_state = s945;
						end
					else if( x70 && ~x2 && x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x70 && ~x2 && ~x1 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x70 && x21 && x16 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x70 && x21 && x16 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s261;
						end
					else if( ~x70 && x21 && ~x16 && x17 && x18 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s1003;
						end
					else if( ~x70 && x21 && ~x16 && x17 && x18 && ~x3 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s810;
						end
					else if( ~x70 && x21 && ~x16 && x17 && x18 && ~x3 && ~x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( ~x70 && x21 && ~x16 && x17 && ~x18 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x70 && x21 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && ~x21 && x22 && x16 && x19 && x18 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && ~x21 && x22 && x16 && x19 && x18 && ~x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s264;
						end
					else if( ~x70 && ~x21 && x22 && x16 && x19 && ~x18 && x13 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x21 && x22 && x16 && x19 && ~x18 && ~x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && ~x21 && x22 && x16 && ~x19 && x13 )
						begin
							y3 = 1'b1;	y16 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && ~x21 && x22 && x16 && ~x19 && ~x13 && x18 && x15 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x21 && x22 && x16 && ~x19 && ~x13 && x18 && ~x15 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && ~x21 && x22 && x16 && ~x19 && ~x13 && ~x18 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && ~x21 && x22 && ~x16 && x17 && x18 && x19 && x10 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s1003;
						end
					else if( ~x70 && ~x21 && x22 && ~x16 && x17 && x18 && x19 && x10 && ~x3 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else if( ~x70 && ~x21 && x22 && ~x16 && x17 && x18 && x19 && ~x10 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && ~x21 && x22 && ~x16 && x17 && x18 && ~x19 && x13 && x3 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s1005;
						end
					else if( ~x70 && ~x21 && x22 && ~x16 && x17 && x18 && ~x19 && x13 && ~x3 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else if( ~x70 && ~x21 && x22 && ~x16 && x17 && x18 && ~x19 && ~x13 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && ~x21 && x22 && ~x16 && x17 && ~x18 && x13 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s1003;
						end
					else if( ~x70 && ~x21 && x22 && ~x16 && x17 && ~x18 && x13 && ~x3 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else if( ~x70 && ~x21 && x22 && ~x16 && x17 && ~x18 && ~x13 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && ~x21 && x22 && ~x16 && x17 && ~x18 && ~x13 && ~x19 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x70 && ~x21 && x22 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && ~x21 && ~x22 && x19 && x17 && x13 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x21 && ~x22 && x19 && x17 && ~x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && ~x21 && ~x22 && x19 && ~x17 && x18 && x13 && x3 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else if( ~x70 && ~x21 && ~x22 && x19 && ~x17 && x18 && x13 && ~x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s1003;
						end
					else if( ~x70 && ~x21 && ~x22 && x19 && ~x17 && x18 && ~x13 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x70 && ~x21 && ~x22 && x19 && ~x17 && ~x18 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x19 && x16 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x19 && x16 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s261;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x19 && ~x16 && x17 && x20 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x19 && ~x16 && x17 && ~x20 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s1003;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x19 && ~x16 && x17 && ~x20 && ~x3 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s810;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x19 && ~x16 && x17 && ~x20 && ~x3 && ~x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x19 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s252;
						end
					else nx_state = s255;
				s256 : if( x65 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x4 )
						nx_state = s1;
					else if( ~x65 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else nx_state = s256;
				s257 : if( x70 && x62 && x64 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x70 && x62 && x64 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x70 && x62 && x64 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x70 && x62 && x64 && ~x19 )
						nx_state = s1;
					else if( x70 && x62 && ~x64 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x70 && x62 && ~x64 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x70 && x62 && ~x64 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( x70 && x62 && ~x64 && ~x27 )
						nx_state = s1;
					else if( x70 && ~x62 && x63 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x70 && ~x62 && x63 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x70 && ~x62 && x63 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && x63 && ~x14 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && x66 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x66 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x66 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && x66 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && x67 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && x67 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && x67 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && x67 && ~x14 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x67 && x12 && x11 && x6 )
						begin
							y5 = 1'b1;	y27 = 1'b1;	y49 = 1'b1;	
							y50 = 1'b1;	
							nx_state = s1006;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x67 && x12 && x11 && ~x6 && x10 )
						begin
							y47 = 1'b1;	
							nx_state = s675;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x67 && x12 && x11 && ~x6 && ~x10 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y29 = 1'b1;	
							y35 = 1'b1;	y36 = 1'b1;	
							nx_state = s749;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x67 && x12 && ~x11 && x6 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y27 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s749;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x67 && x12 && ~x11 && ~x6 && x10 )
						begin
							y56 = 1'b1;	
							nx_state = s1007;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x67 && x12 && ~x11 && ~x6 && ~x10 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y28 = 1'b1;	
							y35 = 1'b1;	y36 = 1'b1;	
							nx_state = s749;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x67 && ~x12 && x11 && x6 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s1008;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x67 && ~x12 && x11 && ~x6 && x10 )
						begin
							y48 = 1'b1;	
							nx_state = s1009;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x67 && ~x12 && x11 && ~x6 && ~x10 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y30 = 1'b1;	
							y35 = 1'b1;	y36 = 1'b1;	
							nx_state = s749;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x67 && ~x12 && ~x11 && x6 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x67 && ~x12 && ~x11 && x6 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x67 && ~x12 && ~x11 && x6 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x67 && ~x12 && ~x11 && x6 && ~x18 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x67 && ~x12 && ~x11 && ~x6 && x10 )
						begin
							y54 = 1'b1;	
							nx_state = s525;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x67 && ~x12 && ~x11 && ~x6 && ~x10 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x67 && ~x12 && ~x11 && ~x6 && ~x10 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x67 && ~x12 && ~x11 && ~x6 && ~x10 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x66 && ~x67 && ~x12 && ~x11 && ~x6 && ~x10 && ~x18 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && x67 && x23 && x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x67 && x23 && x11 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x67 && x23 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && x67 && x23 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && x67 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x67 && x30 )
						begin
							y25 = 1'b1;	
							nx_state = s955;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x67 && ~x30 && x4 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x67 && ~x30 && x4 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x67 && ~x30 && x4 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x67 && ~x30 && x4 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x67 && ~x30 && ~x4 )
						begin
							y5 = 1'b1;	
							nx_state = s950;
						end
					else if( ~x70 && x65 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x4 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x67 && x24 && x26 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x67 && x24 && ~x26 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x65 && x67 && x24 && ~x26 && ~x4 && x19 && x16 && x11 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s368;
						end
					else if( ~x70 && ~x65 && x67 && x24 && ~x26 && ~x4 && x19 && x16 && x11 && ~x12 && x13 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( ~x70 && ~x65 && x67 && x24 && ~x26 && ~x4 && x19 && x16 && x11 && ~x12 && ~x13 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && ~x65 && x67 && x24 && ~x26 && ~x4 && x19 && x16 && ~x11 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s300;
						end
					else if( ~x70 && ~x65 && x67 && x24 && ~x26 && ~x4 && x19 && ~x16 && x17 && x11 && x13 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( ~x70 && ~x65 && x67 && x24 && ~x26 && ~x4 && x19 && ~x16 && x17 && x11 && ~x13 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s122;
						end
					else if( ~x70 && ~x65 && x67 && x24 && ~x26 && ~x4 && x19 && ~x16 && x17 && ~x11 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( ~x70 && ~x65 && x67 && x24 && ~x26 && ~x4 && x19 && ~x16 && ~x17 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && ~x65 && x67 && x24 && ~x26 && ~x4 && ~x19 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x70 && ~x65 && x67 && ~x24 && x25 && x26 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x70 && ~x65 && x67 && ~x24 && x25 && ~x26 && x15 && x10 && x11 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s433;
						end
					else if( ~x70 && ~x65 && x67 && ~x24 && x25 && ~x26 && x15 && x10 && ~x11 && x12 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s432;
						end
					else if( ~x70 && ~x65 && x67 && ~x24 && x25 && ~x26 && x15 && x10 && ~x11 && ~x12 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s300;
						end
					else if( ~x70 && ~x65 && x67 && ~x24 && x25 && ~x26 && x15 && ~x10 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s126;
						end
					else if( ~x70 && ~x65 && x67 && ~x24 && x25 && ~x26 && ~x15 && x16 && x10 && x12 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x70 && ~x65 && x67 && ~x24 && x25 && ~x26 && ~x15 && x16 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x70 && ~x65 && x67 && ~x24 && x25 && ~x26 && ~x15 && x16 && ~x10 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x70 && ~x65 && x67 && ~x24 && x25 && ~x26 && ~x15 && ~x16 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( ~x70 && ~x65 && x67 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x67 && x21 && x9 && x3 )
						nx_state = s47;
					else if( ~x70 && ~x65 && ~x67 && x21 && x9 && ~x3 && x4 )
						nx_state = s47;
					else if( ~x70 && ~x65 && ~x67 && x21 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x67 && x21 && ~x9 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x67 && ~x21 && x22 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x65 && ~x67 && ~x21 && x22 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x65 && ~x67 && ~x21 && x22 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x67 && ~x21 && x22 && ~x5 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x67 && ~x21 && ~x22 )
						nx_state = s1;
					else nx_state = s257;
				s258 : if( x65 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x4 )
						nx_state = s1;
					else if( ~x65 && x24 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( ~x65 && ~x24 && x15 && x10 && x11 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s433;
						end
					else if( ~x65 && ~x24 && x15 && x10 && ~x11 && x12 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s432;
						end
					else if( ~x65 && ~x24 && x15 && x10 && ~x11 && ~x12 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s300;
						end
					else if( ~x65 && ~x24 && x15 && ~x10 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s126;
						end
					else if( ~x65 && ~x24 && ~x15 && x16 && x10 && x12 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s497;
						end
					else if( ~x65 && ~x24 && ~x15 && x16 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x65 && ~x24 && ~x15 && x16 && ~x10 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s497;
						end
					else if( ~x65 && ~x24 && ~x15 && ~x16 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else nx_state = s258;
				s259 : if( x70 && x64 && x12 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y32 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s749;
						end
					else if( x70 && x64 && ~x12 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x70 && x64 && ~x12 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x70 && x64 && ~x12 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x70 && x64 && ~x12 && ~x18 )
						nx_state = s1;
					else if( x70 && ~x64 )
						begin
							y25 = 1'b1;	
							nx_state = s1010;
						end
					else if( ~x70 && x67 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x67 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x67 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x67 && ~x4 )
						nx_state = s1;
					else if( ~x70 && ~x67 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x67 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x67 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x70 && ~x67 && ~x5 )
						nx_state = s1;
					else nx_state = s259;
				s260 : if( x69 && x21 && x66 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x21 && x66 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x21 && x66 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && x21 && x66 && x20 && ~x17 )
						nx_state = s1;
					else if( x69 && x21 && x66 && ~x20 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( x69 && x21 && ~x66 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x21 && ~x66 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x21 && ~x66 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && x21 && ~x66 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x21 && x66 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x21 && ~x66 && x22 && x18 && x19 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x21 && ~x66 && x22 && x18 && x19 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x21 && ~x66 && x22 && x18 && x19 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x21 && ~x66 && x22 && x18 && ~x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x21 && ~x66 && x22 && x18 && ~x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x21 && ~x66 && x22 && x18 && ~x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x21 && ~x66 && x22 && x18 && ~x19 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x21 && ~x66 && x22 && ~x18 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x21 && ~x66 && x22 && ~x18 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x21 && ~x66 && x22 && ~x18 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x21 && ~x66 && x22 && ~x18 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x21 && ~x66 && ~x22 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x21 && ~x66 && ~x22 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && ~x21 && ~x66 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x21 && ~x66 && ~x22 && ~x4 )
						nx_state = s1;
					else if( ~x69 && x10 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s215;
						end
					else if( ~x69 && ~x10 && x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x69 && ~x10 && ~x7 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s280;
						end
					else nx_state = s260;
				s261 : if( x21 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x21 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x21 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x21 && ~x4 )
						nx_state = s1;
					else if( ~x21 && x22 && x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && x22 && x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && x22 && x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && x19 && ~x4 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x18 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && x22 && ~x19 && x18 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && x22 && ~x19 && x18 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x18 && ~x4 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && ~x18 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( ~x21 && ~x22 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s261;
				s262 : if( x70 && x62 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x70 && x62 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x70 && x62 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x70 && x62 && ~x19 )
						nx_state = s1;
					else if( x70 && ~x62 && x64 && x63 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( x70 && ~x62 && x64 && ~x63 && x67 )
						begin
							y5 = 1'b1;	y13 = 1'b1;	y17 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1011;
						end
					else if( x70 && ~x62 && x64 && ~x63 && ~x67 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && x64 && ~x63 && ~x67 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && x64 && ~x63 && ~x67 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && x64 && ~x63 && ~x67 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x64 && x63 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x70 && ~x62 && ~x64 && x63 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x70 && ~x62 && ~x64 && x63 && x19 && ~x14 && ~x13 && x11 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( x70 && ~x62 && ~x64 && x63 && x19 && ~x14 && ~x13 && x11 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( x70 && ~x62 && ~x64 && x63 && x19 && ~x14 && ~x13 && ~x11 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( x70 && ~x62 && ~x64 && x63 && ~x19 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x64 && ~x63 && x65 && x67 && x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x62 && ~x64 && ~x63 && x65 && x67 && x11 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x62 && ~x64 && ~x63 && x65 && x67 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x64 && ~x63 && x65 && x67 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x64 && ~x63 && x65 && ~x67 )
						begin
							y24 = 1'b1;	
							nx_state = s1012;
						end
					else if( x70 && ~x62 && ~x64 && ~x63 && ~x65 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x62 && ~x64 && ~x63 && ~x65 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x62 && ~x64 && ~x63 && ~x65 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x64 && ~x63 && ~x65 && ~x17 )
						nx_state = s1;
					else if( ~x70 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && ~x4 )
						nx_state = s1;
					else nx_state = s262;
				s263 : if( x70 && x11 )
						begin
							y1 = 1'b1;	y22 = 1'b1;	
							nx_state = s1013;
						end
					else if( x70 && ~x11 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && x22 && x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x22 && x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x22 && x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x22 && x19 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x22 && ~x19 && x18 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x22 && ~x19 && x18 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x22 && ~x19 && x18 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x22 && ~x19 && x18 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x22 && ~x19 && ~x18 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && ~x22 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && ~x22 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s263;
				s264 : if( x22 && x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x22 && x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x22 && x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x22 && x19 && ~x4 )
						nx_state = s1;
					else if( x22 && ~x19 && x18 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( x22 && ~x19 && ~x18 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x22 && ~x19 && ~x18 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x22 && ~x19 && ~x18 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x22 && ~x19 && ~x18 && ~x4 )
						nx_state = s1;
					else if( ~x22 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x22 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s264;
				s265 : if( x70 && x63 && x20 && x21 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s1014;
						end
					else if( x70 && x63 && x20 && ~x21 )
						begin
							y6 = 1'b1;	y42 = 1'b1;	y43 = 1'b1;	
							nx_state = s1015;
						end
					else if( x70 && x63 && ~x20 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1016;
						end
					else if( x70 && ~x63 && x67 && x23 )
						begin
							y29 = 1'b1;	
							nx_state = s1017;
						end
					else if( x70 && ~x63 && x67 && ~x23 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x70 && ~x63 && x67 && ~x23 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x70 && ~x63 && x67 && ~x23 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x70 && ~x63 && x67 && ~x23 && ~x20 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x67 && x29 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x63 && ~x67 && x29 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x63 && ~x67 && x29 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x67 && x29 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x67 && ~x29 )
						begin
							y8 = 1'b1;	
							nx_state = s744;
						end
					else if( ~x70 && x65 && x67 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && x67 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && x67 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && x65 && x67 && ~x4 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x67 && x21 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x70 && x65 && ~x67 && ~x21 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x70 && ~x65 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s253;
						end
					else nx_state = s265;
				s266 : if( x70 && x62 && x64 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1018;
						end
					else if( x70 && x62 && ~x64 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y37 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s1019;
						end
					else if( x70 && ~x62 && x63 && x13 && x67 && x11 && x14 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x70 && ~x62 && x63 && x13 && x67 && x11 && ~x14 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s577;
						end
					else if( x70 && ~x62 && x63 && x13 && x67 && ~x11 && x10 && x14 && x3 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s66;
						end
					else if( x70 && ~x62 && x63 && x13 && x67 && ~x11 && x10 && x14 && x3 && ~x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x70 && ~x62 && x63 && x13 && x67 && ~x11 && x10 && x14 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x70 && ~x62 && x63 && x13 && x67 && ~x11 && x10 && ~x14 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s65;
						end
					else if( x70 && ~x62 && x63 && x13 && x67 && ~x11 && x10 && ~x14 && ~x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x70 && ~x62 && x63 && x13 && x67 && ~x11 && ~x10 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x70 && ~x62 && x63 && x13 && x67 && ~x11 && ~x10 && ~x1 && x3 )
						nx_state = s1;
					else if( x70 && ~x62 && x63 && x13 && x67 && ~x11 && ~x10 && ~x1 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x70 && ~x62 && x63 && x13 && ~x67 && x15 && x14 && x10 && x3 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s66;
						end
					else if( x70 && ~x62 && x63 && x13 && ~x67 && x15 && x14 && x10 && x3 && ~x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x70 && ~x62 && x63 && x13 && ~x67 && x15 && x14 && x10 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x70 && ~x62 && x63 && x13 && ~x67 && x15 && x14 && ~x10 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x70 && ~x62 && x63 && x13 && ~x67 && x15 && ~x14 && x10 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s65;
						end
					else if( x70 && ~x62 && x63 && x13 && ~x67 && x15 && ~x14 && x10 && ~x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x70 && ~x62 && x63 && x13 && ~x67 && x15 && ~x14 && ~x10 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s577;
						end
					else if( x70 && ~x62 && x63 && x13 && ~x67 && ~x15 && x11 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && ~x62 && x63 && x13 && ~x67 && ~x15 && x11 && ~x3 && x5 && x7 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x70 && ~x62 && x63 && x13 && ~x67 && ~x15 && x11 && ~x3 && x5 && ~x7 )
						nx_state = s266;
					else if( x70 && ~x62 && x63 && x13 && ~x67 && ~x15 && x11 && ~x3 && ~x5 && x12 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x70 && ~x62 && x63 && x13 && ~x67 && ~x15 && x11 && ~x3 && ~x5 && ~x12 )
						nx_state = s266;
					else if( x70 && ~x62 && x63 && x13 && ~x67 && ~x15 && ~x11 && x10 && x5 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x70 && ~x62 && x63 && x13 && ~x67 && ~x15 && ~x11 && x10 && ~x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x70 && ~x62 && x63 && x13 && ~x67 && ~x15 && ~x11 && ~x10 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( x70 && ~x62 && x63 && x13 && ~x67 && ~x15 && ~x11 && ~x10 && ~x1 && x3 )
						nx_state = s1;
					else if( x70 && ~x62 && x63 && x13 && ~x67 && ~x15 && ~x11 && ~x10 && ~x1 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x70 && ~x62 && x63 && ~x13 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && ~x62 && x63 && ~x13 && ~x3 && x5 && x7 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x70 && ~x62 && x63 && ~x13 && ~x3 && x5 && ~x7 )
						nx_state = s266;
					else if( x70 && ~x62 && x63 && ~x13 && ~x3 && ~x5 && x12 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( x70 && ~x62 && x63 && ~x13 && ~x3 && ~x5 && ~x12 )
						nx_state = s266;
					else if( x70 && ~x62 && ~x63 && x64 && x21 && x20 )
						begin
							y6 = 1'b1;	
							nx_state = s431;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x21 && ~x20 )
						begin
							y6 = 1'b1;	
							nx_state = s659;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x21 )
						begin
							y6 = 1'b1;	
							nx_state = s431;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 )
						begin
							y47 = 1'b1;	y51 = 1'b1;	y61 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s878;
						end
					else if( ~x70 && x68 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x68 && x21 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x68 && ~x21 && x22 && x23 && x15 && x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && ~x68 && ~x21 && x22 && x23 && x15 && ~x10 && x12 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && ~x68 && ~x21 && x22 && x23 && x15 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s366;
						end
					else if( ~x70 && ~x68 && ~x21 && x22 && x23 && ~x15 && x16 && x10 && x12 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x70 && ~x68 && ~x21 && x22 && x23 && ~x15 && x16 && x10 && ~x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x70 && ~x68 && ~x21 && x22 && x23 && ~x15 && x16 && ~x10 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x70 && ~x68 && ~x21 && x22 && x23 && ~x15 && ~x16 )
						nx_state = s47;
					else if( ~x70 && ~x68 && ~x21 && x22 && ~x23 && x6 && x15 && x11 && x10 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x70 && ~x68 && ~x21 && x22 && ~x23 && x6 && x15 && x11 && ~x10 )
						begin
							y14 = 1'b1;	
							nx_state = s366;
						end
					else if( ~x70 && ~x68 && ~x21 && x22 && ~x23 && x6 && x15 && ~x11 && x12 && x10 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x70 && ~x68 && ~x21 && x22 && ~x23 && x6 && x15 && ~x11 && x12 && ~x10 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && ~x68 && ~x21 && x22 && ~x23 && x6 && x15 && ~x11 && ~x12 && x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && ~x68 && ~x21 && x22 && ~x23 && x6 && x15 && ~x11 && ~x12 && ~x10 )
						begin
							y14 = 1'b1;	
							nx_state = s366;
						end
					else if( ~x70 && ~x68 && ~x21 && x22 && ~x23 && x6 && ~x15 && x16 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && ~x68 && ~x21 && x22 && ~x23 && x6 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s362;
						end
					else if( ~x70 && ~x68 && ~x21 && x22 && ~x23 && ~x6 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && ~x68 && ~x21 && ~x22 && x23 && x15 && x7 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s151;
						end
					else if( ~x70 && ~x68 && ~x21 && ~x22 && x23 && x15 && ~x7 && x9 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x68 && ~x21 && ~x22 && x23 && x15 && ~x7 && ~x9 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x68 && ~x21 && ~x22 && x23 && ~x15 && x16 && x7 && x9 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x68 && ~x21 && ~x22 && x23 && ~x15 && x16 && x7 && ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && ~x68 && ~x21 && ~x22 && x23 && ~x15 && x16 && ~x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x68 && ~x21 && ~x22 && x23 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( ~x70 && ~x68 && ~x21 && ~x22 && ~x23 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s151;
						end
					else nx_state = s266;
				s267 : if( x21 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x21 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x21 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x21 && ~x9 )
						nx_state = s1;
					else if( ~x21 && x22 && x8 && x7 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x21 && x22 && x8 && ~x7 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s267;
				s268 : if( x21 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x21 && x22 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x21 && ~x22 )
						begin
							y2 = 1'b1;	y16 = 1'b1;	y24 = 1'b1;	
							nx_state = s270;
						end
					else nx_state = s268;
				s269 : if( 1'b1 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s565;
						end
					else nx_state = s269;
				s270 : if( x65 && x22 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( x65 && ~x22 && ~x23 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s1020;
						end
					else if( ~x65 && x21 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x65 && x21 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x65 && x21 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && x21 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x21 && x22 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x21 && x22 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x7 )
						nx_state = s1;
					else if( ~x65 && ~x21 && ~x22 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x65 && ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x65 && ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s270;
				s271 : if( x70 && x64 && x65 )
						begin
							y6 = 1'b1;	
							nx_state = s431;
						end
					else if( x70 && x64 && ~x65 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y13 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1021;
						end
					else if( x70 && ~x64 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x70 && ~x64 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x70 && ~x64 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x64 && ~x8 )
						nx_state = s1;
					else if( ~x70 && x66 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x70 && ~x66 && x24 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( ~x70 && ~x66 && ~x24 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else nx_state = s271;
				s272 : if( x69 && x66 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x69 && ~x66 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( ~x69 )
						begin
							y8 = 1'b1;	y12 = 1'b1;	
							nx_state = s879;
						end
					else nx_state = s272;
				s273 : if( x21 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x21 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x21 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x21 && ~x9 )
						nx_state = s1;
					else if( ~x21 && x22 )
						nx_state = s1;
					else if( ~x21 && ~x22 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else nx_state = s273;
				s274 : if( x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x18 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x21 && x22 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x21 && x22 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x17 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && x18 && x14 )
						nx_state = s47;
					else if( ~x21 && x22 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s47;
					else if( ~x21 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && x7 && x9 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x23 && x7 && x9 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x23 && x7 && x9 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && x7 && x9 && ~x19 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && x7 && ~x9 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s275;
						end
					else if( ~x21 && ~x22 && x23 && ~x7 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x23 && ~x7 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x23 && ~x7 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x7 && ~x19 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else nx_state = s274;
				s275 : if( x21 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( ~x21 && x22 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x21 && x22 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x21 && x22 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x17 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x19 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 )
						begin
							y3 = 1'b1;	
							nx_state = s835;
						end
					else nx_state = s275;
				s276 : if( x62 && x6 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x62 && ~x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x62 && x15 )
						nx_state = s1;
					else if( ~x62 && ~x15 && x6 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x62 && ~x15 && ~x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else nx_state = s276;
				s277 : if( x62 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x62 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x62 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( x62 && ~x21 )
						nx_state = s1;
					else if( ~x62 && x64 && x63 && x65 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x62 && x64 && x63 && x65 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x62 && x64 && x63 && x65 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x62 && x64 && x63 && x65 && ~x11 )
						nx_state = s1;
					else if( ~x62 && x64 && x63 && ~x65 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x62 && x64 && x63 && ~x65 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x62 && x64 && x63 && ~x65 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x62 && x64 && x63 && ~x65 && ~x14 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x63 && x65 && x6 && x3 && x7 && x9 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && x3 && x7 && ~x9 )
						begin
							y29 = 1'b1;	
							nx_state = s771;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && x3 && ~x7 && x8 && x9 && x11 )
						begin
							y3 = 1'b1;	
							nx_state = s789;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && x3 && ~x7 && x8 && x9 && ~x11 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && x3 && ~x7 && x8 && x9 && ~x11 && x14 && ~x10 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x63 && x65 && x6 && x3 && ~x7 && x8 && x9 && ~x11 && ~x14 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x63 && x65 && x6 && x3 && ~x7 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s789;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && x3 && ~x7 && x8 && ~x9 && ~x10 && x14 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && x3 && ~x7 && x8 && ~x9 && ~x10 && x14 && ~x11 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x63 && x65 && x6 && x3 && ~x7 && x8 && ~x9 && ~x10 && ~x14 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x63 && x65 && x6 && x3 && ~x7 && ~x8 && x9 )
						begin
							y32 = 1'b1;	y33 = 1'b1;	
							nx_state = s396;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && x3 && ~x7 && ~x8 && ~x9 )
						begin
							y30 = 1'b1;	y31 = 1'b1;	
							nx_state = s1022;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && x8 && x9 && x15 && x16 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && x8 && x9 && x15 && x16 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && x8 && x9 && x15 && x16 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && x8 && x9 && x15 && x16 && ~x14 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && x8 && x9 && x15 && ~x16 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && x8 && x9 && ~x15 && x7 )
						begin
							y16 = 1'b1;	
							nx_state = s293;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && x8 && x9 && ~x15 && ~x7 )
						begin
							y25 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s1023;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && x8 && ~x9 && x15 && x17 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && x8 && ~x9 && x15 && ~x17 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && x8 && ~x9 && x15 && ~x17 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && x8 && ~x9 && x15 && ~x17 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && x8 && ~x9 && x15 && ~x17 && ~x14 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && x8 && ~x9 && ~x15 && x7 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && x8 && ~x9 && ~x15 && ~x7 )
						begin
							y22 = 1'b1;	y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s1024;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && ~x8 && x9 && x15 && x18 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && ~x8 && x9 && x15 && ~x18 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && ~x8 && x9 && x15 && ~x18 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && ~x8 && x9 && x15 && ~x18 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && ~x8 && x9 && x15 && ~x18 && ~x14 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && ~x8 && x9 && ~x15 && x7 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && ~x8 && x9 && ~x15 && ~x7 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && ~x8 && ~x9 && x15 && x18 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && ~x8 && ~x9 && x15 && x18 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && ~x8 && ~x9 && x15 && x18 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && ~x8 && ~x9 && x15 && x18 && ~x14 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && ~x8 && ~x9 && x15 && ~x18 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && ~x8 && ~x9 && ~x15 && x7 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x62 && x64 && ~x63 && x65 && x6 && ~x3 && ~x8 && ~x9 && ~x15 && ~x7 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( ~x62 && x64 && ~x63 && x65 && ~x6 && x3 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x62 && x64 && ~x63 && x65 && ~x6 && ~x3 && x12 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s560;
						end
					else if( ~x62 && x64 && ~x63 && x65 && ~x6 && ~x3 && x12 && ~x4 && x5 )
						begin
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s561;
						end
					else if( ~x62 && x64 && ~x63 && x65 && ~x6 && ~x3 && x12 && ~x4 && ~x5 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else if( ~x62 && x64 && ~x63 && x65 && ~x6 && ~x3 && ~x12 && x4 && x5 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x62 && x64 && ~x63 && x65 && ~x6 && ~x3 && ~x12 && x4 && ~x5 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x62 && x64 && ~x63 && x65 && ~x6 && ~x3 && ~x12 && ~x4 )
						begin
							y5 = 1'b1;	
							nx_state = s562;
						end
					else if( ~x62 && x64 && ~x63 && ~x65 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x62 && x64 && ~x63 && ~x65 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x62 && x64 && ~x63 && ~x65 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x63 && ~x65 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x63 && ~x65 && ~x22 )
						nx_state = s1;
					else if( ~x62 && ~x64 && x63 && x16 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x62 && ~x64 && x63 && x16 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x62 && ~x64 && x63 && x16 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x62 && ~x64 && x63 && ~x16 )
						nx_state = s1;
					else if( ~x62 && ~x64 && ~x63 && x65 )
						begin
							y35 = 1'b1;	
							nx_state = s1025;
						end
					else if( ~x62 && ~x64 && ~x63 && ~x65 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x62 && ~x64 && ~x63 && ~x65 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x62 && ~x64 && ~x63 && ~x65 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x62 && ~x64 && ~x63 && ~x65 && ~x8 )
						nx_state = s1;
					else nx_state = s277;
				s278 : if( 1'b1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else nx_state = s278;
				s279 : if( x70 && x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s255;
						end
					else if( x70 && ~x2 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x70 && x67 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x67 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x67 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x67 && x22 && ~x17 )
						nx_state = s1;
					else if( ~x70 && x67 && ~x22 && x18 && x13 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && x67 && ~x22 && x18 && x13 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x67 && ~x22 && x18 && ~x13 && x12 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && x67 && ~x22 && x18 && ~x13 && x12 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x67 && ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && x67 && ~x22 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x67 && x61 && x60 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x70 && ~x67 && x61 && ~x60 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && ~x67 && x61 && ~x60 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && ~x67 && x61 && ~x60 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( ~x70 && ~x67 && x61 && ~x60 && x62 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x67 && x61 && ~x60 && ~x62 && x15 )
						nx_state = s143;
					else if( ~x70 && ~x67 && x61 && ~x60 && ~x62 && ~x15 && x16 )
						begin
							y12 = 1'b1;	
							nx_state = s244;
						end
					else if( ~x70 && ~x67 && x61 && ~x60 && ~x62 && ~x15 && ~x16 )
						nx_state = s143;
					else if( ~x70 && ~x67 && ~x61 && x60 && x15 )
						nx_state = s143;
					else if( ~x70 && ~x67 && ~x61 && x60 && ~x15 && x16 )
						begin
							y12 = 1'b1;	
							nx_state = s244;
						end
					else if( ~x70 && ~x67 && ~x61 && x60 && ~x15 && ~x16 )
						nx_state = s143;
					else if( ~x70 && ~x67 && ~x61 && ~x60 && x62 )
						nx_state = s1;
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && x15 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && x15 && ~x7 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && x15 && ~x7 && ~x11 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && x4 )
						nx_state = s47;
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && ~x4 && x11 && x9 )
						nx_state = s47;
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && ~x4 && x11 && ~x9 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && ~x4 && x11 && ~x9 && ~x7 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s559;
						end
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && ~x4 && ~x11 && x9 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && ~x4 && ~x11 && x9 && ~x7 && x10 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && ~x4 && ~x11 && x9 && ~x7 && ~x10 )
						nx_state = s47;
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && x7 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && x7 && ~x8 )
						nx_state = s47;
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && ~x7 && x12 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && ~x7 && ~x12 )
						nx_state = s47;
					else if( ~x70 && ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else nx_state = s279;
				s280 : if( x69 && x17 && x18 && x6 && x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( x69 && x17 && x18 && x6 && ~x9 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	
							nx_state = s20;
						end
					else if( x69 && x17 && x18 && ~x6 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s215;
						end
					else if( x69 && x17 && ~x18 && x10 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && x17 && ~x18 && ~x10 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x69 && ~x17 && x8 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	
							nx_state = s20;
						end
					else if( x69 && ~x17 && ~x8 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s320;
						end
					else if( ~x69 && x70 && x62 && x16 && x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( ~x69 && x70 && x62 && x16 && ~x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && x70 && x62 && ~x16 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s215;
						end
					else if( ~x69 && x70 && ~x62 && x64 && x63 && x47 && x9 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	y34 = 1'b1;	
							nx_state = s904;
						end
					else if( ~x69 && x70 && ~x62 && x64 && x63 && x47 && ~x9 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s739;
						end
					else if( ~x69 && x70 && ~x62 && x64 && x63 && ~x47 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( ~x69 && x70 && ~x62 && x64 && ~x63 && x16 && x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( ~x69 && x70 && ~x62 && x64 && ~x63 && x16 && ~x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && x70 && ~x62 && x64 && ~x63 && ~x16 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( ~x69 && x70 && ~x62 && ~x64 && x16 && x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( ~x69 && x70 && ~x62 && ~x64 && x16 && ~x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && x70 && ~x62 && ~x64 && ~x16 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x10 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x10 && x11 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x10 && x11 && ~x1 && x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x10 && x11 && ~x1 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x10 && ~x11 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x16 && x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x16 && ~x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x16 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( ~x69 && ~x70 && ~x44 && x10 && x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && ~x70 && ~x44 && x10 && ~x8 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s320;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 && x6 && x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 && x6 && ~x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 && ~x6 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s215;
						end
					else nx_state = s280;
				s281 : if( x63 && x21 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x63 && x21 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x63 && x21 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x63 && x21 && ~x10 )
						nx_state = s1;
					else if( x63 && ~x21 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x63 && x65 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1026;
						end
					else if( ~x63 && ~x65 && x66 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && ~x65 && x66 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && ~x65 && x66 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x63 && ~x65 && x66 && ~x9 )
						nx_state = s1;
					else if( ~x63 && ~x65 && ~x66 )
						begin
							y53 = 1'b1;	
							nx_state = s1027;
						end
					else nx_state = s281;
				s282 : if( x63 && x16 )
						begin
							y47 = 1'b1;	y48 = 1'b1;	
							nx_state = s1028;
						end
					else if( x63 && ~x16 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x63 && ~x16 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x63 && ~x16 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x63 && ~x16 && ~x10 )
						nx_state = s1;
					else if( ~x63 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x63 && ~x9 )
						nx_state = s1;
					else nx_state = s282;
				s283 : if( x65 )
						begin
							y4 = 1'b1;	y20 = 1'b1;	y31 = 1'b1;	
							nx_state = s1029;
						end
					else if( ~x65 && x66 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x66 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x65 && x66 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x66 )
						nx_state = s1;
					else nx_state = s283;
				s284 : if( x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x9 )
						nx_state = s1;
					else nx_state = s284;
				s285 : if( x62 && x33 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s979;
						end
					else if( x62 && ~x33 && x32 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s979;
						end
					else if( x62 && ~x33 && ~x32 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x62 && ~x33 && ~x32 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x62 && ~x33 && ~x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x62 && ~x33 && ~x32 && ~x10 )
						nx_state = s1;
					else if( ~x62 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x62 && ~x9 )
						nx_state = s1;
					else nx_state = s285;
				s286 : if( x62 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x62 && ~x14 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x62 && ~x14 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x62 && ~x14 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( x62 && ~x14 && ~x21 )
						nx_state = s1;
					else if( ~x62 && x63 && x64 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x62 && x63 && x64 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x62 && x63 && x64 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x62 && x63 && x64 && ~x11 )
						nx_state = s1;
					else if( ~x62 && x63 && ~x64 && x65 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x62 && x63 && ~x64 && x65 && ~x18 )
						begin
							y44 = 1'b1;	
							nx_state = s755;
						end
					else if( ~x62 && x63 && ~x64 && ~x65 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x62 && x63 && ~x64 && ~x65 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x62 && x63 && ~x64 && ~x65 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x62 && x63 && ~x64 && ~x65 && ~x1 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x13 )
						begin
							y46 = 1'b1;	
							nx_state = s1030;
						end
					else if( ~x62 && ~x63 && ~x13 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && ~x63 && ~x13 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && ~x63 && ~x13 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x13 && ~x9 )
						nx_state = s1;
					else nx_state = s286;
				s287 : if( x63 && x64 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x63 && x64 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x63 && x64 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x63 && x64 && ~x11 )
						nx_state = s1;
					else if( x63 && ~x64 && x67 )
						begin
							y3 = 1'b1;	y18 = 1'b1;	y52 = 1'b1;	
							nx_state = s1031;
						end
					else if( x63 && ~x64 && ~x67 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x64 && ~x67 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x64 && ~x67 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x63 && ~x64 && ~x67 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x64 && ~x67 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x63 && x66 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x66 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x66 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x63 && x66 && ~x9 )
						nx_state = s1;
					else if( ~x63 && ~x66 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x63 && ~x66 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x63 && ~x66 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( ~x63 && ~x66 && ~x14 )
						nx_state = s1;
					else nx_state = s287;
				s288 : if( x69 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && ~x9 )
						nx_state = s1;
					else if( ~x69 )
						begin
							y3 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s1032;
						end
					else nx_state = s288;
				s289 : if( x63 && x64 && x65 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x63 && x64 && x65 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x63 && x64 && x65 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( x63 && x64 && x65 && ~x22 )
						nx_state = s1;
					else if( x63 && x64 && ~x65 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x63 && x64 && ~x65 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x63 && x64 && ~x65 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x63 && x64 && ~x65 && ~x14 )
						nx_state = s1;
					else if( x63 && ~x64 && x65 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x63 && ~x64 && x65 && ~x15 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x63 && ~x64 && ~x65 )
						nx_state = s1;
					else if( ~x63 && x64 && x65 )
						begin
							y15 = 1'b1;	
							nx_state = s243;
						end
					else if( ~x63 && x64 && ~x65 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x64 && ~x65 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x64 && ~x65 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x63 && x64 && ~x65 && ~x9 )
						nx_state = s1;
					else if( ~x63 && ~x64 && x19 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( ~x63 && ~x64 && ~x19 && x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x64 && ~x19 && x26 && ~x25 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x64 && ~x19 && x26 && ~x25 && ~x24 )
						nx_state = s1;
					else if( ~x63 && ~x64 && ~x19 && ~x26 )
						nx_state = s1;
					else nx_state = s289;
				s290 : if( x64 && x62 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x64 && x62 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x64 && x62 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x64 && x62 && ~x19 )
						nx_state = s1;
					else if( x64 && ~x62 && x63 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x64 && ~x62 && x63 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x64 && ~x62 && x63 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x64 && ~x62 && x63 && ~x14 )
						nx_state = s1;
					else if( x64 && ~x62 && ~x63 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x64 && ~x62 && ~x63 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x64 && ~x62 && ~x63 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x64 && ~x62 && ~x63 && ~x9 )
						nx_state = s1;
					else if( ~x64 && x62 )
						nx_state = s1;
					else if( ~x64 && ~x62 && x65 && x63 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x64 && ~x62 && x65 && ~x63 )
						begin
							y31 = 1'b1;	
							nx_state = s886;
						end
					else if( ~x64 && ~x62 && ~x65 && x63 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x64 && ~x62 && ~x65 && x63 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x64 && ~x62 && ~x65 && x63 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x64 && ~x62 && ~x65 && x63 && ~x1 )
						nx_state = s1;
					else if( ~x64 && ~x62 && ~x65 && ~x63 && x66 && x21 && x22 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x64 && ~x62 && ~x65 && ~x63 && x66 && x21 && ~x22 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x64 && ~x62 && ~x65 && ~x63 && x66 && x21 && ~x22 && ~x23 )
						nx_state = s1;
					else if( ~x64 && ~x62 && ~x65 && ~x63 && x66 && ~x21 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x64 && ~x62 && ~x65 && ~x63 && x66 && ~x21 && ~x23 )
						nx_state = s1;
					else if( ~x64 && ~x62 && ~x65 && ~x63 && ~x66 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( ~x64 && ~x62 && ~x65 && ~x63 && ~x66 && ~x18 && x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x64 && ~x62 && ~x65 && ~x63 && ~x66 && ~x18 && x26 && ~x25 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x64 && ~x62 && ~x65 && ~x63 && ~x66 && ~x18 && x26 && ~x25 && ~x24 )
						nx_state = s1;
					else if( ~x64 && ~x62 && ~x65 && ~x63 && ~x66 && ~x18 && ~x26 )
						nx_state = s1;
					else nx_state = s290;
				s291 : if( x62 && x64 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x62 && x64 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x62 && x64 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( x62 && x64 && ~x21 )
						nx_state = s1;
					else if( x62 && ~x64 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x62 && ~x64 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x62 && ~x64 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( x62 && ~x64 && ~x27 )
						nx_state = s1;
					else if( ~x62 && x63 && x66 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x62 && x63 && ~x66 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( ~x62 && x63 && ~x66 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( ~x62 && x63 && ~x66 && x19 && ~x14 && ~x13 && x11 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( ~x62 && x63 && ~x66 && x19 && ~x14 && ~x13 && x11 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x62 && x63 && ~x66 && x19 && ~x14 && ~x13 && ~x11 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x62 && x63 && ~x66 && ~x19 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && ~x63 && x64 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && ~x63 && x64 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && ~x9 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 && x65 && x67 && x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x62 && ~x63 && ~x64 && x65 && x67 && x11 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x62 && ~x63 && ~x64 && x65 && x67 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 && x65 && x67 && ~x11 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 && x65 && ~x67 )
						begin
							y33 = 1'b1;	
							nx_state = s1033;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x66 && x21 && x22 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x66 && x21 && ~x22 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x66 && x21 && ~x22 && ~x23 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x66 && ~x21 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x66 && ~x21 && ~x23 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 && ~x65 && ~x66 && x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && ~x66 && x26 && ~x25 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && ~x66 && x26 && ~x25 && ~x24 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 && ~x65 && ~x66 && ~x26 )
						nx_state = s1;
					else nx_state = s291;
				s292 : if( x62 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x62 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x62 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( x62 && ~x21 )
						nx_state = s1;
					else if( ~x62 && x65 && x64 && x63 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x62 && x65 && x64 && x63 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x62 && x65 && x64 && x63 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( ~x62 && x65 && x64 && x63 && ~x22 )
						nx_state = s1;
					else if( ~x62 && x65 && x64 && ~x63 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x62 && x65 && ~x64 && x63 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x62 && x65 && ~x64 && ~x63 && x67 )
						nx_state = s1;
					else if( ~x62 && x65 && ~x64 && ~x63 && ~x67 && x4 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x62 && x65 && ~x64 && ~x63 && ~x67 && x4 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x62 && x65 && ~x64 && ~x63 && ~x67 && x4 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x62 && x65 && ~x64 && ~x63 && ~x67 && x4 && ~x23 )
						nx_state = s1;
					else if( ~x62 && x65 && ~x64 && ~x63 && ~x67 && ~x4 )
						begin
							y5 = 1'b1;	
							nx_state = s945;
						end
					else if( ~x62 && ~x65 && x63 )
						nx_state = s1;
					else if( ~x62 && ~x65 && ~x63 && x64 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && ~x65 && ~x63 && x64 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && ~x65 && ~x63 && x64 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x62 && ~x65 && ~x63 && x64 && ~x9 )
						nx_state = s1;
					else if( ~x62 && ~x65 && ~x63 && ~x64 && x66 && x21 && x22 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x62 && ~x65 && ~x63 && ~x64 && x66 && x21 && ~x22 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x62 && ~x65 && ~x63 && ~x64 && x66 && x21 && ~x22 && ~x23 )
						nx_state = s1;
					else if( ~x62 && ~x65 && ~x63 && ~x64 && x66 && ~x21 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x62 && ~x65 && ~x63 && ~x64 && x66 && ~x21 && ~x23 )
						nx_state = s1;
					else if( ~x62 && ~x65 && ~x63 && ~x64 && ~x66 && x20 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( ~x62 && ~x65 && ~x63 && ~x64 && ~x66 && ~x20 && x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x62 && ~x65 && ~x63 && ~x64 && ~x66 && ~x20 && x26 && ~x25 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x62 && ~x65 && ~x63 && ~x64 && ~x66 && ~x20 && x26 && ~x25 && ~x24 )
						nx_state = s1;
					else if( ~x62 && ~x65 && ~x63 && ~x64 && ~x66 && ~x20 && ~x26 )
						nx_state = s1;
					else nx_state = s292;
				s293 : if( x62 && x13 && x4 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	
							nx_state = s231;
						end
					else if( x62 && x13 && ~x4 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x62 && ~x13 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s230;
						end
					else if( x62 && ~x13 && ~x14 && x9 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s230;
						end
					else if( x62 && ~x13 && ~x14 && ~x9 && x7 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s230;
						end
					else if( x62 && ~x13 && ~x14 && ~x9 && ~x7 && x8 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s230;
						end
					else if( x62 && ~x13 && ~x14 && ~x9 && ~x7 && ~x8 )
						nx_state = s293;
					else if( ~x62 && x63 && x15 )
						nx_state = s1;
					else if( ~x62 && x63 && ~x15 && x13 && x4 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	
							nx_state = s231;
						end
					else if( ~x62 && x63 && ~x15 && x13 && ~x4 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( ~x62 && x63 && ~x15 && ~x13 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s230;
						end
					else if( ~x62 && x63 && ~x15 && ~x13 && ~x14 && x9 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s230;
						end
					else if( ~x62 && x63 && ~x15 && ~x13 && ~x14 && ~x9 && x7 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s230;
						end
					else if( ~x62 && x63 && ~x15 && ~x13 && ~x14 && ~x9 && ~x7 && x8 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s230;
						end
					else if( ~x62 && x63 && ~x15 && ~x13 && ~x14 && ~x9 && ~x7 && ~x8 )
						nx_state = s293;
					else if( ~x62 && ~x63 && x65 && x66 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x62 && ~x63 && x65 && x66 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x62 && ~x63 && x65 && x66 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x65 && x66 && ~x14 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x65 && ~x66 )
						begin
							y4 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s1034;
						end
					else if( ~x62 && ~x63 && ~x65 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && ~x63 && ~x65 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && ~x63 && ~x65 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x65 && ~x9 )
						nx_state = s1;
					else nx_state = s293;
				s294 : if( x63 && x64 && x18 && x15 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x63 && x64 && x18 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x63 && x64 && x18 && ~x15 && x16 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x63 && x64 && x18 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s299;
						end
					else if( x63 && x64 && ~x18 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s295;
						end
					else if( x63 && ~x64 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( ~x63 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else nx_state = s294;
				s295 : if( x64 && x63 )
						begin
							y3 = 1'b1;	y22 = 1'b1;	y37 = 1'b1;	
							nx_state = s1035;
						end
					else if( x64 && ~x63 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s102;
						end
					else if( ~x64 && x63 )
						nx_state = s1;
					else if( ~x64 && ~x63 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else nx_state = s295;
				s296 : if( x70 && x63 )
						begin
							y3 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s1036;
						end
					else if( x70 && ~x63 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s1037;
						end
					else if( ~x70 && x65 && x21 && x67 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( ~x70 && x65 && x21 && x67 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( ~x70 && x65 && x21 && x67 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x70 && x65 && x21 && x67 && ~x8 )
						nx_state = s1;
					else if( ~x70 && x65 && x21 && ~x67 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && x65 && x21 && ~x67 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && x21 && ~x67 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x65 && x21 && ~x67 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && x21 && ~x67 && ~x18 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && x23 && x22 && x67 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && x23 && x22 && x67 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && x23 && x22 && x67 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && x23 && x22 && x67 && ~x8 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && x23 && x22 && ~x67 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( ~x70 && x65 && ~x21 && x23 && x22 && ~x67 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x70 && x65 && ~x21 && x23 && x22 && ~x67 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x70 && x65 && ~x21 && x23 && x22 && ~x67 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && x23 && x22 && ~x67 && ~x19 && ~x17 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && x23 && ~x22 && x67 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && x23 && ~x22 && x67 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && x23 && ~x22 && x67 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && x23 && ~x22 && x67 && ~x9 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && x23 && ~x22 && ~x67 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( ~x70 && x65 && ~x21 && x23 && ~x22 && ~x67 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( ~x70 && x65 && ~x21 && x23 && ~x22 && ~x67 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && x23 && ~x22 && ~x67 && ~x20 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && ~x23 && x67 && x8 && x22 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && x67 && x8 && x22 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && x67 && x8 && x22 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && ~x23 && x67 && x8 && ~x22 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && x67 && x8 && ~x22 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && x67 && x8 && ~x22 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && ~x23 && x67 && ~x8 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && ~x23 && ~x67 && x18 && x14 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && ~x67 && x18 && x14 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && ~x67 && x18 && ~x14 && x13 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && ~x67 && x18 && ~x14 && x13 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x70 && x65 && ~x21 && ~x23 && ~x67 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && ~x23 && ~x67 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && ~x65 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && ~x65 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x62 && ~x61 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x65 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && ~x65 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x65 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && ~x65 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x65 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x65 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else nx_state = s296;
				s297 : if( x65 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x65 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x21 && x23 && x22 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( x65 && ~x21 && x23 && x22 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x65 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( x65 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x21 && x23 && x22 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x21 && x23 && ~x22 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x65 && ~x21 && x23 && ~x22 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( x65 && ~x21 && x23 && ~x22 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x21 && x23 && ~x22 && ~x20 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x23 && x18 && x14 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x65 && ~x21 && ~x23 && x18 && x14 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x65 && ~x21 && ~x23 && x18 && ~x14 && x13 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x65 && ~x21 && ~x23 && x18 && ~x14 && x13 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( x65 && ~x21 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x65 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x65 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x62 && ~x61 )
						nx_state = s1;
					else if( ~x65 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x65 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x65 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x65 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x65 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else nx_state = s297;
				s298 : if( x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x62 && ~x61 )
						nx_state = s1;
					else if( ~x62 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else nx_state = s298;
				s299 : if( x62 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s298;
						end
					else if( ~x62 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else nx_state = s299;
				s300 : if( x24 && x26 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x24 && x26 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x24 && x26 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x24 && x26 && ~x18 )
						nx_state = s1;
					else if( x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x24 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x25 && x19 && ~x14 && ~x13 && x26 )
						nx_state = s300;
					else if( ~x24 && x25 && x19 && ~x14 && ~x13 && ~x26 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else nx_state = s300;
				s301 : if( x70 && x7 && x6 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x70 && x7 && ~x6 && x5 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x70 && x7 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x70 && ~x7 )
						nx_state = s1;
					else if( ~x70 && x65 && x21 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x70 && x65 && ~x21 && x22 && x8 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && x22 && x8 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && x22 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && x22 && ~x8 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && ~x22 && x23 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && ~x22 && x23 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && ~x22 && x23 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && ~x22 && x23 && ~x9 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && ~x22 && ~x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && ~x22 && ~x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x21 && ~x22 && ~x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x21 && ~x22 && ~x23 && ~x8 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x24 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s300;
						end
					else if( ~x70 && ~x65 && ~x24 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x70 && ~x65 && ~x24 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x70 && ~x65 && ~x24 && x19 && ~x14 && ~x13 )
						nx_state = s301;
					else if( ~x70 && ~x65 && ~x24 && ~x19 )
						nx_state = s1;
					else nx_state = s301;
				s302 : if( x69 && x24 && x26 )
						nx_state = s1;
					else if( x69 && x24 && ~x26 )
						begin
							y11 = 1'b1;	y16 = 1'b1;	y25 = 1'b1;	
							nx_state = s515;
						end
					else if( x69 && ~x24 && x25 && x15 && x10 && x11 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s300;
						end
					else if( x69 && ~x24 && x25 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s1038;
						end
					else if( x69 && ~x24 && x25 && x15 && x10 && ~x11 && ~x12 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s300;
						end
					else if( x69 && ~x24 && x25 && x15 && ~x10 && x12 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s1039;
						end
					else if( x69 && ~x24 && x25 && x15 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s124;
						end
					else if( x69 && ~x24 && x25 && ~x15 && x16 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( x69 && ~x24 && x25 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( x69 && ~x24 && ~x25 && x26 )
						begin
							y11 = 1'b1;	y16 = 1'b1;	y25 = 1'b1;	
							nx_state = s515;
						end
					else if( x69 && ~x24 && ~x25 && ~x26 && x18 && x15 && x12 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x24 && ~x25 && ~x26 && x18 && x15 && ~x12 && x11 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x24 && ~x25 && ~x26 && x18 && x15 && ~x12 && ~x11 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x69 && ~x24 && ~x25 && ~x26 && x18 && x15 && ~x12 && ~x11 && ~x10 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( x69 && ~x24 && ~x25 && ~x26 && x18 && ~x15 && x16 && x10 && x12 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s497;
						end
					else if( x69 && ~x24 && ~x25 && ~x26 && x18 && ~x15 && x16 && x10 && ~x12 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s899;
						end
					else if( x69 && ~x24 && ~x25 && ~x26 && x18 && ~x15 && x16 && ~x10 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s497;
						end
					else if( x69 && ~x24 && ~x25 && ~x26 && x18 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x69 && ~x24 && ~x25 && ~x26 && ~x18 )
						begin
							y11 = 1'b1;	y16 = 1'b1;	y25 = 1'b1;	
							nx_state = s515;
						end
					else if( ~x69 && x70 && x62 && x3 && x5 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( ~x69 && x70 && x62 && x3 && ~x5 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x69 && x70 && x62 && ~x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && x70 && ~x62 && x64 && x3 && x5 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && x70 && ~x62 && x64 && x3 && ~x5 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x69 && x70 && ~x62 && x64 && ~x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && x70 && ~x62 && ~x64 && x63 && x3 && x5 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && x70 && ~x62 && ~x64 && x63 && x3 && ~x5 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x69 && x70 && ~x62 && ~x64 && x63 && ~x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && x70 && ~x62 && ~x64 && ~x63 && x42 && x5 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && x70 && ~x62 && ~x64 && ~x63 && x42 && ~x5 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s631;
						end
					else if( ~x69 && x70 && ~x62 && ~x64 && ~x63 && ~x42 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else if( ~x69 && ~x70 && x8 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s216;
						end
					else if( ~x69 && ~x70 && x8 && ~x1 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s816;
						end
					else if( ~x69 && ~x70 && x8 && ~x1 && ~x4 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && ~x70 && ~x8 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s733;
						end
					else nx_state = s302;
				s303 : if( x24 && x26 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x24 && x26 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x24 && x26 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x24 && x26 && ~x18 )
						nx_state = s1;
					else if( x24 && ~x26 )
						nx_state = s1;
					else if( ~x24 && x25 && x26 && x18 )
						nx_state = s1;
					else if( ~x24 && x25 && x26 && ~x18 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x24 && x25 && ~x26 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x25 && ~x26 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x25 && ~x26 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x26 && ~x19 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 )
						nx_state = s1;
					else nx_state = s303;
				s304 : if( x24 && x26 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x24 && x26 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x24 && x26 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x24 && x26 && ~x18 )
						nx_state = s1;
					else if( x24 && ~x26 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x24 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x25 && x19 && ~x14 && ~x13 && x26 )
						nx_state = s304;
					else if( ~x24 && x25 && x19 && ~x14 && ~x13 && ~x26 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && x5 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x5 && x18 && x15 && x12 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x5 && x18 && x15 && ~x12 && x11 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x5 && x18 && x15 && ~x12 && ~x11 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x5 && x18 && x15 && ~x12 && ~x11 && ~x10 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x5 && x18 && ~x15 && x16 && x10 && x12 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s497;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x5 && x18 && ~x15 && x16 && x10 && ~x12 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s899;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x5 && x18 && ~x15 && x16 && ~x10 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s497;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x5 && x18 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x5 && ~x18 )
						begin
							y11 = 1'b1;	y16 = 1'b1;	y25 = 1'b1;	
							nx_state = s515;
						end
					else nx_state = s304;
				s305 : if( x24 && x26 && x11 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s300;
						end
					else if( x24 && x26 && ~x11 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x24 && x26 && ~x11 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x24 && x26 && ~x11 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x24 && x26 && ~x11 && ~x18 )
						nx_state = s1;
					else if( x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x24 && x26 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x26 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x26 && x25 && x19 && ~x14 && ~x13 )
						nx_state = s305;
					else if( ~x24 && x26 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x24 && x26 && ~x25 && x10 && x12 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x24 && x26 && ~x25 && x10 && x12 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x24 && x26 && ~x25 && x10 && x12 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && x26 && ~x25 && x10 && x12 && ~x18 )
						nx_state = s1;
					else if( ~x24 && x26 && ~x25 && x10 && ~x12 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s304;
						end
					else if( ~x24 && x26 && ~x25 && ~x10 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x24 && x26 && ~x25 && ~x10 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x24 && x26 && ~x25 && ~x10 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && x26 && ~x25 && ~x10 && ~x18 )
						nx_state = s1;
					else if( ~x24 && ~x26 && x10 && x12 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && ~x26 && x10 && x12 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && ~x26 && x10 && x12 && x25 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x26 && x10 && x12 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x24 && ~x26 && x10 && x12 && ~x25 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x24 && ~x26 && x10 && x12 && ~x25 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x24 && ~x26 && x10 && x12 && ~x25 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x26 && x10 && x12 && ~x25 && ~x17 )
						nx_state = s1;
					else if( ~x24 && ~x26 && x10 && ~x12 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x24 && ~x26 && ~x10 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && ~x26 && ~x10 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && ~x26 && ~x10 && x25 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x26 && ~x10 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x24 && ~x26 && ~x10 && ~x25 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x24 && ~x26 && ~x10 && ~x25 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x24 && ~x26 && ~x10 && ~x25 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x26 && ~x10 && ~x25 && ~x17 )
						nx_state = s1;
					else nx_state = s305;
				s306 : if( x24 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s497;
						end
					else if( ~x24 )
						begin
							y8 = 1'b1;	y17 = 1'b1;	y23 = 1'b1;	
							nx_state = s303;
						end
					else nx_state = s306;
				s307 : if( x66 && x42 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x66 && x42 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x66 && x42 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( x66 && x42 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y28 = 1'b1;	
							nx_state = s299;
						end
					else if( x66 && ~x42 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s1040;
						end
					else if( ~x66 && x24 )
						nx_state = s1;
					else if( ~x66 && ~x24 && x25 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x66 && ~x24 && ~x25 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else nx_state = s307;
				s308 : if( 1'b1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else nx_state = s308;
				s309 : if( x24 && x26 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x24 && x26 && ~x4 && x20 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x24 && x26 && ~x4 && ~x20 && x21 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x24 && x26 && ~x4 && ~x20 && ~x21 && x22 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x24 && x26 && ~x4 && ~x20 && ~x21 && ~x22 && x23 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x24 && x26 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && x16 && x11 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( x24 && x26 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && x16 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x24 && x26 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && x13 && x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x24 && x26 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && x13 && ~x11 && x12 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( x24 && x26 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && x13 && ~x11 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x24 && x26 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && ~x13 && x11 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x24 && x26 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && ~x13 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x24 && x26 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s35;
						end
					else if( x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x24 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x25 && x19 && ~x14 && ~x13 && x26 )
						nx_state = s309;
					else if( ~x24 && x25 && x19 && ~x14 && ~x13 && ~x26 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else nx_state = s309;
				s310 : if( x70 && x63 && x22 && x16 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x70 && x63 && x22 && x16 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x70 && x63 && x22 && x16 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x70 && x63 && x22 && x16 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x70 && x63 && x22 && x16 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x70 && x63 && x22 && ~x16 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y65 = 1'b1;	
							y66 = 1'b1;	
							nx_state = s1041;
						end
					else if( x70 && x63 && ~x22 && x16 && x23 )
						begin
							y3 = 1'b1;	y30 = 1'b1;	y31 = 1'b1;	
							nx_state = s741;
						end
					else if( x70 && x63 && ~x22 && x16 && ~x23 && x7 && x9 && x10 && x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y38 = 1'b1;	
							y46 = 1'b1;	
							nx_state = s741;
						end
					else if( x70 && x63 && ~x22 && x16 && ~x23 && x7 && x9 && x10 && ~x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y38 = 1'b1;	
							y40 = 1'b1;	y41 = 1'b1;	
							nx_state = s741;
						end
					else if( x70 && x63 && ~x22 && x16 && ~x23 && x7 && x9 && ~x10 && x8 )
						begin
							y47 = 1'b1;	
							nx_state = s287;
						end
					else if( x70 && x63 && ~x22 && x16 && ~x23 && x7 && x9 && ~x10 && ~x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y38 = 1'b1;	
							y39 = 1'b1;	y41 = 1'b1;	
							nx_state = s741;
						end
					else if( x70 && x63 && ~x22 && x16 && ~x23 && x7 && ~x9 && x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y42 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s1042;
						end
					else if( x70 && x63 && ~x22 && x16 && ~x23 && x7 && ~x9 && ~x8 )
						begin
							y5 = 1'b1;	y35 = 1'b1;	y36 = 1'b1;	
							y38 = 1'b1;	y41 = 1'b1;	
							nx_state = s741;
						end
					else if( x70 && x63 && ~x22 && x16 && ~x23 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s523;
						end
					else if( x70 && x63 && ~x22 && ~x16 && x23 )
						begin
							y3 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s521;
						end
					else if( x70 && x63 && ~x22 && ~x16 && ~x23 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s524;
						end
					else if( x70 && ~x63 && x67 )
						begin
							y7 = 1'b1;	
							nx_state = s747;
						end
					else if( x70 && ~x63 && ~x67 && x21 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x63 && ~x67 && x21 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x63 && ~x67 && x21 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x67 && x21 && ~x6 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x67 && ~x21 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y62 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s518;
						end
					else if( ~x70 && x67 && x24 && x26 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && x67 && x24 && ~x26 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( ~x70 && x67 && ~x24 && x25 && x26 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && x67 && ~x24 && x25 && ~x26 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x70 && x67 && ~x24 && ~x25 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x70 && ~x67 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && ~x67 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && ~x67 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x70 && ~x67 && ~x3 )
						nx_state = s1;
					else nx_state = s310;
				s311 : if( x70 && x32 && x33 )
						begin
							y3 = 1'b1;	y52 = 1'b1;	
							nx_state = s23;
						end
					else if( x70 && x32 && ~x33 && x14 && x15 && x13 )
						begin
							y6 = 1'b1;	y35 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s338;
						end
					else if( x70 && x32 && ~x33 && x14 && x15 && ~x13 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s352;
						end
					else if( x70 && x32 && ~x33 && x14 && ~x15 && x13 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s349;
						end
					else if( x70 && x32 && ~x33 && x14 && ~x15 && ~x13 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s354;
						end
					else if( x70 && x32 && ~x33 && ~x14 && x15 && x13 && x16 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s347;
						end
					else if( x70 && x32 && ~x33 && ~x14 && x15 && x13 && ~x16 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s348;
						end
					else if( x70 && x32 && ~x33 && ~x14 && x15 && ~x13 && x17 )
						nx_state = s1;
					else if( x70 && x32 && ~x33 && ~x14 && x15 && ~x13 && ~x17 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s353;
						end
					else if( x70 && x32 && ~x33 && ~x14 && ~x15 && x13 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s350;
						end
					else if( x70 && x32 && ~x33 && ~x14 && ~x15 && ~x13 && x18 )
						nx_state = s1;
					else if( x70 && x32 && ~x33 && ~x14 && ~x15 && ~x13 && ~x18 )
						nx_state = s311;
					else if( x70 && ~x32 && x13 && x33 && x15 && x14 && x5 )
						begin
							y6 = 1'b1;	y35 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s338;
						end
					else if( x70 && ~x32 && x13 && x33 && x15 && x14 && ~x5 && x7 )
						begin
							y6 = 1'b1;	y35 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s338;
						end
					else if( x70 && ~x32 && x13 && x33 && x15 && x14 && ~x5 && ~x7 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y27 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s339;
						end
					else if( x70 && ~x32 && x13 && x33 && x15 && ~x14 && x31 && x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s340;
						end
					else if( x70 && ~x32 && x13 && x33 && x15 && ~x14 && x31 && ~x5 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( x70 && ~x32 && x13 && x33 && x15 && ~x14 && ~x31 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x70 && ~x32 && x13 && x33 && x15 && ~x14 && ~x31 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x70 && ~x32 && x13 && x33 && x15 && ~x14 && ~x31 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x32 && x13 && x33 && x15 && ~x14 && ~x31 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x32 && x13 && x33 && ~x15 && x14 && x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s343;
						end
					else if( x70 && ~x32 && x13 && x33 && ~x15 && x14 && ~x5 )
						begin
							y53 = 1'b1;	
							nx_state = s344;
						end
					else if( x70 && ~x32 && x13 && x33 && ~x15 && ~x14 && x16 && x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s340;
						end
					else if( x70 && ~x32 && x13 && x33 && ~x15 && ~x14 && x16 && ~x5 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( x70 && ~x32 && x13 && x33 && ~x15 && ~x14 && ~x16 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x70 && ~x32 && x13 && x33 && ~x15 && ~x14 && ~x16 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x70 && ~x32 && x13 && x33 && ~x15 && ~x14 && ~x16 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x32 && x13 && x33 && ~x15 && ~x14 && ~x16 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x32 && x13 && ~x33 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y35 = 1'b1;	y40 = 1'b1;	
							nx_state = s351;
						end
					else if( x70 && ~x32 && ~x13 && x33 && x14 && x15 && x8 && x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s340;
						end
					else if( x70 && ~x32 && ~x13 && x33 && x14 && x15 && x8 && ~x5 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( x70 && ~x32 && ~x13 && x33 && x14 && x15 && ~x8 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x70 && ~x32 && ~x13 && x33 && x14 && x15 && ~x8 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x70 && ~x32 && ~x13 && x33 && x14 && x15 && ~x8 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x32 && ~x13 && x33 && x14 && x15 && ~x8 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x32 && ~x13 && x33 && x14 && ~x15 && x30 && x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s340;
						end
					else if( x70 && ~x32 && ~x13 && x33 && x14 && ~x15 && x30 && ~x5 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( x70 && ~x32 && ~x13 && x33 && x14 && ~x15 && ~x30 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x70 && ~x32 && ~x13 && x33 && x14 && ~x15 && ~x30 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x70 && ~x32 && ~x13 && x33 && x14 && ~x15 && ~x30 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x32 && ~x13 && x33 && x14 && ~x15 && ~x30 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x32 && ~x13 && x33 && ~x14 && x15 && x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s340;
						end
					else if( x70 && ~x32 && ~x13 && x33 && ~x14 && x15 && ~x5 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( x70 && ~x32 && ~x13 && x33 && ~x14 && ~x15 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s345;
						end
					else if( x70 && ~x32 && ~x13 && ~x33 && x4 && x6 )
						begin
							y6 = 1'b1;	y35 = 1'b1;	y40 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s355;
						end
					else if( x70 && ~x32 && ~x13 && ~x33 && x4 && ~x6 )
						begin
							y15 = 1'b1;	
							nx_state = s22;
						end
					else if( x70 && ~x32 && ~x13 && ~x33 && ~x4 )
						begin
							y15 = 1'b1;	
							nx_state = s356;
						end
					else if( ~x70 && x67 )
						begin
							y15 = 1'b1;	
							nx_state = s243;
						end
					else if( ~x70 && ~x67 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s171;
						end
					else nx_state = s311;
				s312 : if( x70 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x70 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x70 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x24 && x26 )
						begin
							y11 = 1'b1;	y16 = 1'b1;	y25 = 1'b1;	
							nx_state = s515;
						end
					else if( ~x70 && x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x70 && x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x70 && ~x24 && x25 )
						nx_state = s1;
					else if( ~x70 && ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x70 && ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x70 && ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x24 && ~x25 && ~x26 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else nx_state = s312;
				s313 : if( x21 && x9 && x3 )
						nx_state = s47;
					else if( x21 && x9 && ~x3 && x4 )
						nx_state = s47;
					else if( x21 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( x21 && ~x9 )
						nx_state = s1;
					else if( ~x21 && x22 && x10 && x19 && x15 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y17 = 1'b1;	
							nx_state = s314;
						end
					else if( ~x21 && x22 && x10 && x19 && ~x15 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							nx_state = s315;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && x15 && x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s316;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && x15 && ~x14 && x16 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s316;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && x15 && ~x14 && ~x16 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && x15 && ~x14 && ~x16 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && x15 && ~x14 && ~x16 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && x10 && ~x19 && x20 && x15 && ~x14 && ~x16 && ~x5 )
						nx_state = s1;
					else if( ~x21 && x22 && x10 && ~x19 && x20 && ~x15 && x14 && x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s316;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && ~x15 && x14 && ~x18 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && ~x15 && x14 && ~x18 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && ~x15 && x14 && ~x18 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && x10 && ~x19 && x20 && ~x15 && x14 && ~x18 && ~x5 )
						nx_state = s1;
					else if( ~x21 && x22 && x10 && ~x19 && x20 && ~x15 && ~x14 && x17 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s316;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && x10 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && ~x5 )
						nx_state = s1;
					else if( ~x21 && x22 && x10 && ~x19 && ~x20 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( ~x21 && x22 && ~x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x22 && x19 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && ~x22 && x19 && ~x15 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	
							nx_state = s315;
						end
					else if( ~x21 && ~x22 && ~x19 && x20 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( ~x21 && ~x22 && ~x19 && ~x20 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else nx_state = s313;
				s314 : if( x21 && x9 && x3 )
						nx_state = s47;
					else if( x21 && x9 && ~x3 && x4 )
						nx_state = s47;
					else if( x21 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( x21 && ~x9 )
						nx_state = s1;
					else if( ~x21 && x22 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x5 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x19 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && ~x22 && x19 && ~x15 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	
							nx_state = s315;
						end
					else if( ~x21 && ~x22 && ~x19 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else nx_state = s314;
				s315 : if( x21 && x9 && x3 )
						nx_state = s47;
					else if( x21 && x9 && ~x3 && x4 )
						nx_state = s47;
					else if( x21 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( x21 && ~x9 )
						nx_state = s1;
					else if( ~x21 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x5 && ~x4 && x22 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x5 && ~x4 && x22 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x5 && ~x4 && ~x22 )
						nx_state = s1;
					else if( ~x21 && ~x5 && x22 )
						nx_state = s1;
					else if( ~x21 && ~x5 && ~x22 && x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && ~x5 && ~x22 && x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x5 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s315;
				s316 : if( x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x5 )
						nx_state = s1;
					else nx_state = s316;
				s317 : if( x70 && x62 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x70 && x62 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x70 && x62 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( x70 && x62 && ~x27 )
						nx_state = s1;
					else if( x70 && ~x62 && x63 && x65 && x4 && x5 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x62 && x63 && x65 && x4 && ~x5 )
						begin
							y69 = 1'b1;	y73 = 1'b1;	
							nx_state = s1043;
						end
					else if( x70 && ~x62 && x63 && x65 && ~x4 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( x70 && ~x62 && x63 && ~x65 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x62 && x63 && ~x65 && ~x13 )
						begin
							y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s572;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x65 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x65 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x65 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && x65 && ~x14 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x66 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x66 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x66 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && x66 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && ~x66 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && ~x66 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && ~x66 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x65 && ~x66 && ~x18 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && x66 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x66 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x66 && x20 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x66 && x20 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x66 && ~x20 )
						nx_state = s1;
					else if( ~x70 && x66 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && x66 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && x66 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && x66 && x62 && ~x61 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x66 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && x66 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x66 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && x66 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && x66 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && x66 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && x66 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && x66 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else if( ~x70 && ~x66 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s315;
						end
					else nx_state = s317;
				s318 : if( x69 && x21 && x6 )
						begin
							y8 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s172;
						end
					else if( x69 && x21 && ~x6 && x8 && x19 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && x21 && ~x6 && x8 && ~x19 && x20 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s313;
						end
					else if( x69 && x21 && ~x6 && x8 && ~x19 && ~x20 )
						begin
							y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s386;
						end
					else if( x69 && x21 && ~x6 && ~x8 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	
							nx_state = s895;
						end
					else if( x69 && ~x21 && x22 )
						nx_state = s1;
					else if( x69 && ~x21 && ~x22 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x69 && ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x69 && ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else if( ~x69 && x26 && x28 && x9 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( ~x69 && x26 && x28 && ~x9 && x23 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s941;
						end
					else if( ~x69 && x26 && x28 && ~x9 && ~x23 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( ~x69 && x26 && ~x28 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s942;
						end
					else if( ~x69 && ~x26 && x27 && x4 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s942;
						end
					else if( ~x69 && ~x26 && x27 && ~x4 )
						nx_state = s1;
					else if( ~x69 && ~x26 && ~x27 && x28 && x2 && x24 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s612;
						end
					else if( ~x69 && ~x26 && ~x27 && x28 && x2 && ~x24 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s614;
						end
					else if( ~x69 && ~x26 && ~x27 && x28 && ~x2 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s942;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && x18 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s613;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && x18 && ~x3 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && x18 && ~x3 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s614;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && ~x18 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s942;
						end
					else nx_state = s318;
				s319 : if( x64 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s1044;
						end
					else if( ~x64 && x3 && x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s19;
						end
					else if( ~x64 && x3 && ~x6 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x64 && ~x3 && x4 && x5 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x64 && ~x3 && x4 && x5 && ~x1 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( ~x64 && ~x3 && x4 && ~x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x64 && ~x3 && ~x4 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else nx_state = s319;
				s320 : if( x69 && x17 && x18 && x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	
							nx_state = s20;
						end
					else if( x69 && x17 && x18 && ~x1 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x69 && x17 && x18 && ~x1 && ~x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x17 && ~x18 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s320;
						end
					else if( x69 && x17 && ~x18 && ~x2 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( x69 && ~x17 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	
							nx_state = s20;
						end
					else if( ~x69 && x70 && x61 && x2 && x8 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && x70 && x61 && x2 && x8 && ~x1 && x35 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s840;
						end
					else if( ~x69 && x70 && x61 && x2 && x8 && ~x1 && ~x35 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( ~x69 && x70 && x61 && x2 && ~x8 && x32 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s874;
						end
					else if( ~x69 && x70 && x61 && x2 && ~x8 && x32 && ~x1 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x69 && x70 && x61 && x2 && ~x8 && x32 && ~x1 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s875;
						end
					else if( ~x69 && x70 && x61 && x2 && ~x8 && ~x32 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( ~x69 && x70 && x61 && ~x2 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( ~x69 && x70 && ~x61 && x37 && x28 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x69 && x70 && ~x61 && x37 && ~x28 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( ~x69 && x70 && ~x61 && ~x37 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s733;
						end
					else if( ~x69 && ~x70 && x44 && x2 && x10 && x1 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( ~x69 && ~x70 && x44 && x2 && x10 && x1 && ~x3 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x69 && ~x70 && x44 && x2 && x10 && x1 && ~x3 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x69 && ~x70 && x44 && x2 && x10 && ~x1 && x9 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x69 && ~x70 && x44 && x2 && x10 && ~x1 && ~x9 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x69 && ~x70 && x44 && x2 && ~x10 )
						nx_state = s320;
					else if( ~x69 && ~x70 && x44 && ~x2 && x10 && x1 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && ~x70 && x44 && ~x2 && x10 && ~x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x69 && ~x70 && x44 && ~x2 && ~x10 )
						nx_state = s320;
					else if( ~x69 && ~x70 && ~x44 && x10 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 && ~x1 && x3 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 && ~x1 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else nx_state = s320;
				s321 : if( x62 && x61 && x53 && x47 )
						nx_state = s321;
					else if( x62 && x61 && x53 && ~x47 && x59 && x51 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x62 && x61 && x53 && ~x47 && x59 && ~x51 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( x62 && x61 && x53 && ~x47 && ~x59 && x34 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( x62 && x61 && x53 && ~x47 && ~x59 && ~x34 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x62 && x61 && ~x53 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x62 && ~x61 && x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x62 && ~x61 && ~x11 && x1 && x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x62 && ~x61 && ~x11 && x1 && ~x2 && x3 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( x62 && ~x61 && ~x11 && x1 && ~x2 && ~x3 )
						nx_state = s321;
					else if( x62 && ~x61 && ~x11 && ~x1 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x62 && x63 && x55 && x53 && x47 )
						nx_state = s321;
					else if( ~x62 && x63 && x55 && x53 && ~x47 && x59 && x51 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s503;
						end
					else if( ~x62 && x63 && x55 && x53 && ~x47 && x59 && ~x51 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( ~x62 && x63 && x55 && x53 && ~x47 && ~x59 && x34 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( ~x62 && x63 && x55 && x53 && ~x47 && ~x59 && ~x34 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s503;
						end
					else if( ~x62 && x63 && x55 && ~x53 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s503;
						end
					else if( ~x62 && x63 && ~x55 && x11 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s503;
						end
					else if( ~x62 && x63 && ~x55 && ~x11 && x1 && x33 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s503;
						end
					else if( ~x62 && x63 && ~x55 && ~x11 && x1 && ~x33 && x34 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( ~x62 && x63 && ~x55 && ~x11 && x1 && ~x33 && ~x34 )
						nx_state = s321;
					else if( ~x62 && x63 && ~x55 && ~x11 && ~x1 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x62 && ~x63 && x40 && x48 && x42 && x51 && x47 )
						nx_state = s321;
					else if( ~x62 && ~x63 && x40 && x48 && x42 && x51 && ~x47 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x62 && ~x63 && x40 && x48 && x42 && ~x51 && x47 )
						nx_state = s321;
					else if( ~x62 && ~x63 && x40 && x48 && x42 && ~x51 && ~x47 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x62 && ~x63 && x40 && x48 && ~x42 && x47 )
						nx_state = s321;
					else if( ~x62 && ~x63 && x40 && x48 && ~x42 && ~x47 && x34 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x62 && ~x63 && x40 && x48 && ~x42 && ~x47 && ~x34 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x62 && ~x63 && x40 && ~x48 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x62 && ~x63 && ~x40 && x11 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x62 && ~x63 && ~x40 && ~x11 && x1 && x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x62 && ~x63 && ~x40 && ~x11 && x1 && ~x2 && x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x62 && ~x63 && ~x40 && ~x11 && x1 && ~x2 && ~x3 )
						nx_state = s321;
					else if( ~x62 && ~x63 && ~x40 && ~x11 && ~x1 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else nx_state = s321;
				s322 : if( x46 && x16 && x36 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s929;
						end
					else if( x46 && x16 && ~x36 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s932;
						end
					else if( x46 && ~x16 && x43 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s932;
						end
					else if( x46 && ~x16 && ~x43 )
						nx_state = s322;
					else if( ~x46 && x47 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s453;
						end
					else if( ~x46 && ~x47 && x44 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s441;
						end
					else if( ~x46 && ~x47 && ~x44 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s932;
						end
					else nx_state = s322;
				s323 : if( x15 && x16 && x5 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s440;
						end
					else if( x15 && x16 && ~x5 && x37 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x15 && x16 && ~x5 && ~x37 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s440;
						end
					else if( x15 && ~x16 && x37 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x15 && ~x16 && ~x37 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s442;
						end
					else if( ~x15 && x47 && x35 && x36 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x15 && x47 && x35 && ~x36 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x15 && x47 && ~x35 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s932;
						end
					else if( ~x15 && ~x47 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s440;
						end
					else nx_state = s323;
				s324 : if( x69 && x21 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( x69 && ~x21 && x16 && x10 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( x69 && ~x21 && x16 && ~x10 )
						begin
							y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s233;
						end
					else if( x69 && ~x21 && ~x16 && x17 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x21 && ~x16 && ~x17 )
						begin
							y5 = 1'b1;	y17 = 1'b1;	
							nx_state = s721;
						end
					else if( ~x69 && x15 && x16 && x63 && x36 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x15 && x16 && x63 && ~x36 )
						begin
							y21 = 1'b1;	y27 = 1'b1;	
							nx_state = s930;
						end
					else if( ~x69 && x15 && x16 && ~x63 && x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x15 && x16 && ~x63 && ~x5 )
						begin
							y21 = 1'b1;	y27 = 1'b1;	
							nx_state = s930;
						end
					else if( ~x69 && x15 && ~x16 && x13 && x11 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x15 && ~x16 && x13 && ~x11 && x63 && x37 && x4 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x69 && x15 && ~x16 && x13 && ~x11 && x63 && x37 && ~x4 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x69 && x15 && ~x16 && x13 && ~x11 && x63 && x37 && ~x4 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x15 && ~x16 && x13 && ~x11 && x63 && ~x37 && x36 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s440;
						end
					else if( ~x69 && x15 && ~x16 && x13 && ~x11 && x63 && ~x37 && ~x36 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( ~x69 && x15 && ~x16 && x13 && ~x11 && ~x63 && x6 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x69 && x15 && ~x16 && x13 && ~x11 && ~x63 && x6 && ~x4 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x69 && x15 && ~x16 && x13 && ~x11 && ~x63 && x6 && ~x4 && ~x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x15 && ~x16 && x13 && ~x11 && ~x63 && ~x6 && x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s445;
						end
					else if( ~x69 && x15 && ~x16 && x13 && ~x11 && ~x63 && ~x6 && ~x5 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( ~x69 && x15 && ~x16 && ~x13 && x63 && x45 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x15 && ~x16 && ~x13 && x63 && ~x45 && x40 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x15 && ~x16 && ~x13 && x63 && ~x45 && ~x40 && x6 && x2 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x15 && ~x16 && ~x13 && x63 && ~x45 && ~x40 && x6 && ~x2 )
						nx_state = s324;
					else if( ~x69 && x15 && ~x16 && ~x13 && x63 && ~x45 && ~x40 && ~x6 && x8 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x15 && ~x16 && ~x13 && x63 && ~x45 && ~x40 && ~x6 && ~x8 )
						nx_state = s324;
					else if( ~x69 && x15 && ~x16 && ~x13 && ~x63 && x14 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x15 && ~x16 && ~x13 && ~x63 && ~x14 && x9 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x15 && ~x16 && ~x13 && ~x63 && ~x14 && ~x9 && x6 && x2 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x15 && ~x16 && ~x13 && ~x63 && ~x14 && ~x9 && x6 && ~x2 )
						nx_state = s324;
					else if( ~x69 && x15 && ~x16 && ~x13 && ~x63 && ~x14 && ~x9 && ~x6 && x8 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x15 && ~x16 && ~x13 && ~x63 && ~x14 && ~x9 && ~x6 && ~x8 )
						nx_state = s324;
					else if( ~x69 && ~x15 && x63 && x47 && x35 && x5 && x33 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x69 && ~x15 && x63 && x47 && x35 && x5 && ~x33 && x1 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s453;
						end
					else if( ~x69 && ~x15 && x63 && x47 && x35 && x5 && ~x33 && ~x1 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s440;
						end
					else if( ~x69 && ~x15 && x63 && x47 && x35 && ~x5 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x69 && ~x15 && x63 && x47 && ~x35 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x69 && ~x15 && x63 && ~x47 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x69 && ~x15 && ~x63 && x16 && x4 && x5 && x2 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x69 && ~x15 && ~x63 && x16 && x4 && x5 && ~x2 && x1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s455;
						end
					else if( ~x69 && ~x15 && ~x63 && x16 && x4 && x5 && ~x2 && ~x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s445;
						end
					else if( ~x69 && ~x15 && ~x63 && x16 && x4 && ~x5 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x69 && ~x15 && ~x63 && x16 && ~x4 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x69 && ~x15 && ~x63 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else nx_state = s324;
				s325 : if( x63 && x46 && x47 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s442;
						end
					else if( x63 && x46 && ~x47 && x34 && x2 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s322;
						end
					else if( x63 && x46 && ~x47 && x34 && ~x2 )
						nx_state = s325;
					else if( x63 && x46 && ~x47 && ~x34 && x4 && x2 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( x63 && x46 && ~x47 && ~x34 && x4 && ~x2 )
						nx_state = s325;
					else if( x63 && x46 && ~x47 && ~x34 && ~x4 && x32 && x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x63 && x46 && ~x47 && ~x34 && ~x4 && x32 && ~x2 )
						nx_state = s325;
					else if( x63 && x46 && ~x47 && ~x34 && ~x4 && ~x32 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x63 && x46 && ~x47 && ~x34 && ~x4 && ~x32 && ~x2 )
						nx_state = s325;
					else if( x63 && ~x46 && x16 && x4 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s442;
						end
					else if( x63 && ~x46 && x16 && x4 && ~x5 && x1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s442;
						end
					else if( x63 && ~x46 && x16 && x4 && ~x5 && ~x1 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( x63 && ~x46 && x16 && ~x4 && x32 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s442;
						end
					else if( x63 && ~x46 && x16 && ~x4 && ~x32 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s453;
						end
					else if( x63 && ~x46 && ~x16 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s442;
						end
					else if( ~x63 && x16 && x15 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s446;
						end
					else if( ~x63 && x16 && ~x15 && x4 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s446;
						end
					else if( ~x63 && x16 && ~x15 && x4 && ~x5 && x64 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s446;
						end
					else if( ~x63 && x16 && ~x15 && x4 && ~x5 && x64 && ~x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x63 && x16 && ~x15 && x4 && ~x5 && ~x64 && x36 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s446;
						end
					else if( ~x63 && x16 && ~x15 && x4 && ~x5 && ~x64 && ~x36 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x63 && x16 && ~x15 && ~x4 && x64 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s446;
						end
					else if( ~x63 && x16 && ~x15 && ~x4 && x64 && ~x1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s455;
						end
					else if( ~x63 && x16 && ~x15 && ~x4 && ~x64 && x37 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s446;
						end
					else if( ~x63 && x16 && ~x15 && ~x4 && ~x64 && ~x37 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s455;
						end
					else if( ~x63 && ~x16 && x15 && x2 && x64 && x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s326;
						end
					else if( ~x63 && ~x16 && x15 && x2 && x64 && ~x3 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x63 && ~x16 && x15 && x2 && x64 && ~x3 && ~x4 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x63 && ~x16 && x15 && x2 && x64 && ~x3 && ~x4 && ~x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x63 && ~x16 && x15 && x2 && ~x64 && x31 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s326;
						end
					else if( ~x63 && ~x16 && x15 && x2 && ~x64 && ~x31 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x63 && ~x16 && x15 && x2 && ~x64 && ~x31 && ~x4 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x63 && ~x16 && x15 && x2 && ~x64 && ~x31 && ~x4 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x63 && ~x16 && x15 && ~x2 )
						nx_state = s325;
					else if( ~x63 && ~x16 && ~x15 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s446;
						end
					else nx_state = s325;
				s326 : if( x15 && x16 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s929;
						end
					else if( x15 && x16 && ~x5 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s932;
						end
					else if( x15 && ~x16 && x12 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s932;
						end
					else if( x15 && ~x16 && ~x12 )
						nx_state = s326;
					else if( ~x15 && x16 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s455;
						end
					else if( ~x15 && ~x16 && x13 && x64 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s441;
						end
					else if( ~x15 && ~x16 && x13 && ~x64 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s1045;
						end
					else if( ~x15 && ~x16 && ~x13 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s932;
						end
					else nx_state = s326;
				s327 : if( x64 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x64 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x64 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x64 && ~x9 )
						nx_state = s1;
					else if( ~x64 )
						begin
							y9 = 1'b1;	
							nx_state = s83;
						end
					else nx_state = s327;
				s328 : if( x64 && x63 && x4 && x5 && x3 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x64 && x63 && x4 && x5 && ~x3 && x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s651;
						end
					else if( x64 && x63 && x4 && x5 && ~x3 && ~x6 && x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s651;
						end
					else if( x64 && x63 && x4 && x5 && ~x3 && ~x6 && ~x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s652;
						end
					else if( x64 && x63 && x4 && ~x5 && x3 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( x64 && x63 && x4 && ~x5 && ~x3 && x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s653;
						end
					else if( x64 && x63 && x4 && ~x5 && ~x3 && ~x6 && x7 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s653;
						end
					else if( x64 && x63 && x4 && ~x5 && ~x3 && ~x6 && ~x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s654;
						end
					else if( x64 && x63 && ~x4 && x5 && x3 )
						begin
							y51 = 1'b1;	
							nx_state = s655;
						end
					else if( x64 && x63 && ~x4 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s654;
						end
					else if( x64 && x63 && ~x4 && ~x5 && x3 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y48 = 1'b1;	
							y50 = 1'b1;	
							nx_state = s654;
						end
					else if( x64 && x63 && ~x4 && ~x5 && ~x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s654;
						end
					else if( x64 && ~x63 && x66 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s1046;
						end
					else if( x64 && ~x63 && ~x66 && x67 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s938;
						end
					else if( x64 && ~x63 && ~x66 && ~x67 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s1047;
						end
					else if( ~x64 && x63 && x66 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s1048;
						end
					else if( ~x64 && x63 && ~x66 && x67 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s1048;
						end
					else if( ~x64 && x63 && ~x66 && ~x67 )
						begin
							y6 = 1'b1;	
							nx_state = s1049;
						end
					else if( ~x64 && ~x63 && x65 && x67 )
						begin
							y5 = 1'b1;	y42 = 1'b1;	y43 = 1'b1;	
							y68 = 1'b1;	
							nx_state = s1050;
						end
					else if( ~x64 && ~x63 && x65 && ~x67 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s1051;
						end
					else if( ~x64 && ~x63 && ~x65 && x66 && x67 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s1052;
						end
					else if( ~x64 && ~x63 && ~x65 && x66 && ~x67 )
						begin
							y6 = 1'b1;	
							nx_state = s1049;
						end
					else if( ~x64 && ~x63 && ~x65 && ~x66 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s1051;
						end
					else nx_state = s328;
				s329 : if( x69 )
						nx_state = s1;
					else if( ~x69 && x3 )
						nx_state = s1;
					else if( ~x69 && ~x3 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s209;
						end
					else nx_state = s329;
				s330 : if( x61 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( ~x61 && x15 && x12 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s491;
						end
					else if( ~x61 && x15 && x12 && ~x7 )
						begin
							y12 = 1'b1;	
							nx_state = s490;
						end
					else if( ~x61 && x15 && ~x12 && x7 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x61 && x15 && ~x12 && ~x7 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s566;
						end
					else if( ~x61 && ~x15 && x16 && x7 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s490;
						end
					else if( ~x61 && ~x15 && x16 && x7 && ~x12 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s565;
						end
					else if( ~x61 && ~x15 && x16 && ~x7 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s487;
						end
					else if( ~x61 && ~x15 && ~x16 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x61 && ~x15 && ~x16 && ~x7 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else nx_state = s330;
				s331 : if( x60 )
						nx_state = s1;
					else if( ~x60 && x61 )
						nx_state = s1;
					else if( ~x60 && ~x61 && x62 )
						begin
							y2 = 1'b1;	y19 = 1'b1;	y24 = 1'b1;	
							nx_state = s837;
						end
					else if( ~x60 && ~x61 && ~x62 )
						nx_state = s47;
					else nx_state = s331;
				s332 : if( x70 && x63 && x66 && x16 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && x63 && x66 && x16 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && x63 && x66 && x16 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x70 && x63 && x66 && ~x16 )
						nx_state = s1;
					else if( x70 && x63 && ~x66 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && x65 && x66 && x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x70 && ~x63 && x64 && x65 && x66 && x10 && ~x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x70 && ~x63 && x64 && x65 && x66 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && x65 && x66 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && x65 && ~x66 && x6 && x7 && x67 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x70 && ~x63 && x64 && x65 && ~x66 && x6 && x7 && ~x67 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x63 && x64 && x65 && ~x66 && x6 && ~x7 && x8 && x67 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x70 && ~x63 && x64 && x65 && ~x66 && x6 && ~x7 && x8 && ~x67 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x63 && x64 && x65 && ~x66 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && x65 && ~x66 && ~x6 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && ~x65 && x67 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x70 && ~x63 && x64 && ~x65 && x67 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x70 && ~x63 && x64 && ~x65 && x67 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && ~x65 && x67 && x22 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && ~x65 && x67 && ~x22 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && ~x65 && ~x67 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x63 && x64 && ~x65 && ~x67 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x63 && x64 && ~x65 && ~x67 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && ~x65 && ~x67 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x31 && x30 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x70 && ~x63 && ~x64 && x31 && ~x30 )
						begin
							y31 = 1'b1;	
							nx_state = s1053;
						end
					else if( x70 && ~x63 && ~x64 && ~x31 && x30 )
						begin
							y47 = 1'b1;	y49 = 1'b1;	y58 = 1'b1;	
							y61 = 1'b1;	y68 = 1'b1;	
							nx_state = s857;
						end
					else if( x70 && ~x63 && ~x64 && ~x31 && ~x30 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x70 && x21 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x70 && ~x21 && x23 && x22 && x5 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x70 && ~x21 && x23 && x22 && ~x5 && x18 && x15 && x9 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x21 && x23 && x22 && ~x5 && x18 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && ~x21 && x23 && x22 && ~x5 && x18 && ~x15 && x16 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x70 && ~x21 && x23 && x22 && ~x5 && x18 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s495;
						end
					else if( ~x70 && ~x21 && x23 && x22 && ~x5 && ~x18 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							nx_state = s165;
						end
					else if( ~x70 && ~x21 && x23 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x70 && ~x21 && ~x23 && x22 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x23 && ~x22 && x15 && x9 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && ~x21 && ~x23 && ~x22 && x15 && ~x9 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x70 && ~x21 && ~x23 && ~x22 && ~x15 && x16 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && ~x21 && ~x23 && ~x22 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s495;
						end
					else nx_state = s332;
				s333 : if( x21 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x21 && x22 && x23 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x21 && x22 && ~x23 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s406;
						end
					else if( ~x21 && ~x22 && x23 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s406;
						end
					else if( ~x21 && ~x22 && ~x23 && x18 && x14 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x21 && ~x22 && ~x23 && x18 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x21 && ~x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 && ~x18 )
						nx_state = s1;
					else nx_state = s333;
				s334 : if( x65 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x65 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else nx_state = s334;
				s335 : if( x70 )
						begin
							y14 = 1'b1;	
							nx_state = s124;
						end
					else if( ~x70 && x21 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x21 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && x21 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x9 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x22 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && ~x21 && ~x22 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else nx_state = s335;
				s336 : if( 1'b1 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else nx_state = s336;
				s337 : if( 1'b1 )
						begin
							y6 = 1'b1;	y47 = 1'b1;	
							nx_state = s1054;
						end
					else nx_state = s337;
				s338 : if( x32 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x32 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x32 && ~x10 )
						nx_state = s1;
					else if( ~x32 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s349;
						end
					else nx_state = s338;
				s339 : if( 1'b1 )
						begin
							y8 = 1'b1;	y31 = 1'b1;	
							nx_state = s1055;
						end
					else nx_state = s339;
				s340 : if( 1'b1 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s1056;
						end
					else nx_state = s340;
				s341 : if( x32 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x32 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x32 && ~x10 )
						nx_state = s1;
					else if( ~x32 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s974;
						end
					else nx_state = s341;
				s342 : if( x62 )
						nx_state = s1;
					else if( ~x62 && x63 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( ~x62 && x63 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( ~x62 && x63 && x19 && ~x14 && ~x13 && x11 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( ~x62 && x63 && x19 && ~x14 && ~x13 && x11 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x62 && x63 && x19 && ~x14 && ~x13 && ~x11 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x62 && x63 && ~x19 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && x65 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && ~x63 && x64 && x65 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && ~x63 && x64 && x65 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && x65 && ~x6 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && ~x65 && x66 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x62 && ~x63 && x64 && ~x65 && x66 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x62 && ~x63 && x64 && ~x65 && x66 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && ~x65 && x66 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && ~x65 && x66 && ~x22 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && ~x65 && ~x66 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x62 && ~x63 && x64 && ~x65 && ~x66 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x62 && ~x63 && x64 && ~x65 && ~x66 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && ~x65 && ~x66 && ~x18 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 )
						begin
							y5 = 1'b1;	y42 = 1'b1;	y43 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s1057;
						end
					else nx_state = s342;
				s343 : if( 1'b1 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s1058;
						end
					else nx_state = s343;
				s344 : if( x62 && x32 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x62 && x32 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x62 && x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x62 && x32 && ~x10 )
						nx_state = s1;
					else if( x62 && ~x32 && x33 )
						begin
							y8 = 1'b1;	y36 = 1'b1;	y42 = 1'b1;	
							nx_state = s969;
						end
					else if( x62 && ~x32 && ~x33 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x62 && ~x32 && ~x33 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x62 && ~x32 && ~x33 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x62 && ~x32 && ~x33 && ~x10 )
						nx_state = s1;
					else if( ~x62 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x62 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x62 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( ~x62 && ~x14 )
						nx_state = s1;
					else nx_state = s344;
				s345 : if( x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x10 )
						nx_state = s1;
					else nx_state = s345;
				s346 : if( x33 && x32 && x10 && x11 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s470;
						end
					else if( x33 && x32 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s470;
						end
					else if( x33 && x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x33 && x32 && ~x10 )
						nx_state = s1;
					else if( x33 && ~x32 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s311;
						end
					else if( ~x33 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s311;
						end
					else nx_state = s346;
				s347 : if( x32 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x32 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x32 && ~x10 )
						nx_state = s1;
					else if( ~x32 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s348;
						end
					else nx_state = s347;
				s348 : if( x32 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x32 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x32 && ~x10 )
						nx_state = s1;
					else if( ~x32 && x33 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y12 = 1'b1;	
							y37 = 1'b1;	y38 = 1'b1;	
							nx_state = s1059;
						end
					else if( ~x32 && ~x33 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y35 = 1'b1;	y40 = 1'b1;	
							nx_state = s351;
						end
					else nx_state = s348;
				s349 : if( x32 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x32 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x32 && ~x10 )
						nx_state = s1;
					else if( ~x32 && x33 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s347;
						end
					else if( ~x32 && ~x33 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x32 && ~x33 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x32 && ~x33 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x32 && ~x33 && ~x10 )
						nx_state = s1;
					else nx_state = s349;
				s350 : if( 1'b1 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s1060;
						end
					else nx_state = s350;
				s351 : if( x33 && x32 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s1061;
						end
					else if( x33 && ~x32 && x30 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s1061;
						end
					else if( x33 && ~x32 && ~x30 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x33 && ~x32 && ~x30 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x33 && ~x32 && ~x30 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x33 && ~x32 && ~x30 && ~x10 )
						nx_state = s1;
					else if( ~x33 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s1061;
						end
					else nx_state = s351;
				s352 : if( 1'b1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	y40 = 1'b1;	
							nx_state = s1062;
						end
					else nx_state = s352;
				s353 : if( 1'b1 )
						begin
							y30 = 1'b1;	
							nx_state = s416;
						end
					else nx_state = s353;
				s354 : if( 1'b1 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s1063;
						end
					else nx_state = s354;
				s355 : if( x32 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x32 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x32 && ~x10 )
						nx_state = s1;
					else if( ~x32 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s973;
						end
					else nx_state = s355;
				s356 : if( x62 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1064;
						end
					else if( ~x62 && x20 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y45 = 1'b1;	
							y49 = 1'b1;	
							nx_state = s1065;
						end
					else if( ~x62 && ~x20 && x21 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1066;
						end
					else if( ~x62 && ~x20 && ~x21 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else nx_state = s356;
				s357 : if( x21 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x21 && x22 && x15 && x10 && x16 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x21 && x22 && x15 && x10 && x16 && ~x12 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s363;
						end
					else if( ~x21 && x22 && x15 && x10 && ~x16 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x21 && x22 && x15 && x10 && ~x16 && ~x3 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && x22 && x15 && x10 && ~x16 && ~x3 && ~x2 && x11 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s358;
						end
					else if( ~x21 && x22 && x15 && x10 && ~x16 && ~x3 && ~x2 && ~x11 && x12 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s851;
						end
					else if( ~x21 && x22 && x15 && x10 && ~x16 && ~x3 && ~x2 && ~x11 && ~x12 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s274;
						end
					else if( ~x21 && x22 && x15 && ~x10 && x11 && x12 && x16 )
						begin
							y14 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x21 && x22 && x15 && ~x10 && x11 && x12 && ~x16 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x21 && x22 && x15 && ~x10 && x11 && x12 && ~x16 && ~x3 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && x22 && x15 && ~x10 && x11 && x12 && ~x16 && ~x3 && ~x2 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s367;
						end
					else if( ~x21 && x22 && x15 && ~x10 && x11 && ~x12 && x16 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && x15 && ~x10 && x11 && ~x12 && ~x16 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s275;
						end
					else if( ~x21 && x22 && x15 && ~x10 && ~x11 && x16 && x12 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( ~x21 && x22 && x15 && ~x10 && ~x11 && x16 && x12 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x22 && x15 && ~x10 && ~x11 && x16 && ~x12 && x14 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( ~x21 && x22 && x15 && ~x10 && ~x11 && x16 && ~x12 && ~x14 )
						nx_state = s1;
					else if( ~x21 && x22 && x15 && ~x10 && ~x11 && ~x16 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x21 && x22 && x15 && ~x10 && ~x11 && ~x16 && ~x3 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && x22 && x15 && ~x10 && ~x11 && ~x16 && ~x3 && ~x2 && x12 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x21 && x22 && x15 && ~x10 && ~x11 && ~x16 && ~x3 && ~x2 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s124;
						end
					else if( ~x21 && x22 && ~x15 && x16 && x12 && x10 && x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x15 && x16 && x12 && x10 && ~x8 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x21 && x22 && ~x15 && x16 && x12 && x10 && ~x8 && ~x3 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && x22 && ~x15 && x16 && x12 && x10 && ~x8 && ~x3 && ~x2 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x21 && x22 && ~x15 && x16 && x12 && ~x10 && x11 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x21 && x22 && ~x15 && x16 && x12 && ~x10 && x11 && ~x3 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && x22 && ~x15 && x16 && x12 && ~x10 && x11 && ~x3 && ~x2 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x21 && x22 && ~x15 && x16 && x12 && ~x10 && ~x11 && x7 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x21 && x22 && ~x15 && x16 && x12 && ~x10 && ~x11 && x7 && ~x3 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x21 && x22 && ~x15 && x16 && x12 && ~x10 && ~x11 && x7 && ~x3 && ~x2 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x21 && x22 && ~x15 && x16 && x12 && ~x10 && ~x11 && ~x7 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && x10 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && x10 && ~x3 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s567;
						end
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && x10 && ~x3 && ~x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && ~x10 && x11 && x9 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && ~x10 && x11 && x9 && ~x3 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && ~x10 && x11 && x9 && ~x3 && ~x2 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && ~x10 && x11 && ~x9 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && ~x10 && ~x11 && x8 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && ~x10 && ~x11 && x8 && ~x3 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && ~x10 && ~x11 && x8 && ~x3 && ~x2 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && ~x10 && ~x11 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x15 && ~x16 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x21 && x22 && ~x15 && ~x16 && ~x3 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && x22 && ~x15 && ~x16 && ~x3 && ~x2 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x19 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else nx_state = s357;
				s358 : if( x70 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x70 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x70 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x65 && x67 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && x67 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && x67 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x65 && x67 && x22 && ~x17 )
						nx_state = s1;
					else if( ~x70 && x65 && x67 && ~x22 && x18 && x13 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && x65 && x67 && ~x22 && x18 && x13 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x65 && x67 && ~x22 && x18 && ~x13 && x12 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && x65 && x67 && ~x22 && x18 && ~x13 && x12 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x65 && x67 && ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && x65 && x67 && ~x22 && ~x18 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x67 && x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x67 && x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x65 && ~x67 && x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x67 && x21 && x20 && ~x17 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x67 && x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x65 && ~x67 && x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x65 && ~x67 && x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x67 && x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x67 && ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x65 && ~x67 && ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x65 && ~x67 && ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x67 && ~x21 && ~x19 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && x21 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s67;
						end
					else if( ~x70 && ~x65 && x66 && ~x21 && x23 && x22 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && ~x65 && x66 && ~x21 && x23 && ~x22 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x70 && ~x65 && x66 && ~x21 && x23 && ~x22 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x70 && ~x65 && x66 && ~x21 && x23 && ~x22 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && ~x21 && x23 && ~x22 && ~x19 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x66 && ~x21 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x65 && ~x66 && x67 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && ~x66 && x67 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x65 && ~x66 && x67 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && x67 && x20 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && x67 && ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x70 && ~x65 && ~x66 && x67 && ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x70 && ~x65 && ~x66 && x67 && ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && x67 && ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && x67 && ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x70 && ~x65 && ~x66 && x67 && ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x70 && ~x65 && ~x66 && x67 && ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && x67 && ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && ~x67 && x21 && x19 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && x21 && ~x19 && x20 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s313;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && x21 && ~x19 && ~x20 )
						begin
							y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s386;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && x13 && x20 && x15 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && x13 && x20 && ~x15 )
						begin
							y22 = 1'b1;	y25 = 1'b1;	
							nx_state = s315;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && x13 && ~x20 )
						begin
							y2 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s385;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && x20 && x14 && x15 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	y23 = 1'b1;	
							nx_state = s383;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && x20 && x14 && ~x15 )
						begin
							y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s386;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && x20 && ~x14 && x15 && x6 )
						begin
							y12 = 1'b1;	
							nx_state = s493;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && x20 && ~x14 && x15 && ~x6 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && x20 && ~x14 && x15 && ~x6 && x5 && ~x4 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && x20 && ~x14 && x15 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && x20 && ~x14 && ~x15 && x4 )
						begin
							y12 = 1'b1;	
							nx_state = s493;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && x20 && ~x14 && ~x15 && ~x4 && x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && x20 && ~x14 && ~x15 && ~x4 && x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && x20 && ~x14 && ~x15 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && ~x20 && x14 )
						begin
							y2 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s385;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && ~x20 && ~x14 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s850;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && ~x20 && ~x14 && ~x7 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s169;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && ~x20 && ~x14 && ~x7 && ~x8 && x15 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	
							nx_state = s895;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && ~x20 && ~x14 && ~x7 && ~x8 && ~x15 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	
							nx_state = s315;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && ~x19 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s850;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && ~x19 && ~x7 && x20 && x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && ~x19 && ~x7 && x20 && x15 && ~x14 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s169;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && ~x19 && ~x7 && x20 && ~x15 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s169;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && ~x19 && ~x7 && ~x20 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s169;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && x22 && ~x19 && ~x7 && ~x20 && ~x8 )
						begin
							y21 = 1'b1;	y24 = 1'b1;	
							nx_state = s684;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && ~x22 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x66 && ~x67 && ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s358;
				s359 : if( x21 && x65 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x21 && x65 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x21 && x65 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x65 && x20 && ~x17 )
						nx_state = s1;
					else if( x21 && x65 && ~x20 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( x21 && ~x65 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x21 && ~x65 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x21 && ~x65 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x65 && ~x18 )
						nx_state = s1;
					else if( ~x21 && x65 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && ~x65 && x22 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x21 && ~x65 && x22 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x21 && ~x65 && x22 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x65 && x22 && x23 && ~x17 )
						nx_state = s1;
					else if( ~x21 && ~x65 && x22 && ~x23 && x18 && x14 )
						nx_state = s47;
					else if( ~x21 && ~x65 && x22 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s47;
					else if( ~x21 && ~x65 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x65 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x21 && ~x65 && ~x22 && x23 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s362;
						end
					else if( ~x21 && ~x65 && ~x22 && ~x23 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s1067;
						end
					else nx_state = s359;
				s360 : if( 1'b1 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else nx_state = s360;
				s361 : if( x21 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x21 && x22 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x21 && x22 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x21 && x22 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x17 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s365;
						end
					else if( ~x21 && ~x22 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s362;
						end
					else nx_state = s361;
				s362 : if( x21 && x16 && x15 && x10 && x12 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x21 && x16 && x15 && x10 && ~x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x21 && x16 && x15 && ~x10 && x11 && x12 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s363;
						end
					else if( x21 && x16 && x15 && ~x10 && x11 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s5;
						end
					else if( x21 && x16 && x15 && ~x10 && ~x11 && x12 && x13 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s852;
						end
					else if( x21 && x16 && x15 && ~x10 && ~x11 && x12 && ~x13 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x21 && x16 && x15 && ~x10 && ~x11 && x12 && ~x13 && x18 && ~x14 )
						nx_state = s1;
					else if( x21 && x16 && x15 && ~x10 && ~x11 && x12 && ~x13 && ~x18 )
						nx_state = s1;
					else if( x21 && x16 && x15 && ~x10 && ~x11 && ~x12 && x14 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s852;
						end
					else if( x21 && x16 && x15 && ~x10 && ~x11 && ~x12 && ~x14 && x18 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x21 && x16 && x15 && ~x10 && ~x11 && ~x12 && ~x14 && x18 && ~x13 )
						nx_state = s1;
					else if( x21 && x16 && x15 && ~x10 && ~x11 && ~x12 && ~x14 && ~x18 )
						nx_state = s1;
					else if( x21 && x16 && ~x15 && x12 && x10 && x8 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x21 && x16 && ~x15 && x12 && x10 && x8 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x21 && x16 && ~x15 && x12 && x10 && x8 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x16 && ~x15 && x12 && x10 && x8 && ~x18 )
						nx_state = s1;
					else if( x21 && x16 && ~x15 && x12 && x10 && ~x8 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x21 && x16 && ~x15 && x12 && x10 && ~x8 && ~x3 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x21 && x16 && ~x15 && x12 && x10 && ~x8 && ~x3 && ~x5 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x21 && x16 && ~x15 && x12 && ~x10 && x7 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x21 && x16 && ~x15 && x12 && ~x10 && x7 && ~x3 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x21 && x16 && ~x15 && x12 && ~x10 && x7 && ~x3 && ~x5 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x21 && x16 && ~x15 && x12 && ~x10 && ~x7 && x11 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x21 && x16 && ~x15 && x12 && ~x10 && ~x7 && x11 && ~x3 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x21 && x16 && ~x15 && x12 && ~x10 && ~x7 && x11 && ~x3 && ~x5 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x21 && x16 && ~x15 && x12 && ~x10 && ~x7 && ~x11 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x21 && x16 && ~x15 && x12 && ~x10 && ~x7 && ~x11 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x21 && x16 && ~x15 && x12 && ~x10 && ~x7 && ~x11 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x16 && ~x15 && x12 && ~x10 && ~x7 && ~x11 && ~x18 )
						nx_state = s1;
					else if( x21 && x16 && ~x15 && ~x12 && x10 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x21 && x16 && ~x15 && ~x12 && x10 && ~x3 && x5 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s706;
						end
					else if( x21 && x16 && ~x15 && ~x12 && x10 && ~x3 && ~x5 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s361;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && x11 && x9 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && x11 && x9 && ~x3 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && x11 && x9 && ~x3 && ~x5 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && ~x18 )
						nx_state = s1;
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && ~x11 && x8 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && ~x11 && x8 && ~x3 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && ~x11 && x8 && ~x3 && ~x5 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && ~x18 )
						nx_state = s1;
					else if( x21 && ~x16 && x15 && x10 && x11 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x21 && ~x16 && x15 && x10 && ~x11 && x12 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s358;
						end
					else if( x21 && ~x16 && x15 && x10 && ~x11 && ~x12 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x21 && ~x16 && x15 && x10 && ~x11 && ~x12 && ~x3 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x21 && ~x16 && x15 && x10 && ~x11 && ~x12 && ~x3 && ~x5 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x21 && ~x16 && x15 && ~x10 && x11 && x12 )
						begin
							y14 = 1'b1;	
							nx_state = s366;
						end
					else if( x21 && ~x16 && x15 && ~x10 && x11 && ~x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x21 && ~x16 && x15 && ~x10 && ~x11 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x21 && ~x16 && x15 && ~x10 && ~x11 && ~x3 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x21 && ~x16 && x15 && ~x10 && ~x11 && ~x3 && ~x5 && x12 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s275;
						end
					else if( x21 && ~x16 && x15 && ~x10 && ~x11 && ~x3 && ~x5 && ~x12 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s851;
						end
					else if( x21 && ~x16 && ~x15 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x21 && ~x16 && ~x15 && ~x3 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x21 && ~x16 && ~x15 && ~x3 && ~x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s57;
						end
					else if( ~x21 && x22 && x23 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x21 && x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x19 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 && x18 && x14 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x21 && ~x22 && ~x23 && x18 && ~x14 && x13 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x21 && ~x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 && ~x18 )
						nx_state = s1;
					else nx_state = s362;
				s363 : if( x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x18 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x21 && x22 && x23 && ~x4 && x18 && x15 && x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x21 && x22 && x23 && ~x4 && x18 && x15 && ~x10 && x12 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x21 && x22 && x23 && ~x4 && x18 && x15 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s366;
						end
					else if( ~x21 && x22 && x23 && ~x4 && x18 && ~x15 && x16 && x10 && x12 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else if( ~x21 && x22 && x23 && ~x4 && x18 && ~x15 && x16 && x10 && ~x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x21 && x22 && x23 && ~x4 && x18 && ~x15 && x16 && ~x10 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else if( ~x21 && x22 && x23 && ~x4 && x18 && ~x15 && ~x16 )
						nx_state = s47;
					else if( ~x21 && x22 && x23 && ~x4 && ~x18 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && x22 && ~x23 && x18 && x14 )
						nx_state = s47;
					else if( ~x21 && x22 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s47;
					else if( ~x21 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x19 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else nx_state = s363;
				s364 : if( x65 && x66 && x22 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	
							nx_state = s486;
						end
					else if( x65 && x66 && ~x22 && x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x65 && x66 && ~x22 && ~x23 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x65 && ~x66 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && ~x66 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && ~x66 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x5 )
						nx_state = s1;
					else if( ~x65 && x66 && x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x65 && x66 && x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x65 && x66 && x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x66 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x21 && x22 && x23 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else if( ~x65 && x66 && ~x21 && x22 && ~x23 && x18 && x14 )
						nx_state = s47;
					else if( ~x65 && x66 && ~x21 && x22 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s47;
					else if( ~x65 && x66 && ~x21 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x21 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x21 && ~x22 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x21 && ~x22 && x23 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x21 && ~x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x65 && ~x66 && x20 && x15 && x16 && x8 && x14 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x65 && ~x66 && x20 && x15 && x16 && x8 && ~x14 && x7 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s358;
						end
					else if( ~x65 && ~x66 && x20 && x15 && x16 && x8 && ~x14 && ~x7 && x12 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( ~x65 && ~x66 && x20 && x15 && x16 && x8 && ~x14 && ~x7 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x20 && x15 && x16 && ~x8 && x14 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x65 && ~x66 && x20 && x15 && x16 && ~x8 && ~x14 && x7 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	y20 = 1'b1;	
							nx_state = s781;
						end
					else if( ~x65 && ~x66 && x20 && x15 && x16 && ~x8 && ~x14 && ~x7 && x13 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( ~x65 && ~x66 && x20 && x15 && x16 && ~x8 && ~x14 && ~x7 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x20 && x15 && ~x16 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( ~x65 && ~x66 && x20 && x15 && ~x16 && ~x7 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( ~x65 && ~x66 && x20 && x15 && ~x16 && ~x7 && ~x5 && x8 && x1 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x65 && ~x66 && x20 && x15 && ~x16 && ~x7 && ~x5 && x8 && ~x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x65 && ~x66 && x20 && x15 && ~x16 && ~x7 && ~x5 && ~x8 && x1 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x65 && ~x66 && x20 && x15 && ~x16 && ~x7 && ~x5 && ~x8 && ~x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && x7 && x8 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && x7 && x8 && ~x5 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && x7 && ~x8 && x11 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && x7 && ~x8 && x11 && ~x5 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && x7 && ~x8 && ~x11 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && x7 && ~x8 && ~x11 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && x7 && ~x8 && ~x11 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && x7 && ~x8 && ~x11 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && x8 && x9 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && x8 && x9 && ~x5 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && x8 && ~x9 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && x8 && ~x9 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && x8 && ~x9 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && x8 && ~x9 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && ~x8 && x10 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && ~x8 && x10 && ~x5 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && ~x8 && ~x10 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && ~x8 && ~x10 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && ~x8 && ~x10 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && ~x8 && ~x10 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x20 && ~x15 && ~x16 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && ~x16 && ~x5 && x1 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && ~x16 && ~x5 && ~x1 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else if( ~x65 && ~x66 && ~x20 )
						nx_state = s1;
					else nx_state = s364;
				s365 : if( x68 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x68 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x68 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( x68 && ~x7 )
						nx_state = s1;
					else if( ~x68 && x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x68 && x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x68 && x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x68 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x68 && ~x21 && x22 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x68 && ~x21 && x22 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x68 && ~x21 && x22 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x68 && ~x21 && x22 && x23 && ~x17 )
						nx_state = s1;
					else if( ~x68 && ~x21 && x22 && ~x23 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s605;
						end
					else if( ~x68 && ~x21 && ~x22 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x68 && ~x21 && ~x22 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x68 && ~x21 && ~x22 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x68 && ~x21 && ~x22 && x23 && ~x19 )
						nx_state = s1;
					else if( ~x68 && ~x21 && ~x22 && ~x23 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s362;
						end
					else nx_state = s365;
				s366 : if( x70 && x62 )
						begin
							y5 = 1'b1;	
							nx_state = s64;
						end
					else if( x70 && ~x62 && x63 )
						begin
							y6 = 1'b1;	y17 = 1'b1;	y34 = 1'b1;	
							nx_state = s1068;
						end
					else if( x70 && ~x62 && ~x63 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x70 && x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x22 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x70 && ~x21 && x22 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x70 && ~x21 && x22 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x22 && x23 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x22 && ~x23 && x18 && x14 )
						nx_state = s47;
					else if( ~x70 && ~x21 && x22 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s47;
					else if( ~x70 && ~x21 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s362;
						end
					else nx_state = s366;
				s367 : if( x68 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x68 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x68 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( x68 && ~x7 )
						nx_state = s1;
					else if( ~x68 && x21 )
						begin
							y5 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x68 && ~x21 && x22 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x68 && ~x21 && x22 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x68 && ~x21 && x22 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x68 && ~x21 && x22 && x23 && ~x17 )
						nx_state = s1;
					else if( ~x68 && ~x21 && x22 && ~x23 && x18 && x14 )
						nx_state = s47;
					else if( ~x68 && ~x21 && x22 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s47;
					else if( ~x68 && ~x21 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x68 && ~x21 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x68 && ~x21 && ~x22 && x23 )
						nx_state = s1;
					else if( ~x68 && ~x21 && ~x22 && ~x23 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s362;
						end
					else nx_state = s367;
				s368 : if( x70 && x62 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s536;
						end
					else if( x70 && ~x62 && x65 )
						begin
							y7 = 1'b1;	
							nx_state = s748;
						end
					else if( x70 && ~x62 && ~x65 )
						begin
							y12 = 1'b1;	y48 = 1'b1;	
							nx_state = s1069;
						end
					else if( ~x70 && x66 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x70 && ~x66 && x24 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else if( ~x70 && ~x66 && ~x24 && x26 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x66 && ~x24 && ~x26 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else nx_state = s368;
				s369 : if( x68 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	y22 = 1'b1;	
							nx_state = s1070;
						end
					else if( ~x68 && x26 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x68 && ~x26 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s122;
						end
					else nx_state = s369;
				s370 : if( x26 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s304;
						end
					else if( ~x26 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else nx_state = s370;
				s371 : if( x70 )
						begin
							y53 = 1'b1;	
							nx_state = s1071;
						end
					else if( ~x70 && x65 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( ~x70 && ~x65 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s35;
						end
					else nx_state = s371;
				s372 : if( 1'b1 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else nx_state = s372;
				s373 : if( x70 && x64 && x21 && x3 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else if( x70 && x64 && x21 && ~x3 )
						begin
							y31 = 1'b1;	
							nx_state = s1072;
						end
					else if( x70 && x64 && ~x21 && x3 )
						begin
							y14 = 1'b1;	
							nx_state = s366;
						end
					else if( x70 && x64 && ~x21 && ~x3 )
						begin
							y31 = 1'b1;	
							nx_state = s1073;
						end
					else if( x70 && ~x64 )
						begin
							y48 = 1'b1;	y57 = 1'b1;	y61 = 1'b1;	
							nx_state = s954;
						end
					else if( ~x70 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else nx_state = s373;
				s374 : if( 1'b1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else nx_state = s374;
				s375 : if( 1'b1 )
						begin
							y18 = 1'b1;	
							nx_state = s981;
						end
					else nx_state = s375;
				s376 : if( x70 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && x20 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && x20 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x20 )
						nx_state = s1;
					else if( ~x70 && x21 && x8 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s576;
						end
					else if( ~x70 && x21 && ~x8 && x19 && x18 && x17 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s574;
						end
					else if( ~x70 && x21 && ~x8 && x19 && x18 && x17 && ~x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s574;
						end
					else if( ~x70 && x21 && ~x8 && x19 && x18 && ~x17 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x21 && ~x8 && x19 && x18 && ~x17 && ~x12 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s377;
						end
					else if( ~x70 && x21 && ~x8 && x19 && ~x18 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s575;
						end
					else if( ~x70 && x21 && ~x8 && ~x19 && x9 && x20 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s574;
						end
					else if( ~x70 && x21 && ~x8 && ~x19 && x9 && x20 && ~x12 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s171;
						end
					else if( ~x70 && x21 && ~x8 && ~x19 && x9 && ~x20 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s573;
						end
					else if( ~x70 && x21 && ~x8 && ~x19 && x9 && ~x20 && ~x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x70 && x21 && ~x8 && ~x19 && ~x9 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s575;
						end
					else if( ~x70 && ~x21 && x22 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s168;
						end
					else nx_state = s376;
				s377 : if( x21 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x21 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x21 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x21 && ~x3 )
						nx_state = s1;
					else if( ~x21 && x22 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x21 && x22 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x21 && x22 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x21 && ~x22 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x21 && ~x22 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x8 )
						nx_state = s1;
					else nx_state = s377;
				s378 : if( x21 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( ~x21 && x22 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	
							nx_state = s594;
						end
					else if( ~x21 && ~x22 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else nx_state = s378;
				s379 : if( 1'b1 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else nx_state = s379;
				s380 : if( x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x6 )
						nx_state = s1;
					else nx_state = s380;
				s381 : if( 1'b1 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s382;
						end
					else nx_state = s381;
				s382 : if( 1'b1 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else nx_state = s382;
				s383 : if( x21 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s315;
						end
					else if( ~x21 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x5 && ~x4 && x22 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x5 && ~x4 && x22 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x5 && ~x4 && ~x22 )
						nx_state = s1;
					else if( ~x21 && ~x5 && x22 )
						nx_state = s1;
					else if( ~x21 && ~x5 && ~x22 && x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && ~x5 && ~x22 && x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x5 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s383;
				s384 : if( x65 && x60 && x61 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s117;
						end
					else if( x65 && x60 && ~x61 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s139;
						end
					else if( x65 && ~x60 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s139;
						end
					else if( ~x65 && x68 && x19 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s894;
						end
					else if( ~x65 && x68 && ~x19 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && ~x68 && x21 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && ~x68 && ~x21 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	
							nx_state = s895;
						end
					else nx_state = s384;
				s385 : if( x22 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s315;
						end
					else if( ~x22 && x21 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s315;
						end
					else if( ~x22 && ~x21 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x22 && ~x21 && x4 && ~x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x22 && ~x21 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x22 && ~x21 && ~x4 )
						nx_state = s1;
					else nx_state = s385;
				s386 : if( x22 && x21 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s315;
						end
					else if( x22 && ~x21 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x22 && ~x21 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x22 && ~x21 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( x22 && ~x21 && ~x5 )
						nx_state = s1;
					else if( ~x22 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s315;
						end
					else nx_state = s386;
				s387 : if( x44 && x28 && x18 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( x44 && x28 && ~x18 )
						nx_state = s387;
					else if( x44 && ~x28 && x27 && x8 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( x44 && ~x28 && x27 && ~x8 && x37 )
						nx_state = s1;
					else if( x44 && ~x28 && x27 && ~x8 && ~x37 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x44 && ~x28 && ~x27 && x41 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x44 && ~x28 && ~x27 && ~x41 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s387;
						end
					else if( ~x44 && x10 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x44 && x10 && ~x4 )
						nx_state = s387;
					else if( ~x44 && ~x10 && x5 && x6 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x44 && ~x10 && x5 && ~x6 && x7 )
						nx_state = s1;
					else if( ~x44 && ~x10 && x5 && ~x6 && ~x7 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x44 && ~x10 && ~x5 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x44 && ~x10 && ~x5 && ~x4 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s387;
						end
					else nx_state = s387;
				s388 : if( x62 )
						nx_state = s1;
					else if( ~x62 && x14 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x62 && x14 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x62 && x14 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x62 && x14 && ~x23 )
						nx_state = s1;
					else if( ~x62 && ~x14 )
						begin
							y48 = 1'b1;	y57 = 1'b1;	y61 = 1'b1;	
							nx_state = s954;
						end
					else nx_state = s388;
				s389 : if( x62 && x20 && x18 && x17 && x19 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y17 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s389;
						end
					else if( x62 && x20 && x18 && x17 && ~x19 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x62 && x20 && x18 && ~x17 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x62 && x20 && ~x18 && x17 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x62 && x20 && ~x18 && ~x17 && x19 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x62 && x20 && ~x18 && ~x17 && ~x19 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x62 && ~x20 && x22 && x18 && x17 && x19 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y17 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s389;
						end
					else if( x62 && ~x20 && x22 && x18 && x17 && ~x19 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x62 && ~x20 && x22 && x18 && ~x17 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x62 && ~x20 && x22 && ~x18 && x17 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x62 && ~x20 && x22 && ~x18 && ~x17 && x19 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x62 && ~x20 && x22 && ~x18 && ~x17 && ~x19 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x62 && ~x20 && ~x22 && x21 && x18 && x17 && x19 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y17 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s389;
						end
					else if( x62 && ~x20 && ~x22 && x21 && x18 && x17 && ~x19 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x62 && ~x20 && ~x22 && x21 && x18 && ~x17 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x62 && ~x20 && ~x22 && x21 && ~x18 && x17 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x62 && ~x20 && ~x22 && x21 && ~x18 && ~x17 && x19 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x62 && ~x20 && ~x22 && x21 && ~x18 && ~x17 && ~x19 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x62 && ~x20 && ~x22 && ~x21 && x24 && x2 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x62 && ~x20 && ~x22 && ~x21 && x24 && x2 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x62 && ~x20 && ~x22 && ~x21 && x24 && ~x2 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x62 && ~x20 && ~x22 && ~x21 && ~x24 && x2 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( x62 && ~x20 && ~x22 && ~x21 && ~x24 && ~x2 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( x62 && ~x20 && ~x22 && ~x21 && ~x24 && ~x2 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x62 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s1074;
						end
					else nx_state = s389;
				s390 : if( x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x24 )
						begin
							y60 = 1'b1;	
							nx_state = s424;
						end
					else nx_state = s390;
				s391 : if( x63 )
						begin
							y53 = 1'b1;	
							nx_state = s1071;
						end
					else if( ~x63 && x65 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y54 = 1'b1;	
							nx_state = s1075;
						end
					else if( ~x63 && ~x65 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s1075;
						end
					else nx_state = s391;
				s392 : if( x63 && x19 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( x63 && ~x19 && x4 && x22 )
						begin
							y51 = 1'b1;	
							nx_state = s391;
						end
					else if( x63 && ~x19 && x4 && ~x22 )
						begin
							y44 = 1'b1;	y45 = 1'b1;	
							nx_state = s392;
						end
					else if( x63 && ~x19 && ~x4 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x63 && ~x19 && ~x4 && ~x18 )
						begin
							y44 = 1'b1;	y45 = 1'b1;	
							nx_state = s392;
						end
					else if( ~x63 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x63 && ~x6 )
						nx_state = s1;
					else nx_state = s392;
				s393 : if( x63 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x63 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && x20 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && x20 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x63 && ~x20 )
						nx_state = s1;
					else nx_state = s393;
				s394 : if( x63 )
						begin
							y23 = 1'b1;	y65 = 1'b1;	y72 = 1'b1;	
							nx_state = s1076;
						end
					else if( ~x63 && x21 && x22 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x63 && x21 && ~x22 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x63 && x21 && ~x22 && ~x23 )
						nx_state = s1;
					else if( ~x63 && ~x21 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x63 && ~x21 && ~x23 )
						nx_state = s1;
					else nx_state = s394;
				s395 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1077;
						end
					else nx_state = s395;
				s396 : if( x63 )
						nx_state = s1;
					else if( ~x63 && x14 && x65 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x63 && x14 && x65 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x63 && x14 && x65 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x63 && x14 && ~x65 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x63 && x14 && ~x65 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x63 && x14 && ~x65 && ~x15 && ~x16 )
						nx_state = s1;
					else if( ~x63 && ~x14 )
						nx_state = s1;
					else nx_state = s396;
				s397 : if( 1'b1 )
						begin
							y24 = 1'b1;	
							nx_state = s1012;
						end
					else nx_state = s397;
				s398 : if( 1'b1 )
						begin
							y21 = 1'b1;	
							nx_state = s822;
						end
					else nx_state = s398;
				s399 : if( x69 && x67 && x11 )
						nx_state = s1;
					else if( x69 && x67 && ~x11 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s64;
						end
					else if( x69 && x67 && ~x11 && ~x4 )
						nx_state = s399;
					else if( x69 && ~x67 && x10 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s64;
						end
					else if( x69 && ~x67 && x10 && ~x4 )
						nx_state = s399;
					else if( x69 && ~x67 && ~x10 && x15 )
						nx_state = s1;
					else if( x69 && ~x67 && ~x10 && ~x15 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s64;
						end
					else if( x69 && ~x67 && ~x10 && ~x15 && ~x4 )
						nx_state = s399;
					else if( ~x69 && x70 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x45 && x46 && x4 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x69 && ~x70 && x45 && x46 && ~x4 )
						nx_state = s399;
					else if( ~x69 && ~x70 && x45 && ~x46 && x12 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x45 && ~x46 && ~x12 && x4 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x69 && ~x70 && x45 && ~x46 && ~x12 && ~x4 )
						nx_state = s399;
					else if( ~x69 && ~x70 && ~x45 && x46 && x47 && x4 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x69 && ~x70 && ~x45 && x46 && x47 && ~x4 )
						nx_state = s399;
					else if( ~x69 && ~x70 && ~x45 && x46 && ~x47 && x4 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x69 && ~x70 && ~x45 && x46 && ~x47 && ~x4 )
						nx_state = s399;
					else if( ~x69 && ~x70 && ~x45 && ~x46 && x10 && x11 && x4 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x46 && x10 && x11 && ~x4 )
						nx_state = s399;
					else if( ~x69 && ~x70 && ~x45 && ~x46 && x10 && ~x11 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x45 && ~x46 && ~x10 && x12 && x4 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x69 && ~x70 && ~x45 && ~x46 && ~x10 && x12 && ~x4 )
						nx_state = s399;
					else if( ~x69 && ~x70 && ~x45 && ~x46 && ~x10 && ~x12 )
						nx_state = s1;
					else nx_state = s399;
				s400 : if( x63 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x63 && x65 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x63 && ~x65 && x66 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y57 = 1'b1;	
							nx_state = s1078;
						end
					else if( ~x63 && ~x65 && ~x66 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else nx_state = s400;
				s401 : if( x12 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( ~x12 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x12 && ~x13 )
						begin
							y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s572;
						end
					else nx_state = s401;
				s402 : if( x10 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x10 && x11 )
						begin
							y14 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s401;
						end
					else if( ~x10 && ~x11 )
						begin
							y10 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s402;
						end
					else nx_state = s402;
				s403 : if( x70 && x62 && x12 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && x62 && ~x12 )
						nx_state = s403;
					else if( x70 && ~x62 && x63 && x15 )
						begin
							y11 = 1'b1;	y24 = 1'b1;	
							nx_state = s1079;
						end
					else if( x70 && ~x62 && x63 && ~x15 && x12 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && ~x62 && x63 && ~x15 && ~x12 )
						nx_state = s403;
					else if( x70 && ~x62 && ~x63 && x64 && x20 && x7 && x6 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x20 && x7 && ~x6 && x5 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x20 && x7 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && x20 && ~x7 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x20 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && x65 && x66 && x68 && x21 && x20 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s1080;
						end
					else if( ~x70 && x65 && x66 && x68 && x21 && ~x20 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && x65 && x66 && x68 && ~x21 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && x65 && x66 && ~x68 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x70 && x65 && ~x66 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && ~x65 && x16 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && ~x65 && ~x16 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else nx_state = s403;
				s404 : if( x70 && x62 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x70 && x62 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x70 && x62 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x70 && x62 && ~x19 )
						nx_state = s1;
					else if( x70 && ~x62 && x63 && x23 && x22 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x70 && ~x62 && x63 && x23 && x22 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x70 && ~x62 && x63 && x23 && x22 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x70 && ~x62 && x63 && x23 && x22 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x70 && ~x62 && x63 && x23 && x22 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x70 && ~x62 && x63 && x23 && ~x22 && x19 && x20 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s523;
						end
					else if( x70 && ~x62 && x63 && x23 && ~x22 && x19 && ~x20 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s743;
						end
					else if( x70 && ~x62 && x63 && x23 && ~x22 && ~x19 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s742;
						end
					else if( x70 && ~x62 && x63 && ~x23 )
						begin
							y32 = 1'b1;	y33 = 1'b1;	
							nx_state = s396;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && x64 && ~x14 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && x65 && x67 && x24 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x65 && x67 && ~x24 && x11 && x12 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x65 && x67 && ~x24 && x11 && ~x12 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x65 && x67 && ~x24 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && x65 && x67 && ~x24 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && x65 && ~x67 && x29 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x65 && ~x67 && x29 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x65 && ~x67 && x29 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && x65 && ~x67 && x29 && ~x23 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && x65 && ~x67 && ~x29 )
						begin
							y8 = 1'b1;	
							nx_state = s373;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x65 && x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x65 && x26 && ~x25 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x65 && x26 && ~x25 && ~x24 )
						nx_state = s1;
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x65 && ~x26 )
						nx_state = s1;
					else if( ~x70 && x64 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x70 && ~x64 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s295;
						end
					else nx_state = s404;
				s405 : if( x69 && x70 && x63 && x23 && x22 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s1081;
						end
					else if( x69 && x70 && x63 && x23 && ~x22 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	y26 = 1'b1;	
							nx_state = s418;
						end
					else if( x69 && x70 && x63 && ~x23 && x22 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	y26 = 1'b1;	
							nx_state = s418;
						end
					else if( x69 && x70 && x63 && ~x23 && ~x22 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	y26 = 1'b1;	
							nx_state = s419;
						end
					else if( x69 && x70 && ~x63 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x69 && x70 && ~x63 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x69 && x70 && ~x63 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x69 && x70 && ~x63 && x22 && ~x23 )
						nx_state = s1;
					else if( x69 && x70 && ~x63 && ~x22 )
						nx_state = s1;
					else if( x69 && ~x70 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x69 && x25 )
						nx_state = s1;
					else if( ~x69 && ~x25 && x28 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s941;
						end
					else if( ~x69 && ~x25 && ~x28 )
						nx_state = s1;
					else nx_state = s405;
				s406 : if( x21 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x21 && x23 && x22 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x21 && x23 && ~x22 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( ~x21 && x23 && ~x22 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( ~x21 && x23 && ~x22 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x23 && ~x22 && ~x20 )
						nx_state = s1;
					else if( ~x21 && ~x23 && x18 && x14 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x21 && ~x23 && x18 && x14 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x21 && ~x23 && x18 && ~x14 && x13 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x21 && ~x23 && x18 && ~x14 && x13 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x21 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x23 && ~x18 )
						nx_state = s1;
					else nx_state = s406;
				s407 : if( x20 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( ~x20 && x21 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x20 && ~x21 )
						nx_state = s1;
					else nx_state = s407;
				s408 : if( x44 && x37 && x28 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x44 && x37 && ~x28 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x44 && ~x37 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x44 && x10 && x1 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x44 && x10 && ~x1 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x44 && ~x10 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else nx_state = s408;
				s409 : if( 1'b1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y40 = 1'b1;	
							y42 = 1'b1;	
							nx_state = s1082;
						end
					else nx_state = s409;
				s410 : if( x62 )
						nx_state = s1;
					else if( ~x62 && x63 && x20 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x62 && x63 && ~x20 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x62 && x63 && ~x20 && ~x18 )
						begin
							y44 = 1'b1;	y45 = 1'b1;	
							nx_state = s392;
						end
					else if( ~x62 && ~x63 && x64 && x65 && x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x62 && ~x63 && x64 && x65 && x10 && ~x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x62 && ~x63 && x64 && x65 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && x65 && ~x10 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && ~x65 && x66 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && ~x63 && x64 && ~x65 && x66 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && ~x63 && x64 && ~x65 && x66 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && ~x65 && x66 && ~x9 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && ~x65 && ~x66 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x62 && ~x63 && x64 && ~x65 && ~x66 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x62 && ~x63 && x64 && ~x65 && ~x66 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && ~x65 && ~x66 && ~x18 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 )
						begin
							y38 = 1'b1;	
							nx_state = s845;
						end
					else nx_state = s410;
				s411 : if( 1'b1 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s693;
						end
					else nx_state = s411;
				s412 : if( x21 && x12 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x21 && x12 && ~x8 && x7 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x21 && x12 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x21 && ~x12 )
						nx_state = s1;
					else if( ~x21 && x7 && x6 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && x7 && ~x6 && x5 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && x7 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x21 && ~x7 )
						nx_state = s1;
					else nx_state = s412;
				s413 : if( x63 )
						begin
							y27 = 1'b1;	
							nx_state = s1083;
						end
					else if( ~x63 && x65 && x21 && x17 && x16 && x19 && x11 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x63 && x65 && x21 && x17 && x16 && x19 && ~x11 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x65 && x21 && x17 && x16 && ~x19 && x18 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x63 && x65 && x21 && x17 && x16 && ~x19 && ~x18 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x65 && x21 && x17 && ~x16 && x11 )
						begin
							y3 = 1'b1;	
							nx_state = s788;
						end
					else if( ~x63 && x65 && x21 && x17 && ~x16 && ~x11 )
						begin
							y32 = 1'b1;	
							nx_state = s854;
						end
					else if( ~x63 && x65 && x21 && ~x17 && x16 && x19 && x14 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x63 && x65 && x21 && ~x17 && x16 && x19 && ~x14 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x65 && x21 && ~x17 && x16 && ~x19 && x13 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x63 && x65 && x21 && ~x17 && x16 && ~x19 && ~x13 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x65 && x21 && ~x17 && ~x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x65 && ~x21 )
						begin
							y30 = 1'b1;	
							nx_state = s416;
						end
					else if( ~x63 && ~x65 )
						begin
							y5 = 1'b1;	y13 = 1'b1;	y17 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1084;
						end
					else nx_state = s413;
				s414 : if( x64 && x17 && x16 && x19 && x11 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x64 && x17 && x16 && x19 && ~x11 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x64 && x17 && x16 && ~x19 && x18 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x64 && x17 && x16 && ~x19 && ~x18 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x64 && x17 && ~x16 && x11 )
						begin
							y3 = 1'b1;	
							nx_state = s788;
						end
					else if( x64 && x17 && ~x16 && ~x11 )
						begin
							y32 = 1'b1;	
							nx_state = s854;
						end
					else if( x64 && ~x17 && x16 && x19 && x14 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x64 && ~x17 && x16 && x19 && ~x14 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x64 && ~x17 && x16 && ~x19 && x13 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x64 && ~x17 && x16 && ~x19 && ~x13 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x64 && ~x17 && ~x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x64 && x30 )
						begin
							y3 = 1'b1;	
							nx_state = s788;
						end
					else if( ~x64 && ~x30 && x4 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x64 && ~x30 && ~x4 )
						begin
							y5 = 1'b1;	
							nx_state = s791;
						end
					else nx_state = s414;
				s415 : if( x7 && x6 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x7 && ~x6 && x5 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x7 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x7 )
						nx_state = s1;
					else nx_state = s415;
				s416 : if( x62 )
						begin
							y6 = 1'b1;	y47 = 1'b1;	
							nx_state = s1085;
						end
					else if( ~x62 && x64 )
						nx_state = s47;
					else if( ~x62 && ~x64 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else nx_state = s416;
				s417 : if( x63 )
						begin
							y60 = 1'b1;	
							nx_state = s424;
						end
					else if( ~x63 )
						nx_state = s1;
					else nx_state = s417;
				s418 : if( x23 && x17 && x22 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s1086;
						end
					else if( x23 && x17 && ~x22 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s1087;
						end
					else if( x23 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1088;
						end
					else if( ~x23 && x22 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s1087;
						end
					else if( ~x23 && x22 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1088;
						end
					else if( ~x23 && ~x22 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s1086;
						end
					else if( ~x23 && ~x22 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1089;
						end
					else nx_state = s418;
				s419 : if( x22 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s1086;
						end
					else if( x22 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1090;
						end
					else if( ~x22 && x23 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s1086;
						end
					else if( ~x22 && x23 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1091;
						end
					else if( ~x22 && ~x23 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s1092;
						end
					else if( ~x22 && ~x23 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1088;
						end
					else nx_state = s419;
				s420 : if( x24 )
						nx_state = s1;
					else if( ~x24 && x23 && x10 )
						begin
							y25 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x24 && x23 && ~x10 )
						begin
							y23 = 1'b1;	
							nx_state = s588;
						end
					else if( ~x24 && ~x23 )
						nx_state = s1;
					else nx_state = s420;
				s421 : if( x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( ~x21 && x15 && x10 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x21 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s605;
						end
					else if( ~x21 && x15 && x10 && ~x11 && ~x12 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s606;
						end
					else if( ~x21 && x15 && ~x10 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( ~x21 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s600;
						end
					else if( ~x21 && ~x15 && x16 && x10 && x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y11 = 1'b1;	
							nx_state = s600;
						end
					else if( ~x21 && ~x15 && x16 && x10 && ~x12 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( ~x21 && ~x15 && x16 && ~x10 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y11 = 1'b1;	
							nx_state = s600;
						end
					else if( ~x21 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s607;
						end
					else nx_state = s421;
				s422 : if( x69 && x63 && x19 && x18 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1093;
						end
					else if( x69 && x63 && x19 && ~x18 )
						begin
							y25 = 1'b1;	y29 = 1'b1;	y48 = 1'b1;	
							nx_state = s820;
						end
					else if( x69 && x63 && ~x19 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1094;
						end
					else if( x69 && ~x63 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y20 = 1'b1;	
							nx_state = s1095;
						end
					else if( ~x69 && x38 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( ~x69 && ~x38 )
						nx_state = s422;
					else nx_state = s422;
				s423 : if( x69 && x66 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x69 && ~x66 && x22 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s1096;
						end
					else if( x69 && ~x66 && ~x22 && x23 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s1081;
						end
					else if( x69 && ~x66 && ~x22 && ~x23 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s1096;
						end
					else if( ~x69 && x10 && x61 && x12 && x23 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x69 && x10 && x61 && x12 && ~x23 && x4 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x69 && x10 && x61 && x12 && ~x23 && ~x4 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( ~x69 && x10 && x61 && ~x12 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s215;
						end
					else if( ~x69 && x10 && ~x61 && x39 && x46 && x51 && x36 )
						nx_state = s423;
					else if( ~x69 && x10 && ~x61 && x39 && x46 && x51 && ~x36 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x69 && x10 && ~x61 && x39 && x46 && ~x51 && x36 )
						nx_state = s423;
					else if( ~x69 && x10 && ~x61 && x39 && x46 && ~x51 && ~x36 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s840;
						end
					else if( ~x69 && x10 && ~x61 && x39 && ~x46 && x36 )
						nx_state = s423;
					else if( ~x69 && x10 && ~x61 && x39 && ~x46 && ~x36 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s1097;
						end
					else if( ~x69 && x10 && ~x61 && ~x39 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s874;
						end
					else if( ~x69 && ~x10 && x61 && x1 && x22 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							nx_state = s869;
						end
					else if( ~x69 && ~x10 && x61 && x1 && ~x22 && x2 && x11 && x5 && x3 )
						nx_state = s423;
					else if( ~x69 && ~x10 && x61 && x1 && ~x22 && x2 && x11 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s840;
						end
					else if( ~x69 && ~x10 && x61 && x1 && ~x22 && x2 && x11 && ~x5 && x3 )
						nx_state = s423;
					else if( ~x69 && ~x10 && x61 && x1 && ~x22 && x2 && x11 && ~x5 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( ~x69 && ~x10 && x61 && x1 && ~x22 && x2 && ~x11 && x3 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( ~x69 && ~x10 && x61 && x1 && ~x22 && x2 && ~x11 && ~x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x69 && ~x10 && x61 && x1 && ~x22 && ~x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s1097;
						end
					else if( ~x69 && ~x10 && x61 && ~x1 && x11 && x4 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( ~x69 && ~x10 && x61 && ~x1 && x11 && ~x4 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( ~x69 && ~x10 && x61 && ~x1 && ~x11 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( ~x69 && ~x10 && ~x61 && x11 && x34 && x8 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s733;
						end
					else if( ~x69 && ~x10 && ~x61 && x11 && x34 && ~x8 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x69 && ~x10 && ~x61 && x11 && x34 && ~x8 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( ~x69 && ~x10 && ~x61 && x11 && ~x34 && x32 && x7 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s733;
						end
					else if( ~x69 && ~x10 && ~x61 && x11 && ~x34 && x32 && ~x7 && x54 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x69 && ~x10 && ~x61 && x11 && ~x34 && x32 && ~x7 && x54 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( ~x69 && ~x10 && ~x61 && x11 && ~x34 && x32 && ~x7 && ~x54 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s1097;
						end
					else if( ~x69 && ~x10 && ~x61 && x11 && ~x34 && ~x32 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( ~x69 && ~x10 && ~x61 && ~x11 && x12 && x20 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s1097;
						end
					else if( ~x69 && ~x10 && ~x61 && ~x11 && x12 && ~x20 && x2 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( ~x69 && ~x10 && ~x61 && ~x11 && x12 && ~x20 && ~x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x69 && ~x10 && ~x61 && ~x11 && ~x12 && x13 && x1 && x3 && x6 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s215;
						end
					else if( ~x69 && ~x10 && ~x61 && ~x11 && ~x12 && x13 && x1 && x3 && ~x6 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( ~x69 && ~x10 && ~x61 && ~x11 && ~x12 && x13 && x1 && ~x3 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( ~x69 && ~x10 && ~x61 && ~x11 && ~x12 && x13 && ~x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s1097;
						end
					else if( ~x69 && ~x10 && ~x61 && ~x11 && ~x12 && ~x13 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s840;
						end
					else nx_state = s423;
				s424 : if( x63 && x65 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x63 && ~x65 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x65 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x65 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x63 && ~x65 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x65 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x63 )
						begin
							y61 = 1'b1;	
							nx_state = s1098;
						end
					else nx_state = s424;
				s425 : if( 1'b1 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1099;
						end
					else nx_state = s425;
				s426 : if( x70 && x64 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( x70 && ~x64 && x1 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x70 && ~x64 && x1 && ~x2 && x5 && x3 )
						nx_state = s426;
					else if( x70 && ~x64 && x1 && ~x2 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x70 && ~x64 && x1 && ~x2 && ~x5 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	
							nx_state = s7;
						end
					else if( x70 && ~x64 && ~x1 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( ~x70 && x67 && x22 )
						begin
							y2 = 1'b1;	y16 = 1'b1;	y24 = 1'b1;	
							nx_state = s270;
						end
					else if( ~x70 && x67 && ~x22 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( ~x70 && ~x67 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else nx_state = s426;
				s427 : if( 1'b1 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else nx_state = s427;
				s428 : if( x69 && x21 && x15 && x16 && x9 && x7 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && x21 && x15 && x16 && x9 && ~x7 && x8 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s296;
						end
					else if( x69 && x21 && x15 && x16 && x9 && ~x7 && ~x8 && x13 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x69 && x21 && x15 && x16 && x9 && ~x7 && ~x8 && ~x13 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && x21 && x15 && x16 && x9 && ~x7 && ~x8 && ~x13 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x21 && x15 && x16 && x9 && ~x7 && ~x8 && ~x13 && ~x18 && x19 && ~x14 )
						nx_state = s1;
					else if( x69 && x21 && x15 && x16 && x9 && ~x7 && ~x8 && ~x13 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && x21 && x15 && x16 && ~x9 && x7 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && x21 && x15 && x16 && ~x9 && ~x7 && x8 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s297;
						end
					else if( x69 && x21 && x15 && x16 && ~x9 && ~x7 && ~x8 && x14 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x69 && x21 && x15 && x16 && ~x9 && ~x7 && ~x8 && ~x14 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && x21 && x15 && ~x16 && x7 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s406;
						end
					else if( x69 && x21 && x15 && ~x16 && ~x7 && x8 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s406;
						end
					else if( x69 && x21 && x15 && ~x16 && ~x7 && ~x8 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x69 && x21 && x15 && ~x16 && ~x7 && ~x8 && ~x2 && x5 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && x21 && x15 && ~x16 && ~x7 && ~x8 && ~x2 && ~x5 && x9 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x69 && x21 && x15 && ~x16 && ~x7 && ~x8 && ~x2 && ~x5 && ~x9 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x69 && x21 && ~x15 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x69 && x21 && ~x15 && ~x2 && x16 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x21 && ~x15 && ~x2 && x16 && x9 && ~x10 && x8 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x21 && ~x15 && ~x2 && x16 && x9 && ~x10 && ~x8 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && x21 && ~x15 && ~x2 && x16 && x9 && ~x10 && ~x8 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x21 && ~x15 && ~x2 && x16 && x9 && ~x10 && ~x8 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x21 && ~x15 && ~x2 && x16 && x9 && ~x10 && ~x8 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && x21 && ~x15 && ~x2 && x16 && x9 && ~x10 && ~x8 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && x21 && ~x15 && ~x2 && x16 && ~x9 && x8 && x12 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x21 && ~x15 && ~x2 && x16 && ~x9 && x8 && ~x12 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && x21 && ~x15 && ~x2 && x16 && ~x9 && x8 && ~x12 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x21 && ~x15 && ~x2 && x16 && ~x9 && x8 && ~x12 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x21 && ~x15 && ~x2 && x16 && ~x9 && x8 && ~x12 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && x21 && ~x15 && ~x2 && x16 && ~x9 && x8 && ~x12 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && x21 && ~x15 && ~x2 && x16 && ~x9 && ~x8 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x21 && ~x15 && ~x2 && x16 && ~x9 && ~x8 && ~x11 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x69 && x21 && ~x15 && ~x2 && x16 && ~x9 && ~x8 && ~x11 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x21 && ~x15 && ~x2 && x16 && ~x9 && ~x8 && ~x11 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x21 && ~x15 && ~x2 && x16 && ~x9 && ~x8 && ~x11 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && x21 && ~x15 && ~x2 && x16 && ~x9 && ~x8 && ~x11 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x69 && x21 && ~x15 && ~x2 && ~x16 && x5 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && x21 && ~x15 && ~x2 && ~x16 && ~x5 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s495;
						end
					else if( x69 && ~x21 && x22 && x18 && x14 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x21 && x22 && x18 && ~x14 && x13 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x21 && x22 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x21 && x22 && ~x18 )
						nx_state = s1;
					else if( x69 && ~x21 && ~x22 )
						nx_state = s1;
					else if( ~x69 && x12 && x15 && x13 && x3 )
						begin
							y13 = 1'b1;	
							nx_state = s763;
						end
					else if( ~x69 && x12 && x15 && x13 && ~x3 && x14 )
						begin
							y13 = 1'b1;	
							nx_state = s763;
						end
					else if( ~x69 && x12 && x15 && x13 && ~x3 && ~x14 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s764;
						end
					else if( ~x69 && x12 && x15 && ~x13 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s765;
						end
					else if( ~x69 && x12 && ~x15 )
						begin
							y10 = 1'b1;	
							nx_state = s766;
						end
					else if( ~x69 && ~x12 )
						begin
							y10 = 1'b1;	
							nx_state = s766;
						end
					else nx_state = s428;
				s429 : if( x68 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x68 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x68 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x68 && x20 && ~x18 )
						nx_state = s1;
					else if( x68 && ~x20 && x21 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x68 && ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( x68 && ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( x68 && ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x68 && ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else if( ~x68 && x24 && x26 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x68 && x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x68 && x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x68 && x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x68 && x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x68 && ~x24 && x25 && x26 && x15 && x10 && x11 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s300;
						end
					else if( ~x68 && ~x24 && x25 && x26 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s1038;
						end
					else if( ~x68 && ~x24 && x25 && x26 && x15 && x10 && ~x11 && ~x12 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s300;
						end
					else if( ~x68 && ~x24 && x25 && x26 && x15 && ~x10 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s1039;
						end
					else if( ~x68 && ~x24 && x25 && x26 && ~x15 && x16 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s497;
						end
					else if( ~x68 && ~x24 && x25 && x26 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( ~x68 && ~x24 && x25 && ~x26 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && x19 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && x20 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && ~x20 && x21 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && ~x20 && ~x21 && x22 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && ~x20 && ~x21 && ~x22 && x16 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && ~x20 && ~x21 && ~x22 && x16 && ~x11 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && ~x20 && ~x21 && ~x22 && x16 && ~x11 && ~x12 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && ~x20 && ~x21 && ~x22 && x16 && ~x11 && ~x12 && ~x10 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && ~x20 && ~x21 && ~x22 && ~x16 && x17 && x10 && x12 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && ~x20 && ~x21 && ~x22 && ~x16 && x17 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && ~x20 && ~x21 && ~x22 && ~x16 && x17 && ~x10 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && ~x20 && ~x21 && ~x22 && ~x16 && ~x17 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x68 && ~x24 && ~x25 && ~x26 && x15 && x12 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x68 && ~x24 && ~x25 && ~x26 && x15 && ~x12 && x11 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x68 && ~x24 && ~x25 && ~x26 && x15 && ~x12 && ~x11 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x68 && ~x24 && ~x25 && ~x26 && x15 && ~x12 && ~x11 && ~x10 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( ~x68 && ~x24 && ~x25 && ~x26 && ~x15 && x16 && x10 && x12 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s497;
						end
					else if( ~x68 && ~x24 && ~x25 && ~x26 && ~x15 && x16 && x10 && ~x12 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s899;
						end
					else if( ~x68 && ~x24 && ~x25 && ~x26 && ~x15 && x16 && ~x10 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s497;
						end
					else if( ~x68 && ~x24 && ~x25 && ~x26 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else nx_state = s429;
				s430 : if( x24 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( x24 && ~x4 && x20 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x24 && ~x4 && ~x20 && x21 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x24 && ~x4 && ~x20 && ~x21 && x22 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x24 && ~x4 && ~x20 && ~x21 && ~x22 && x23 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x24 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && x16 && x11 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( x24 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && x16 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x24 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && x13 && x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x24 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && x13 && ~x11 && x12 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( x24 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && x13 && ~x11 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x24 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && ~x13 && x11 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x24 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && ~x13 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x24 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s35;
						end
					else if( ~x24 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x19 && ~x14 && ~x13 )
						nx_state = s430;
					else if( ~x24 && ~x19 )
						nx_state = s1;
					else nx_state = s430;
				s431 : if( x70 && x62 )
						begin
							y5 = 1'b1;	
							nx_state = s791;
						end
					else if( x70 && ~x62 && x63 && x16 && x22 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1100;
						end
					else if( x70 && ~x62 && x63 && x16 && x22 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s523;
						end
					else if( x70 && ~x62 && x63 && x16 && ~x22 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s442;
						end
					else if( x70 && ~x62 && x63 && ~x16 && x22 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s524;
						end
					else if( x70 && ~x62 && x63 && ~x16 && ~x22 )
						begin
							y3 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s520;
						end
					else if( x70 && ~x62 && ~x63 )
						begin
							y7 = 1'b1;	
							nx_state = s82;
						end
					else if( ~x70 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else nx_state = s431;
				s432 : if( x26 )
						begin
							y14 = 1'b1;	
							nx_state = s124;
						end
					else if( ~x26 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else nx_state = s432;
				s433 : if( 1'b1 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else nx_state = s433;
				s434 : if( x69 && x65 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( x69 && ~x65 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s225;
						end
					else if( ~x69 && x62 && x61 && x19 && x28 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && x62 && x61 && x19 && x28 && ~x1 && x35 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s840;
						end
					else if( ~x69 && x62 && x61 && x19 && x28 && ~x1 && ~x35 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( ~x69 && x62 && x61 && x19 && ~x28 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( ~x69 && x62 && x61 && ~x19 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( ~x69 && x62 && ~x61 && x13 && x23 && x51 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x69 && x62 && ~x61 && x13 && x23 && ~x51 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s840;
						end
					else if( ~x69 && x62 && ~x61 && x13 && ~x23 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x69 && x62 && ~x61 && ~x13 && x28 && x35 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x69 && x62 && ~x61 && ~x13 && x28 && x35 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( ~x69 && x62 && ~x61 && ~x13 && x28 && ~x35 && x60 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( ~x69 && x62 && ~x61 && ~x13 && x28 && ~x35 && ~x60 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( ~x69 && x62 && ~x61 && ~x13 && ~x28 && x6 && x35 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x69 && x62 && ~x61 && ~x13 && ~x28 && x6 && ~x35 && x60 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( ~x69 && x62 && ~x61 && ~x13 && ~x28 && x6 && ~x35 && ~x60 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( ~x69 && x62 && ~x61 && ~x13 && ~x28 && ~x6 && x39 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( ~x69 && x62 && ~x61 && ~x13 && ~x28 && ~x6 && ~x39 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x69 && ~x62 && x55 && x50 && x28 && x32 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s739;
						end
					else if( ~x69 && ~x62 && x55 && x50 && x28 && ~x32 && x35 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && ~x62 && x55 && x50 && x28 && ~x32 && ~x35 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( ~x69 && ~x62 && x55 && x50 && ~x28 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( ~x69 && ~x62 && x55 && ~x50 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( ~x69 && ~x62 && ~x55 && x13 && x23 && x51 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s906;
						end
					else if( ~x69 && ~x62 && ~x55 && x13 && x23 && ~x51 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && ~x62 && ~x55 && x13 && ~x23 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s906;
						end
					else if( ~x69 && ~x62 && ~x55 && ~x13 && x28 && x35 && x36 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s906;
						end
					else if( ~x69 && ~x62 && ~x55 && ~x13 && x28 && x35 && ~x36 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( ~x69 && ~x62 && ~x55 && ~x13 && x28 && ~x35 && x58 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( ~x69 && ~x62 && ~x55 && ~x13 && x28 && ~x35 && ~x58 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( ~x69 && ~x62 && ~x55 && ~x13 && ~x28 && x6 && x35 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s443;
						end
					else if( ~x69 && ~x62 && ~x55 && ~x13 && ~x28 && x6 && ~x35 && x58 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( ~x69 && ~x62 && ~x55 && ~x13 && ~x28 && x6 && ~x35 && ~x58 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( ~x69 && ~x62 && ~x55 && ~x13 && ~x28 && ~x6 && x39 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( ~x69 && ~x62 && ~x55 && ~x13 && ~x28 && ~x6 && ~x39 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s734;
						end
					else nx_state = s434;
				s435 : if( x66 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x66 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s306;
						end
					else nx_state = s435;
				s436 : if( x15 && x16 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x15 && ~x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x15 && x16 && x4 && x5 && x1 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s448;
						end
					else if( ~x15 && x16 && x4 && x5 && ~x1 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else if( ~x15 && x16 && x4 && ~x5 && x2 && x3 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s928;
						end
					else if( ~x15 && x16 && x4 && ~x5 && x2 && ~x3 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else if( ~x15 && x16 && x4 && ~x5 && ~x2 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s900;
						end
					else if( ~x15 && x16 && ~x4 && x2 && x3 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s194;
						end
					else if( ~x15 && x16 && ~x4 && x2 && ~x3 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else if( ~x15 && x16 && ~x4 && ~x2 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s900;
						end
					else if( ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s194;
						end
					else nx_state = s436;
				s437 : if( x69 && x63 && x19 && x18 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1101;
						end
					else if( x69 && x63 && x19 && ~x18 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1102;
						end
					else if( x69 && x63 && ~x19 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s821;
						end
					else if( x69 && ~x63 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							nx_state = s1103;
						end
					else if( ~x69 && x15 && x16 && x5 && x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s451;
						end
					else if( ~x69 && x15 && x16 && x5 && ~x1 && x2 && x3 && x4 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s448;
						end
					else if( ~x69 && x15 && x16 && x5 && ~x1 && x2 && x3 && ~x4 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x15 && x16 && x5 && ~x1 && x2 && ~x3 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x15 && x16 && x5 && ~x1 && ~x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x15 && x16 && ~x5 && x6 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x15 && x16 && ~x5 && ~x6 && x1 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s436;
						end
					else if( ~x69 && x15 && x16 && ~x5 && ~x6 && ~x1 && x2 && x3 && x4 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s448;
						end
					else if( ~x69 && x15 && x16 && ~x5 && ~x6 && ~x1 && x2 && x3 && ~x4 )
						begin
							y10 = 1'b1;	
							nx_state = s193;
						end
					else if( ~x69 && x15 && x16 && ~x5 && ~x6 && ~x1 && x2 && ~x3 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x15 && x16 && ~x5 && ~x6 && ~x1 && ~x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x15 && ~x16 && x6 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && x15 && ~x16 && ~x6 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s438;
						end
					else if( ~x69 && ~x15 && x16 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s901;
						end
					else if( ~x69 && ~x15 && ~x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else nx_state = s437;
				s438 : if( x69 )
						begin
							y8 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s172;
						end
					else if( ~x69 && x16 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x16 && x15 && x8 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && ~x16 && x15 && ~x8 && x9 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && ~x16 && x15 && ~x8 && ~x9 && x10 && x6 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x16 && x15 && ~x8 && ~x9 && x10 && ~x6 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s438;
						end
					else if( ~x69 && ~x16 && x15 && ~x8 && ~x9 && ~x10 && x11 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s436;
						end
					else if( ~x69 && ~x16 && x15 && ~x8 && ~x9 && ~x10 && ~x11 )
						nx_state = s438;
					else if( ~x69 && ~x16 && ~x15 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else nx_state = s438;
				s439 : if( x63 && x46 && x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x63 && x46 && x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x63 && x46 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x63 && ~x46 && x47 && x4 && x5 && x1 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s453;
						end
					else if( x63 && ~x46 && x47 && x4 && x5 && ~x1 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s440;
						end
					else if( x63 && ~x46 && x47 && x4 && ~x5 && x2 && x3 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s932;
						end
					else if( x63 && ~x46 && x47 && x4 && ~x5 && x2 && ~x3 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s440;
						end
					else if( x63 && ~x46 && x47 && x4 && ~x5 && ~x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( x63 && ~x46 && x47 && ~x4 && x33 && x34 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( x63 && ~x46 && x47 && ~x4 && x33 && ~x34 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s440;
						end
					else if( x63 && ~x46 && x47 && ~x4 && ~x33 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( x63 && ~x46 && ~x47 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x63 && x16 && x15 && x64 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x63 && x16 && x15 && x64 && ~x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x63 && x16 && x15 && ~x64 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x63 && x16 && x15 && ~x64 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x63 && x16 && ~x15 && x4 && x5 && x1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s455;
						end
					else if( ~x63 && x16 && ~x15 && x4 && x5 && ~x1 && x64 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s445;
						end
					else if( ~x63 && x16 && ~x15 && x4 && x5 && ~x1 && ~x64 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s931;
						end
					else if( ~x63 && x16 && ~x15 && x4 && ~x5 && x2 && x3 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s932;
						end
					else if( ~x63 && x16 && ~x15 && x4 && ~x5 && x2 && ~x3 && x64 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s445;
						end
					else if( ~x63 && x16 && ~x15 && x4 && ~x5 && x2 && ~x3 && ~x64 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s931;
						end
					else if( ~x63 && x16 && ~x15 && x4 && ~x5 && ~x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( ~x63 && x16 && ~x15 && ~x4 && x64 && x2 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x63 && x16 && ~x15 && ~x4 && x64 && x2 && ~x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s445;
						end
					else if( ~x63 && x16 && ~x15 && ~x4 && x64 && ~x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( ~x63 && x16 && ~x15 && ~x4 && ~x64 && x34 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x63 && x16 && ~x15 && ~x4 && ~x64 && x34 && ~x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s931;
						end
					else if( ~x63 && x16 && ~x15 && ~x4 && ~x64 && ~x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( ~x63 && ~x16 && x15 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x63 && ~x16 && ~x15 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else nx_state = s439;
				s440 : if( x46 && x16 && x36 && x1 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s322;
						end
					else if( x46 && x16 && x36 && ~x1 && x2 && x3 && x35 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s453;
						end
					else if( x46 && x16 && x36 && ~x1 && x2 && x3 && ~x35 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x46 && x16 && x36 && ~x1 && x2 && ~x3 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x46 && x16 && x36 && ~x1 && ~x2 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x46 && x16 && ~x36 && x6 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x46 && x16 && ~x36 && ~x6 && x32 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( x46 && x16 && ~x36 && ~x6 && ~x32 && x33 && x34 && x4 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s453;
						end
					else if( x46 && x16 && ~x36 && ~x6 && ~x32 && x33 && x34 && ~x4 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( x46 && x16 && ~x36 && ~x6 && ~x32 && x33 && ~x34 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x46 && x16 && ~x36 && ~x6 && ~x32 && ~x33 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x46 && ~x16 && x37 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x46 && ~x16 && ~x37 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s442;
						end
					else if( ~x46 && x47 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( ~x46 && ~x47 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else nx_state = s440;
				s441 : if( x69 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x69 && x63 && x46 && x16 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && x63 && x46 && ~x16 && x42 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x63 && x46 && ~x16 && ~x42 && x10 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s453;
						end
					else if( ~x69 && x63 && x46 && ~x16 && ~x42 && ~x10 )
						nx_state = s441;
					else if( ~x69 && x63 && ~x46 && x47 && x3 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s322;
						end
					else if( ~x69 && x63 && ~x46 && x47 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s929;
						end
					else if( ~x69 && x63 && ~x46 && ~x47 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x69 && ~x63 && x16 && x15 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && ~x63 && x16 && ~x15 && x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s326;
						end
					else if( ~x69 && ~x63 && x16 && ~x15 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s929;
						end
					else if( ~x69 && ~x63 && ~x16 && x15 && x11 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && ~x63 && ~x16 && x15 && ~x11 && x10 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s455;
						end
					else if( ~x69 && ~x63 && ~x16 && x15 && ~x11 && ~x10 )
						nx_state = s441;
					else if( ~x69 && ~x63 && ~x16 && ~x15 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else nx_state = s441;
				s442 : if( x69 && x23 )
						begin
							y19 = 1'b1;	
							nx_state = s13;
						end
					else if( x69 && ~x23 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( ~x69 && x16 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x16 && x15 && x39 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s441;
						end
					else if( ~x69 && ~x16 && x15 && ~x39 && x9 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s441;
						end
					else if( ~x69 && ~x16 && x15 && ~x39 && ~x9 && x41 && x37 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x16 && x15 && ~x39 && ~x9 && x41 && ~x37 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s442;
						end
					else if( ~x69 && ~x16 && x15 && ~x39 && ~x9 && ~x41 && x42 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && ~x16 && x15 && ~x39 && ~x9 && ~x41 && ~x42 )
						nx_state = s442;
					else if( ~x69 && ~x16 && ~x15 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else nx_state = s442;
				s443 : if( x69 && x21 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x69 && ~x21 && x22 && x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x21 && x22 && ~x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s107;
						end
					else if( x69 && ~x21 && ~x22 && x8 && x16 && x15 && x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x21 && ~x22 && x8 && x16 && x15 && ~x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s828;
						end
					else if( x69 && ~x21 && ~x22 && x8 && x16 && ~x15 && x10 )
						begin
							y2 = 1'b1;	y16 = 1'b1;	y24 = 1'b1;	
							nx_state = s270;
						end
					else if( x69 && ~x21 && ~x22 && x8 && x16 && ~x15 && ~x10 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s267;
						end
					else if( x69 && ~x21 && ~x22 && x8 && ~x16 && x17 && x10 && x15 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x21 && ~x22 && x8 && ~x16 && x17 && x10 && ~x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s827;
						end
					else if( x69 && ~x21 && ~x22 && x8 && ~x16 && x17 && ~x10 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s149;
						end
					else if( x69 && ~x21 && ~x22 && x8 && ~x16 && ~x17 && x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x21 && ~x22 && x8 && ~x16 && ~x17 && ~x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s829;
						end
					else if( x69 && ~x21 && ~x22 && ~x8 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( ~x69 && x70 && x63 && x64 && x55 && x40 )
						begin
							y13 = 1'b1;	
							nx_state = s450;
						end
					else if( ~x69 && x70 && x63 && x64 && x55 && ~x40 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && x70 && x63 && x64 && x55 && ~x40 && ~x3 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s734;
						end
					else if( ~x69 && x70 && x63 && x64 && ~x55 && x29 && x50 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s910;
						end
					else if( ~x69 && x70 && x63 && x64 && ~x55 && x29 && ~x50 )
						nx_state = s443;
					else if( ~x69 && x70 && x63 && x64 && ~x55 && ~x29 && x58 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( ~x69 && x70 && x63 && x64 && ~x55 && ~x29 && ~x58 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( ~x69 && x70 && x63 && ~x64 && x15 && x9 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && x70 && x63 && ~x64 && x15 && ~x9 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && x70 && x63 && ~x64 && x15 && ~x9 && ~x3 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x70 && x63 && ~x64 && ~x15 && x29 && x49 )
						begin
							y12 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s912;
						end
					else if( ~x69 && x70 && x63 && ~x64 && ~x15 && x29 && ~x49 )
						nx_state = s443;
					else if( ~x69 && x70 && x63 && ~x64 && ~x15 && ~x29 && x21 )
						nx_state = s1;
					else if( ~x69 && x70 && x63 && ~x64 && ~x15 && ~x29 && ~x21 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && x70 && ~x63 && x40 && x9 )
						begin
							y13 = 1'b1;	
							nx_state = s450;
						end
					else if( ~x69 && x70 && ~x63 && x40 && ~x9 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && x70 && ~x63 && x40 && ~x9 && ~x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s736;
						end
					else if( ~x69 && x70 && ~x63 && ~x40 && x29 && x50 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s910;
						end
					else if( ~x69 && x70 && ~x63 && ~x40 && x29 && ~x50 )
						nx_state = s443;
					else if( ~x69 && x70 && ~x63 && ~x40 && ~x29 && x41 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x69 && x70 && ~x63 && ~x40 && ~x29 && ~x41 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( ~x69 && ~x70 && x9 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && ~x70 && ~x9 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && ~x70 && ~x9 && ~x3 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else nx_state = s443;
				s444 : if( x69 && x62 && x13 && x20 )
						nx_state = s1;
					else if( x69 && x62 && x13 && ~x20 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && x62 && ~x13 && x12 )
						nx_state = s1;
					else if( x69 && x62 && ~x13 && ~x12 && x10 && x3 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && x62 && ~x13 && ~x12 && x10 && ~x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s540;
						end
					else if( x69 && x62 && ~x13 && ~x12 && ~x10 && x19 && x16 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( x69 && x62 && ~x13 && ~x12 && ~x10 && x19 && ~x16 )
						nx_state = s1;
					else if( x69 && x62 && ~x13 && ~x12 && ~x10 && ~x19 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( x69 && ~x62 && x18 && x17 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && ~x62 && x18 && x17 && ~x1 && x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && x18 && x17 && ~x1 && ~x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && ~x62 && x18 && ~x17 && x3 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && ~x62 && x18 && ~x17 && ~x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s540;
						end
					else if( x69 && ~x62 && ~x18 && x17 && x7 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( x69 && ~x62 && ~x18 && x17 && ~x7 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && ~x18 && ~x17 && x15 )
						nx_state = s1;
					else if( x69 && ~x62 && ~x18 && ~x17 && ~x15 && x1 && x2 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( x69 && ~x62 && ~x18 && ~x17 && ~x15 && x1 && ~x2 )
						nx_state = s1;
					else if( x69 && ~x62 && ~x18 && ~x17 && ~x15 && ~x1 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x69 && x70 && x64 && x11 && x43 && x9 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x70 && x64 && x11 && x43 && ~x9 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x70 && x64 && x11 && x43 && ~x9 && ~x34 && x1 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x69 && x70 && x64 && x11 && x43 && ~x9 && ~x34 && ~x1 && x38 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s801;
						end
					else if( ~x69 && x70 && x64 && x11 && x43 && ~x9 && ~x34 && ~x1 && ~x38 )
						nx_state = s444;
					else if( ~x69 && x70 && x64 && x11 && ~x43 && x44 && x10 && x35 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && x64 && x11 && ~x43 && x44 && x10 && ~x35 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x70 && x64 && x11 && ~x43 && x44 && ~x10 && x9 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x70 && x64 && x11 && ~x43 && x44 && ~x10 && ~x9 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x70 && x64 && x11 && ~x43 && x44 && ~x10 && ~x9 && ~x34 && x1 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x69 && x70 && x64 && x11 && ~x43 && x44 && ~x10 && ~x9 && ~x34 && ~x1 && x38 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s801;
						end
					else if( ~x69 && x70 && x64 && x11 && ~x43 && x44 && ~x10 && ~x9 && ~x34 && ~x1 && ~x38 )
						nx_state = s444;
					else if( ~x69 && x70 && x64 && x11 && ~x43 && ~x44 && x9 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x70 && x64 && x11 && ~x43 && ~x44 && ~x9 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x70 && x64 && x11 && ~x43 && ~x44 && ~x9 && ~x34 && x1 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x69 && x70 && x64 && x11 && ~x43 && ~x44 && ~x9 && ~x34 && ~x1 && x38 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s801;
						end
					else if( ~x69 && x70 && x64 && x11 && ~x43 && ~x44 && ~x9 && ~x34 && ~x1 && ~x38 )
						nx_state = s444;
					else if( ~x69 && x70 && x64 && ~x11 && x12 && x9 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x70 && x64 && ~x11 && x12 && ~x9 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x70 && x64 && ~x11 && x12 && ~x9 && ~x34 && x1 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x69 && x70 && x64 && ~x11 && x12 && ~x9 && ~x34 && ~x1 && x38 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s801;
						end
					else if( ~x69 && x70 && x64 && ~x11 && x12 && ~x9 && ~x34 && ~x1 && ~x38 )
						nx_state = s444;
					else if( ~x69 && x70 && x64 && ~x11 && ~x12 && x13 && x45 && x41 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x69 && x70 && x64 && ~x11 && ~x12 && x13 && x45 && ~x41 && x9 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x70 && x64 && ~x11 && ~x12 && x13 && x45 && ~x41 && ~x9 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x70 && x64 && ~x11 && ~x12 && x13 && x45 && ~x41 && ~x9 && ~x34 && x1 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x69 && x70 && x64 && ~x11 && ~x12 && x13 && x45 && ~x41 && ~x9 && ~x34 && ~x1 && x38 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s801;
						end
					else if( ~x69 && x70 && x64 && ~x11 && ~x12 && x13 && x45 && ~x41 && ~x9 && ~x34 && ~x1 && ~x38 )
						nx_state = s444;
					else if( ~x69 && x70 && x64 && ~x11 && ~x12 && x13 && ~x45 && x9 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x70 && x64 && ~x11 && ~x12 && x13 && ~x45 && ~x9 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x70 && x64 && ~x11 && ~x12 && x13 && ~x45 && ~x9 && ~x34 && x1 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x69 && x70 && x64 && ~x11 && ~x12 && x13 && ~x45 && ~x9 && ~x34 && ~x1 && x38 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s801;
						end
					else if( ~x69 && x70 && x64 && ~x11 && ~x12 && x13 && ~x45 && ~x9 && ~x34 && ~x1 && ~x38 )
						nx_state = s444;
					else if( ~x69 && x70 && x64 && ~x11 && ~x12 && ~x13 && x9 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x70 && x64 && ~x11 && ~x12 && ~x13 && ~x9 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x70 && x64 && ~x11 && ~x12 && ~x13 && ~x9 && ~x34 && x1 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x69 && x70 && x64 && ~x11 && ~x12 && ~x13 && ~x9 && ~x34 && ~x1 && x38 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s801;
						end
					else if( ~x69 && x70 && x64 && ~x11 && ~x12 && ~x13 && ~x9 && ~x34 && ~x1 && ~x38 )
						nx_state = s444;
					else if( ~x69 && x70 && ~x64 && x15 && x25 && x22 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x64 && x15 && x25 && ~x22 && x6 && x8 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && x70 && ~x64 && x15 && x25 && ~x22 && x6 && ~x8 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x64 && x15 && x25 && ~x22 && ~x6 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x69 && x70 && ~x64 && x15 && ~x25 && x29 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s190;
						end
					else if( ~x69 && x70 && ~x64 && x15 && ~x25 && ~x29 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x69 && x70 && ~x64 && ~x15 && x38 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x69 && x70 && ~x64 && ~x15 && ~x38 && x49 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && ~x64 && ~x15 && ~x38 && ~x49 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && ~x70 && x25 && x22 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x25 && ~x22 && x6 && x8 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && ~x70 && x25 && ~x22 && x6 && ~x8 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x25 && ~x22 && ~x6 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x69 && ~x70 && ~x25 && x29 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s190;
						end
					else if( ~x69 && ~x70 && ~x25 && ~x29 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else nx_state = s444;
				s445 : if( x15 && x16 && x5 && x1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s326;
						end
					else if( x15 && x16 && x5 && ~x1 && x2 && x3 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s455;
						end
					else if( x15 && x16 && x5 && ~x1 && x2 && x3 && ~x4 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x15 && x16 && x5 && ~x1 && x2 && ~x3 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x15 && x16 && x5 && ~x1 && ~x2 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x15 && x16 && ~x5 && x6 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x15 && x16 && ~x5 && ~x6 && x1 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( x15 && x16 && ~x5 && ~x6 && ~x1 && x2 && x3 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s455;
						end
					else if( x15 && x16 && ~x5 && ~x6 && ~x1 && x2 && x3 && ~x4 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( x15 && x16 && ~x5 && ~x6 && ~x1 && x2 && ~x3 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x15 && x16 && ~x5 && ~x6 && ~x1 && ~x2 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x15 && ~x16 && x6 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x15 && ~x16 && ~x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s446;
						end
					else if( ~x15 && x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( ~x15 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else nx_state = s445;
				s446 : if( x15 && x16 && x64 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x15 && x16 && ~x64 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s540;
						end
					else if( x15 && ~x16 && x8 && x64 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s441;
						end
					else if( x15 && ~x16 && x8 && ~x64 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s1045;
						end
					else if( x15 && ~x16 && ~x8 && x9 && x64 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s441;
						end
					else if( x15 && ~x16 && ~x8 && x9 && ~x64 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s1045;
						end
					else if( x15 && ~x16 && ~x8 && ~x9 && x10 && x6 && x64 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x15 && ~x16 && ~x8 && ~x9 && x10 && x6 && ~x64 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s540;
						end
					else if( x15 && ~x16 && ~x8 && ~x9 && x10 && ~x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s446;
						end
					else if( x15 && ~x16 && ~x8 && ~x9 && ~x10 && x11 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( x15 && ~x16 && ~x8 && ~x9 && ~x10 && ~x11 )
						nx_state = s446;
					else if( ~x15 && x64 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x15 && ~x64 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s540;
						end
					else nx_state = s446;
				s447 : if( x62 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s449;
						end
					else if( ~x62 && x64 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s456;
						end
					else if( ~x62 && ~x64 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s670;
						end
					else nx_state = s447;
				s448 : if( x16 && x15 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x16 && ~x15 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s193;
						end
					else if( x16 && ~x15 && x4 && ~x5 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( x16 && ~x15 && ~x4 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s436;
						end
					else if( ~x16 && x15 )
						begin
							y10 = 1'b1;	
							nx_state = s193;
						end
					else if( ~x16 && ~x15 && x12 && x13 && x3 )
						begin
							y13 = 1'b1;	
							nx_state = s450;
						end
					else if( ~x16 && ~x15 && x12 && x13 && ~x3 && x14 )
						begin
							y13 = 1'b1;	
							nx_state = s450;
						end
					else if( ~x16 && ~x15 && x12 && x13 && ~x3 && ~x14 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s451;
						end
					else if( ~x16 && ~x15 && x12 && ~x13 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s195;
						end
					else if( ~x16 && ~x15 && ~x12 )
						begin
							y10 = 1'b1;	
							nx_state = s193;
						end
					else nx_state = s448;
				s449 : if( x62 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s1105;
						end
					else if( ~x62 && x64 && x40 && x29 && x50 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1106;
						end
					else if( ~x62 && x64 && x40 && x29 && ~x50 )
						nx_state = s449;
					else if( ~x62 && x64 && x40 && ~x29 && x41 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x62 && x64 && x40 && ~x29 && ~x41 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x62 && x64 && ~x40 && x11 && x6 && x9 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x62 && x64 && ~x40 && x11 && x6 && ~x9 )
						begin
							y3 = 1'b1;	y13 = 1'b1;	y18 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s639;
						end
					else if( ~x62 && x64 && ~x40 && x11 && ~x6 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s510;
						end
					else if( ~x62 && x64 && ~x40 && ~x11 && x8 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x62 && x64 && ~x40 && ~x11 && ~x8 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else if( ~x62 && ~x64 && x44 && x29 && x50 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s1107;
						end
					else if( ~x62 && ~x64 && x44 && x29 && ~x50 )
						nx_state = s449;
					else if( ~x62 && ~x64 && x44 && ~x29 && x45 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x62 && ~x64 && x44 && ~x29 && ~x45 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x62 && ~x64 && ~x44 && x11 && x6 && x9 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x62 && ~x64 && ~x44 && x11 && x6 && ~x9 )
						begin
							y3 = 1'b1;	y13 = 1'b1;	y22 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s640;
						end
					else if( ~x62 && ~x64 && ~x44 && x11 && ~x6 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s510;
						end
					else if( ~x62 && ~x64 && ~x44 && ~x11 && x8 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x62 && ~x64 && ~x44 && ~x11 && ~x8 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else nx_state = s449;
				s450 : if( x62 && x69 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s1108;
						end
					else if( x62 && x69 && ~x17 )
						begin
							y1 = 1'b1;	y12 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s647;
						end
					else if( x62 && ~x69 && x15 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s194;
						end
					else if( x62 && ~x69 && ~x15 && x16 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x62 && ~x69 && ~x15 && ~x16 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s627;
						end
					else if( ~x62 && x69 && x64 )
						begin
							y29 = 1'b1;	
							nx_state = s1109;
						end
					else if( ~x62 && x69 && ~x64 )
						begin
							y22 = 1'b1;	
							nx_state = s683;
						end
					else if( ~x62 && ~x69 && x63 && x55 && x33 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s908;
						end
					else if( ~x62 && ~x69 && x63 && x55 && ~x33 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x62 && ~x69 && x63 && x55 && ~x33 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x62 && ~x69 && x63 && ~x55 && x50 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s910;
						end
					else if( ~x62 && ~x69 && x63 && ~x55 && ~x50 )
						nx_state = s450;
					else if( ~x62 && ~x69 && ~x63 && x64 && x40 && x33 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( ~x62 && ~x69 && ~x63 && x64 && x40 && ~x33 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x62 && ~x69 && ~x63 && x64 && x40 && ~x33 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x62 && ~x69 && ~x63 && x64 && ~x40 && x50 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s910;
						end
					else if( ~x62 && ~x69 && ~x63 && x64 && ~x40 && ~x50 )
						nx_state = s450;
					else if( ~x62 && ~x69 && ~x63 && ~x64 && x44 && x33 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( ~x62 && ~x69 && ~x63 && ~x64 && x44 && ~x33 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x62 && ~x69 && ~x63 && ~x64 && x44 && ~x33 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x62 && ~x69 && ~x63 && ~x64 && ~x44 && x50 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s910;
						end
					else if( ~x62 && ~x69 && ~x63 && ~x64 && ~x44 && ~x50 )
						nx_state = s450;
					else nx_state = s450;
				s451 : if( x16 && x15 && x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s927;
						end
					else if( x16 && x15 && ~x5 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s928;
						end
					else if( x16 && ~x15 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s448;
						end
					else if( ~x16 && x15 && x12 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s928;
						end
					else if( ~x16 && x15 && ~x12 )
						nx_state = s451;
					else if( ~x16 && ~x15 && x13 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x16 && ~x15 && ~x13 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s928;
						end
					else nx_state = s451;
				s452 : if( 1'b1 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y29 = 1'b1;	
							nx_state = s288;
						end
					else nx_state = s452;
				s453 : if( x15 && x16 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x15 && ~x16 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x15 && x47 && x4 && x5 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x15 && x47 && x4 && ~x5 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s441;
						end
					else if( ~x15 && x47 && ~x4 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x15 && ~x47 && x43 && x44 && x34 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x15 && ~x47 && x43 && x44 && ~x34 && x14 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x15 && ~x47 && x43 && x44 && ~x34 && ~x14 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s322;
						end
					else if( ~x15 && ~x47 && x43 && ~x44 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x15 && ~x47 && ~x43 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else nx_state = s453;
				s454 : if( x69 && x62 && x13 && x8 && x1 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && x62 && x13 && x8 && ~x1 && x14 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && x62 && x13 && x8 && ~x1 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && x62 && x13 && ~x8 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( x69 && x62 && ~x13 && x10 )
						nx_state = s1;
					else if( x69 && x62 && ~x13 && ~x10 && x6 && x7 && x5 && x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s540;
						end
					else if( x69 && x62 && ~x13 && ~x10 && x6 && x7 && x5 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x69 && x62 && ~x13 && ~x10 && x6 && x7 && x5 && ~x3 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && x62 && ~x13 && ~x10 && x6 && x7 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && x62 && ~x13 && ~x10 && x6 && ~x7 && x8 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( x69 && x62 && ~x13 && ~x10 && x6 && ~x7 && ~x8 && x5 && x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s540;
						end
					else if( x69 && x62 && ~x13 && ~x10 && x6 && ~x7 && ~x8 && x5 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x69 && x62 && ~x13 && ~x10 && x6 && ~x7 && ~x8 && x5 && ~x3 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && x62 && ~x13 && ~x10 && x6 && ~x7 && ~x8 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && x62 && ~x13 && ~x10 && ~x6 && x16 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( x69 && x62 && ~x13 && ~x10 && ~x6 && ~x16 )
						nx_state = s1;
					else if( x69 && ~x62 && x17 && x18 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x5 && x6 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x5 && ~x6 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && x17 && ~x18 && x9 && x10 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && ~x62 && x17 && ~x18 && x9 && ~x10 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && ~x62 && x17 && ~x18 && ~x9 && x6 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( x69 && ~x62 && x17 && ~x18 && ~x9 && ~x6 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && ~x62 && ~x17 && x18 )
						nx_state = s1;
					else if( x69 && ~x62 && ~x17 && ~x18 && x6 && x7 && x2 && x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 && x6 && x7 && x2 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 && x6 && x7 && x2 && ~x3 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 && x6 && x7 && ~x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 && x6 && ~x7 && x8 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 && x6 && ~x7 && ~x8 && x2 && x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 && x6 && ~x7 && ~x8 && x2 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 && x6 && ~x7 && ~x8 && x2 && ~x3 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 && x6 && ~x7 && ~x8 && ~x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 && ~x6 && x2 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 && ~x6 && ~x2 )
						nx_state = s1;
					else if( ~x69 && x70 && x63 && x64 && x42 && x43 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && x63 && x64 && x42 && ~x43 && x44 && x10 && x36 && x6 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x69 && x70 && x63 && x64 && x42 && ~x43 && x44 && x10 && x36 && ~x6 && x7 && x15 && x47 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x69 && x70 && x63 && x64 && x42 && ~x43 && x44 && x10 && x36 && ~x6 && x7 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && x63 && x64 && x42 && ~x43 && x44 && x10 && x36 && ~x6 && x7 && x15 && ~x47 && ~x1 )
						nx_state = s454;
					else if( ~x69 && x70 && x63 && x64 && x42 && ~x43 && x44 && x10 && x36 && ~x6 && x7 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && x63 && x64 && x42 && ~x43 && x44 && x10 && x36 && ~x6 && x7 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x69 && x70 && x63 && x64 && x42 && ~x43 && x44 && x10 && x36 && ~x6 && x7 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x69 && x70 && x63 && x64 && x42 && ~x43 && x44 && x10 && x36 && ~x6 && ~x7 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s902;
						end
					else if( ~x69 && x70 && x63 && x64 && x42 && ~x43 && x44 && x10 && ~x36 && x35 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && x63 && x64 && x42 && ~x43 && x44 && x10 && ~x36 && ~x35 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x70 && x63 && x64 && x42 && ~x43 && x44 && ~x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && x63 && x64 && x42 && ~x43 && ~x44 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && x63 && x64 && ~x42 && x12 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && x63 && x64 && ~x42 && ~x12 && x13 && x14 && x41 && x4 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x69 && x70 && x63 && x64 && ~x42 && ~x12 && x13 && x14 && x41 && ~x4 )
						nx_state = s454;
					else if( ~x69 && x70 && x63 && x64 && ~x42 && ~x12 && x13 && x14 && ~x41 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && x63 && x64 && ~x42 && ~x12 && x13 && ~x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && x63 && x64 && ~x42 && ~x12 && ~x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x69 && x70 && x63 && ~x64 && x15 && x16 && x19 && x33 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && x70 && x63 && ~x64 && x15 && x16 && x19 && ~x33 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && x70 && x63 && ~x64 && x15 && x16 && x19 && ~x33 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && x70 && x63 && ~x64 && x15 && x16 && ~x19 && x30 && x26 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x69 && x70 && x63 && ~x64 && x15 && x16 && ~x19 && x30 && x26 && ~x1 )
						nx_state = s454;
					else if( ~x69 && x70 && x63 && ~x64 && x15 && x16 && ~x19 && x30 && ~x26 && x3 )
						nx_state = s454;
					else if( ~x69 && x70 && x63 && ~x64 && x15 && x16 && ~x19 && x30 && ~x26 && ~x3 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x69 && x70 && x63 && ~x64 && x15 && x16 && ~x19 && x30 && ~x26 && ~x3 && ~x1 )
						nx_state = s454;
					else if( ~x69 && x70 && x63 && ~x64 && x15 && x16 && ~x19 && ~x30 )
						nx_state = s454;
					else if( ~x69 && x70 && x63 && ~x64 && x15 && ~x16 )
						nx_state = s1;
					else if( ~x69 && x70 && x63 && ~x64 && ~x15 && x28 && x41 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x69 && x70 && x63 && ~x64 && ~x15 && x28 && ~x41 )
						nx_state = s454;
					else if( ~x69 && x70 && x63 && ~x64 && ~x15 && ~x28 && x27 && x8 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x69 && x70 && x63 && ~x64 && ~x15 && ~x28 && x27 && ~x8 && x37 )
						nx_state = s1;
					else if( ~x69 && x70 && x63 && ~x64 && ~x15 && ~x28 && x27 && ~x8 && ~x37 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && x70 && x63 && ~x64 && ~x15 && ~x28 && ~x27 && x49 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x70 && x63 && ~x64 && ~x15 && ~x28 && ~x27 && ~x49 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x70 && ~x63 && x17 && x18 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( ~x69 && x70 && ~x63 && x17 && x18 && ~x5 && x6 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x70 && ~x63 && x17 && x18 && ~x5 && ~x6 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x70 && ~x63 && x17 && ~x18 && x9 && x10 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( ~x69 && x70 && ~x63 && x17 && ~x18 && x9 && ~x10 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x70 && ~x63 && x17 && ~x18 && ~x9 && x6 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( ~x69 && x70 && ~x63 && x17 && ~x18 && ~x9 && ~x6 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && x18 && x15 && x16 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && x18 && x15 && x16 && ~x5 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && x18 && x15 && x16 && ~x5 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && x18 && x15 && ~x16 && x1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && x18 && x15 && ~x16 && ~x1 )
						nx_state = s454;
					else if( ~x69 && x70 && ~x63 && ~x17 && x18 && ~x15 && x16 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && x18 && ~x15 && ~x16 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && x18 && ~x15 && ~x16 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && ~x18 && x6 && x7 && x39 && x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && ~x18 && x6 && x7 && x39 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && ~x18 && x6 && x7 && x39 && ~x3 && ~x4 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s543;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && ~x18 && x6 && x7 && ~x39 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && ~x18 && x6 && ~x7 && x8 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && ~x18 && x6 && ~x7 && ~x8 && x39 && x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && ~x18 && x6 && ~x7 && ~x8 && x39 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && ~x18 && x6 && ~x7 && ~x8 && x39 && ~x3 && ~x4 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s543;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && ~x18 && x6 && ~x7 && ~x8 && ~x39 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && ~x18 && ~x6 && x32 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && ~x18 && ~x6 && ~x32 && x15 && x16 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && ~x18 && ~x6 && ~x32 && x15 && x16 && ~x5 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && ~x18 && ~x6 && ~x32 && x15 && ~x16 && x1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && ~x18 && ~x6 && ~x32 && x15 && ~x16 && ~x1 )
						nx_state = s454;
					else if( ~x69 && x70 && ~x63 && ~x17 && ~x18 && ~x6 && ~x32 && ~x15 && x16 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && ~x18 && ~x6 && ~x32 && ~x15 && ~x16 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x69 && x70 && ~x63 && ~x17 && ~x18 && ~x6 && ~x32 && ~x15 && ~x16 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x70 && x16 && x19 && x20 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && ~x70 && x16 && x19 && ~x20 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && ~x70 && x16 && x19 && ~x20 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && ~x70 && x16 && ~x19 && x30 && x26 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x69 && ~x70 && x16 && ~x19 && x30 && x26 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && ~x70 && x16 && ~x19 && x30 && ~x26 && x3 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && ~x70 && x16 && ~x19 && x30 && ~x26 && ~x3 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x69 && ~x70 && x16 && ~x19 && x30 && ~x26 && ~x3 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && ~x70 && x16 && ~x19 && ~x30 && x8 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && ~x70 && x16 && ~x19 && ~x30 && ~x8 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x16 )
						nx_state = s1;
					else nx_state = s454;
				s455 : if( x16 && x15 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x16 && ~x15 && x4 && x64 && x5 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( x16 && ~x15 && x4 && x64 && ~x5 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s441;
						end
					else if( x16 && ~x15 && x4 && ~x64 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( x16 && ~x15 && x4 && ~x64 && ~x5 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s1045;
						end
					else if( x16 && ~x15 && ~x4 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x16 && x12 && x15 && x64 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x16 && x12 && x15 && ~x64 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x16 && x12 && ~x15 && x13 && x3 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x16 && x12 && ~x15 && x13 && ~x3 && x14 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x16 && x12 && ~x15 && x13 && ~x3 && ~x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s326;
						end
					else if( ~x16 && x12 && ~x15 && ~x13 && x64 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x16 && x12 && ~x15 && ~x13 && ~x64 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x16 && ~x12 && x64 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x16 && ~x12 && ~x64 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else nx_state = s455;
				s456 : if( x69 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s689;
						end
					else if( ~x69 && x63 && x55 && x46 && x3 && x23 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( ~x69 && x63 && x55 && x46 && x3 && ~x23 )
						nx_state = s456;
					else if( ~x69 && x63 && x55 && x46 && ~x3 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && x63 && x55 && ~x46 && x2 && x23 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( ~x69 && x63 && x55 && ~x46 && x2 && ~x23 )
						nx_state = s456;
					else if( ~x69 && x63 && x55 && ~x46 && ~x2 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && x63 && ~x55 && x10 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && x63 && ~x55 && ~x10 && x11 && x5 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s818;
						end
					else if( ~x69 && x63 && ~x55 && ~x10 && x11 && ~x5 && x37 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( ~x69 && x63 && ~x55 && ~x10 && x11 && ~x5 && ~x37 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && x63 && ~x55 && ~x10 && ~x11 && x1 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && x63 && ~x55 && ~x10 && ~x11 && ~x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( ~x69 && ~x63 && x64 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s498;
						end
					else if( ~x69 && ~x63 && ~x64 )
						begin
							y19 = 1'b1;	y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s1032;
						end
					else nx_state = s456;
				s457 : if( x3 && x1 && x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s46;
						end
					else if( x3 && x1 && ~x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s557;
						end
					else if( x3 && ~x1 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	
							nx_state = s594;
						end
					else if( ~x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else nx_state = s457;
				s458 : if( x65 && x67 && x22 && x15 && x8 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && x67 && x22 && x15 && ~x8 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x65 && x67 && x22 && ~x15 && x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s126;
						end
					else if( x65 && x67 && x22 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( x65 && x67 && ~x22 && x15 && x8 && x23 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && x67 && ~x22 && x15 && x8 && ~x23 )
						begin
							y11 = 1'b1;	
							nx_state = s91;
						end
					else if( x65 && x67 && ~x22 && x15 && ~x8 && x23 && x6 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s591;
						end
					else if( x65 && x67 && ~x22 && x15 && ~x8 && x23 && ~x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && x67 && ~x22 && x15 && ~x8 && ~x23 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s591;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && x8 && x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && x8 && ~x7 && x9 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && x8 && ~x7 && ~x9 && x18 && x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && x8 && ~x7 && ~x9 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && x8 && ~x7 && ~x9 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && x8 && ~x7 && ~x9 && ~x18 )
						nx_state = s1;
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && ~x8 && x7 && x11 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && ~x8 && x7 && ~x11 && x18 && x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && ~x8 && x7 && ~x11 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && ~x8 && x7 && ~x11 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && ~x8 && x7 && ~x11 && ~x18 )
						nx_state = s1;
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && ~x8 && ~x7 && x10 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && ~x8 && ~x7 && ~x10 && x18 && x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && ~x8 && ~x7 && ~x10 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && ~x8 && ~x7 && ~x10 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && ~x8 && ~x7 && ~x10 && ~x18 )
						nx_state = s1;
					else if( x65 && x67 && ~x22 && ~x15 && x16 && ~x23 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( x65 && x67 && ~x22 && ~x15 && ~x16 && x23 && x6 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x65 && x67 && ~x22 && ~x15 && ~x16 && x23 && ~x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && x67 && ~x22 && ~x15 && ~x16 && ~x23 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x65 && ~x67 && x61 && x60 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( x65 && ~x67 && x61 && ~x60 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x65 && ~x67 && ~x61 && x60 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x65 && ~x67 && ~x61 && ~x60 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x65 && x22 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x22 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else nx_state = s458;
				s459 : if( 1'b1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s46;
						end
					else nx_state = s459;
				s460 : if( x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y8 = 1'b1;	
							nx_state = s2;
						end
					else if( ~x5 && x2 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s459;
						end
					else if( ~x5 && x2 && ~x1 )
						begin
							y3 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							nx_state = s460;
						end
					else if( ~x5 && ~x2 && x1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s461;
						end
					else if( ~x5 && ~x2 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y8 = 1'b1;	
							nx_state = s2;
						end
					else nx_state = s460;
				s461 : if( x70 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x70 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s805;
						end
					else nx_state = s461;
				s462 : if( x62 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x62 && x30 )
						begin
							y33 = 1'b1;	
							nx_state = s589;
						end
					else if( ~x62 && ~x30 && x31 )
						begin
							y47 = 1'b1;	y56 = 1'b1;	y61 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s1110;
						end
					else if( ~x62 && ~x30 && ~x31 )
						begin
							y47 = 1'b1;	y52 = 1'b1;	y61 = 1'b1;	
							y66 = 1'b1;	
							nx_state = s54;
						end
					else nx_state = s462;
				s463 : if( x19 && x18 )
						begin
							y2 = 1'b1;	
							nx_state = s1111;
						end
					else if( x19 && ~x18 )
						begin
							y2 = 1'b1;	
							nx_state = s1112;
						end
					else if( ~x19 )
						begin
							y2 = 1'b1;	
							nx_state = s768;
						end
					else nx_state = s463;
				s464 : if( x16 && x15 && x10 && x12 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x16 && x15 && x10 && ~x12 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x16 && x15 && ~x10 && x11 && x12 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s358;
						end
					else if( x16 && x15 && ~x10 && x11 && ~x12 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s600;
						end
					else if( x16 && x15 && ~x10 && ~x11 && x12 && x13 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s426;
						end
					else if( x16 && x15 && ~x10 && ~x11 && x12 && ~x13 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x16 && x15 && ~x10 && ~x11 && x12 && ~x13 && x17 && ~x14 )
						nx_state = s1;
					else if( x16 && x15 && ~x10 && ~x11 && x12 && ~x13 && ~x17 )
						nx_state = s1;
					else if( x16 && x15 && ~x10 && ~x11 && ~x12 && x14 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s426;
						end
					else if( x16 && x15 && ~x10 && ~x11 && ~x12 && ~x14 && x17 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x16 && x15 && ~x10 && ~x11 && ~x12 && ~x14 && x17 && ~x13 )
						nx_state = s1;
					else if( x16 && x15 && ~x10 && ~x11 && ~x12 && ~x14 && ~x17 )
						nx_state = s1;
					else if( x16 && ~x15 && x12 && x10 && x8 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x16 && ~x15 && x12 && x10 && x8 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x16 && ~x15 && x12 && x10 && x8 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x16 && ~x15 && x12 && x10 && x8 && ~x17 )
						nx_state = s1;
					else if( x16 && ~x15 && x12 && x10 && ~x8 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( x16 && ~x15 && x12 && x10 && ~x8 && ~x5 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s731;
						end
					else if( x16 && ~x15 && x12 && x10 && ~x8 && ~x5 && ~x2 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s603;
						end
					else if( x16 && ~x15 && x12 && ~x10 && x11 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( x16 && ~x15 && x12 && ~x10 && x11 && ~x5 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s731;
						end
					else if( x16 && ~x15 && x12 && ~x10 && x11 && ~x5 && ~x2 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s603;
						end
					else if( x16 && ~x15 && x12 && ~x10 && ~x11 && x7 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( x16 && ~x15 && x12 && ~x10 && ~x11 && x7 && ~x5 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s731;
						end
					else if( x16 && ~x15 && x12 && ~x10 && ~x11 && x7 && ~x5 && ~x2 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s603;
						end
					else if( x16 && ~x15 && x12 && ~x10 && ~x11 && ~x7 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x16 && ~x15 && x12 && ~x10 && ~x11 && ~x7 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x16 && ~x15 && x12 && ~x10 && ~x11 && ~x7 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x16 && ~x15 && x12 && ~x10 && ~x11 && ~x7 && ~x17 )
						nx_state = s1;
					else if( x16 && ~x15 && ~x12 && x10 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( x16 && ~x15 && ~x12 && x10 && ~x5 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s778;
						end
					else if( x16 && ~x15 && ~x12 && x10 && ~x5 && ~x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s731;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && x11 && x9 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && x11 && x9 && ~x5 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s731;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && x11 && x9 && ~x5 && ~x2 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s603;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x16 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && ~x17 )
						nx_state = s1;
					else if( x16 && ~x15 && ~x12 && ~x10 && ~x11 && x8 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && ~x11 && x8 && ~x5 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s731;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && ~x11 && x8 && ~x5 && ~x2 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s603;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x16 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && ~x17 )
						nx_state = s1;
					else if( ~x16 && x15 && x10 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x16 && x15 && x10 && ~x5 && x11 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s731;
						end
					else if( ~x16 && x15 && x10 && ~x5 && x11 && ~x2 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x16 && x15 && x10 && ~x5 && ~x11 && x12 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s731;
						end
					else if( ~x16 && x15 && x10 && ~x5 && ~x11 && x12 && ~x2 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s601;
						end
					else if( ~x16 && x15 && x10 && ~x5 && ~x11 && ~x12 && x2 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s606;
						end
					else if( ~x16 && x15 && x10 && ~x5 && ~x11 && ~x12 && ~x2 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y13 = 1'b1;	
							nx_state = s600;
						end
					else if( ~x16 && x15 && ~x10 && x11 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x16 && x15 && ~x10 && ~x11 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x16 && x15 && ~x10 && ~x11 && ~x5 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s731;
						end
					else if( ~x16 && x15 && ~x10 && ~x11 && ~x5 && ~x2 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( ~x16 && x15 && ~x10 && ~x11 && ~x5 && ~x2 && ~x12 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s556;
						end
					else if( ~x16 && ~x15 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x16 && ~x15 && ~x5 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s731;
						end
					else if( ~x16 && ~x15 && ~x5 && ~x2 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s209;
						end
					else nx_state = s464;
				s465 : if( x21 && x18 && x4 && x15 && x17 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x21 && x18 && x4 && x15 && ~x17 )
						begin
							y12 = 1'b1;	
							nx_state = s245;
						end
					else if( x21 && x18 && x4 && ~x15 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s797;
						end
					else if( x21 && x18 && ~x4 )
						begin
							y12 = 1'b1;	
							nx_state = s245;
						end
					else if( x21 && ~x18 && x19 && x15 && x4 && x17 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x21 && ~x18 && x19 && x15 && x4 && ~x17 )
						begin
							y12 = 1'b1;	
							nx_state = s245;
						end
					else if( x21 && ~x18 && x19 && x15 && ~x4 )
						begin
							y12 = 1'b1;	
							nx_state = s245;
						end
					else if( x21 && ~x18 && x19 && ~x15 && x16 && x14 )
						begin
							y12 = 1'b1;	
							nx_state = s245;
						end
					else if( x21 && ~x18 && x19 && ~x15 && x16 && ~x14 && x17 )
						begin
							y12 = 1'b1;	
							nx_state = s245;
						end
					else if( x21 && ~x18 && x19 && ~x15 && x16 && ~x14 && ~x17 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && ~x18 && x19 && ~x15 && x16 && ~x14 && ~x17 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && ~x18 && x19 && ~x15 && x16 && ~x14 && ~x17 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x18 && x19 && ~x15 && x16 && ~x14 && ~x17 && ~x8 )
						nx_state = s1;
					else if( x21 && ~x18 && x19 && ~x15 && ~x16 && x17 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s245;
						end
					else if( x21 && ~x18 && x19 && ~x15 && ~x16 && x17 && ~x12 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && ~x18 && x19 && ~x15 && ~x16 && x17 && ~x12 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && ~x18 && x19 && ~x15 && ~x16 && x17 && ~x12 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x18 && x19 && ~x15 && ~x16 && x17 && ~x12 && ~x8 )
						nx_state = s1;
					else if( x21 && ~x18 && x19 && ~x15 && ~x16 && ~x17 && x13 )
						begin
							y12 = 1'b1;	
							nx_state = s245;
						end
					else if( x21 && ~x18 && x19 && ~x15 && ~x16 && ~x17 && ~x13 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && ~x18 && x19 && ~x15 && ~x16 && ~x17 && ~x13 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && ~x18 && x19 && ~x15 && ~x16 && ~x17 && ~x13 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x18 && x19 && ~x15 && ~x16 && ~x17 && ~x13 && ~x8 )
						nx_state = s1;
					else if( x21 && ~x18 && ~x19 && x4 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s115;
						end
					else if( x21 && ~x18 && ~x19 && ~x4 )
						begin
							y12 = 1'b1;	
							nx_state = s245;
						end
					else if( ~x21 && x23 && x22 && x6 )
						begin
							y12 = 1'b1;	
							nx_state = s245;
						end
					else if( ~x21 && x23 && x22 && ~x6 && x7 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && x23 && x22 && ~x6 && x7 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && x23 && x22 && ~x6 && x7 && ~x18 && x19 && x15 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s666;
						end
					else if( ~x21 && x23 && x22 && ~x6 && x7 && ~x18 && x19 && ~x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( ~x21 && x23 && x22 && ~x6 && x7 && ~x18 && ~x19 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x21 && x23 && x22 && ~x6 && ~x7 )
						begin
							y3 = 1'b1;	y12 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s113;
						end
					else if( ~x21 && x23 && ~x22 )
						begin
							y12 = 1'b1;	y19 = 1'b1;	
							nx_state = s794;
						end
					else if( ~x21 && ~x23 && x22 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s301;
						end
					else if( ~x21 && ~x23 && ~x22 && x6 )
						begin
							y12 = 1'b1;	
							nx_state = s245;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x6 && x7 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x6 && x7 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x6 && x7 && ~x18 && x19 && x15 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s666;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x6 && x7 && ~x18 && x19 && ~x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x6 && x7 && ~x18 && ~x19 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x6 && ~x7 )
						begin
							y3 = 1'b1;	y12 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s113;
						end
					else nx_state = s465;
				s466 : if( 1'b1 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							nx_state = s1113;
						end
					else nx_state = s466;
				s467 : if( x21 && x20 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x21 && ~x20 )
						begin
							y15 = 1'b1;	
							nx_state = s1114;
						end
					else if( ~x21 && x20 )
						begin
							y15 = 1'b1;	
							nx_state = s1115;
						end
					else if( ~x21 && ~x20 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else nx_state = s467;
				s468 : if( 1'b1 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else nx_state = s468;
				s469 : if( x62 )
						begin
							y29 = 1'b1;	
							nx_state = s771;
						end
					else if( ~x62 && x20 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && ~x20 && x9 )
						begin
							y15 = 1'b1;	
							nx_state = s1116;
						end
					else if( ~x62 && ~x20 && ~x9 )
						begin
							y14 = 1'b1;	
							nx_state = s366;
						end
					else nx_state = s469;
				s470 : if( x33 && x32 )
						nx_state = s1;
					else if( x33 && ~x32 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s968;
						end
					else if( ~x33 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s968;
						end
					else nx_state = s470;
				s471 : if( 1'b1 )
						begin
							y3 = 1'b1;	y53 = 1'b1;	
							nx_state = s1117;
						end
					else nx_state = s471;
				s472 : if( x13 && x10 && x12 && x11 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s27;
						end
					else if( x13 && x10 && x12 && ~x11 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x13 && x10 && x12 && ~x11 && ~x3 && x6 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s29;
						end
					else if( x13 && x10 && x12 && ~x11 && ~x3 && ~x6 )
						nx_state = s472;
					else if( x13 && x10 && ~x12 && x11 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x13 && x10 && ~x12 && x11 && ~x3 && x6 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s29;
						end
					else if( x13 && x10 && ~x12 && x11 && ~x3 && ~x6 )
						nx_state = s472;
					else if( x13 && x10 && ~x12 && ~x11 && x14 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x13 && x10 && ~x12 && ~x11 && x14 && ~x3 && x6 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s29;
						end
					else if( x13 && x10 && ~x12 && ~x11 && x14 && ~x3 && ~x6 )
						nx_state = s472;
					else if( x13 && x10 && ~x12 && ~x11 && ~x14 && x1 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s476;
						end
					else if( x13 && x10 && ~x12 && ~x11 && ~x14 && ~x1 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x13 && ~x10 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x13 && ~x10 && ~x3 && x6 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s29;
						end
					else if( x13 && ~x10 && ~x3 && ~x6 )
						nx_state = s472;
					else if( ~x13 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( ~x13 && ~x3 && x6 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x13 && ~x3 && ~x6 )
						nx_state = s472;
					else nx_state = s472;
				s473 : if( x2 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	
							nx_state = s474;
						end
					else if( ~x2 )
						nx_state = s473;
					else nx_state = s473;
				s474 : if( x12 && x11 && x10 && x13 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x12 && x11 && x10 && x13 && ~x8 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x12 && x11 && x10 && x13 && ~x8 && ~x1 )
						nx_state = s474;
					else if( x12 && x11 && x10 && ~x13 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s27;
						end
					else if( x12 && x11 && ~x10 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x12 && x11 && ~x10 && ~x8 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x12 && x11 && ~x10 && ~x8 && ~x1 )
						nx_state = s474;
					else if( x12 && ~x11 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x12 && ~x11 && ~x8 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x12 && ~x11 && ~x8 && ~x1 )
						nx_state = s474;
					else if( ~x12 && x11 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x12 && x11 && ~x8 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x12 && x11 && ~x8 && ~x1 )
						nx_state = s474;
					else if( ~x12 && ~x11 && x14 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x12 && ~x11 && x14 && ~x8 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x12 && ~x11 && x14 && ~x8 && ~x1 )
						nx_state = s474;
					else if( ~x12 && ~x11 && ~x14 && x13 && x10 && x9 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x12 && ~x11 && ~x14 && x13 && x10 && ~x9 && x7 )
						nx_state = s1;
					else if( ~x12 && ~x11 && ~x14 && x13 && x10 && ~x9 && ~x7 )
						begin
							y15 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s475;
						end
					else if( ~x12 && ~x11 && ~x14 && x13 && ~x10 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x12 && ~x11 && ~x14 && x13 && ~x10 && ~x8 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x12 && ~x11 && ~x14 && x13 && ~x10 && ~x8 && ~x1 )
						nx_state = s474;
					else if( ~x12 && ~x11 && ~x14 && ~x13 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x12 && ~x11 && ~x14 && ~x13 && ~x8 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x12 && ~x11 && ~x14 && ~x13 && ~x8 && ~x1 )
						nx_state = s474;
					else nx_state = s474;
				s475 : if( x11 && x12 && x4 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s31;
						end
					else if( x11 && x12 && ~x4 )
						nx_state = s475;
					else if( x11 && ~x12 && x13 )
						nx_state = s1;
					else if( x11 && ~x12 && ~x13 && x4 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s31;
						end
					else if( x11 && ~x12 && ~x13 && ~x4 )
						nx_state = s475;
					else if( ~x11 && x14 && x4 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s31;
						end
					else if( ~x11 && x14 && ~x4 )
						nx_state = s475;
					else if( ~x11 && ~x14 && x12 && x4 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s31;
						end
					else if( ~x11 && ~x14 && x12 && ~x4 )
						nx_state = s475;
					else if( ~x11 && ~x14 && ~x12 && x13 )
						nx_state = s1;
					else if( ~x11 && ~x14 && ~x12 && ~x13 && x4 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s31;
						end
					else if( ~x11 && ~x14 && ~x12 && ~x13 && ~x4 )
						nx_state = s475;
					else nx_state = s475;
				s476 : if( x70 && x10 && x13 && x11 && x12 && x3 && x6 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s24;
						end
					else if( x70 && x10 && x13 && x11 && x12 && x3 && ~x6 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x70 && x10 && x13 && x11 && x12 && ~x3 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x70 && x10 && x13 && x11 && ~x12 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x70 && x10 && x13 && ~x11 && x12 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x70 && x10 && x13 && ~x11 && x12 && ~x3 && x1 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x70 && x10 && x13 && ~x11 && x12 && ~x3 && ~x1 && x7 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	
							nx_state = s474;
						end
					else if( x70 && x10 && x13 && ~x11 && x12 && ~x3 && ~x1 && ~x7 )
						nx_state = s476;
					else if( x70 && x10 && x13 && ~x11 && ~x12 && x14 && x5 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y13 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s29;
						end
					else if( x70 && x10 && x13 && ~x11 && ~x12 && x14 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x70 && x10 && x13 && ~x11 && ~x12 && ~x14 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s28;
						end
					else if( x70 && x10 && ~x13 && x12 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x70 && x10 && ~x13 && x12 && ~x3 && x1 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x70 && x10 && ~x13 && x12 && ~x3 && ~x1 && x7 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	
							nx_state = s474;
						end
					else if( x70 && x10 && ~x13 && x12 && ~x3 && ~x1 && ~x7 )
						nx_state = s476;
					else if( x70 && x10 && ~x13 && ~x12 && x14 && x5 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s28;
						end
					else if( x70 && x10 && ~x13 && ~x12 && x14 && ~x5 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x70 && x10 && ~x13 && ~x12 && ~x14 && x1 )
						begin
							y5 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s26;
						end
					else if( x70 && x10 && ~x13 && ~x12 && ~x14 && ~x1 && x3 )
						nx_state = s1;
					else if( x70 && x10 && ~x13 && ~x12 && ~x14 && ~x1 && ~x3 )
						begin
							y14 = 1'b1;	y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s25;
						end
					else if( x70 && ~x10 && x3 )
						begin
							y22 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s32;
						end
					else if( x70 && ~x10 && ~x3 && x1 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x70 && ~x10 && ~x3 && ~x1 && x7 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	
							nx_state = s474;
						end
					else if( x70 && ~x10 && ~x3 && ~x1 && ~x7 )
						nx_state = s476;
					else if( ~x70 && x21 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( ~x70 && x21 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( ~x70 && x21 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x8 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x22 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s724;
						end
					else if( ~x70 && ~x21 && x22 && ~x12 && x8 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && x22 && ~x12 && x8 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && x22 && ~x12 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x22 && ~x12 && ~x8 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 && x12 && x23 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s666;
						end
					else if( ~x70 && ~x21 && ~x22 && x12 && ~x23 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x12 && x23 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x12 && x23 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x12 && x23 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 && ~x12 && x23 && ~x9 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 && ~x12 && ~x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x12 && ~x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x12 && ~x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 && ~x12 && ~x23 && ~x8 )
						nx_state = s1;
					else nx_state = s476;
				s477 : if( x69 && x62 && x1 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s636;
						end
					else if( x69 && x62 && ~x1 && x4 && x5 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s636;
						end
					else if( x69 && x62 && ~x1 && x4 && ~x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s60;
						end
					else if( x69 && x62 && ~x1 && ~x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( x69 && ~x62 && x15 && x16 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s636;
						end
					else if( x69 && ~x62 && x15 && ~x16 && x3 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( x69 && ~x62 && x15 && ~x16 && x3 && ~x2 )
						nx_state = s477;
					else if( x69 && ~x62 && x15 && ~x16 && ~x3 && x4 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s60;
						end
					else if( x69 && ~x62 && x15 && ~x16 && ~x3 && x4 && ~x2 )
						nx_state = s477;
					else if( x69 && ~x62 && x15 && ~x16 && ~x3 && ~x4 && x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( x69 && ~x62 && x15 && ~x16 && ~x3 && ~x4 && ~x2 )
						nx_state = s477;
					else if( x69 && ~x62 && ~x15 && x1 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s636;
						end
					else if( x69 && ~x62 && ~x15 && ~x1 && x16 && x4 && x5 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s636;
						end
					else if( x69 && ~x62 && ~x15 && ~x1 && x16 && x4 && ~x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s60;
						end
					else if( x69 && ~x62 && ~x15 && ~x1 && x16 && ~x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( x69 && ~x62 && ~x15 && ~x1 && ~x16 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s636;
						end
					else if( ~x69 && x15 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s705;
						end
					else if( ~x69 && ~x15 && x3 && x64 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( ~x69 && ~x15 && x3 && x64 && ~x2 )
						nx_state = s477;
					else if( ~x69 && ~x15 && x3 && ~x64 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s700;
						end
					else if( ~x69 && ~x15 && x3 && ~x64 && ~x2 )
						nx_state = s477;
					else if( ~x69 && ~x15 && ~x3 && x4 && x64 && x2 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s997;
						end
					else if( ~x69 && ~x15 && ~x3 && x4 && x64 && ~x2 )
						nx_state = s477;
					else if( ~x69 && ~x15 && ~x3 && x4 && ~x64 && x2 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s999;
						end
					else if( ~x69 && ~x15 && ~x3 && x4 && ~x64 && ~x2 )
						nx_state = s477;
					else if( ~x69 && ~x15 && ~x3 && ~x4 && x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1000;
						end
					else if( ~x69 && ~x15 && ~x3 && ~x4 && ~x2 )
						nx_state = s477;
					else nx_state = s477;
				s478 : if( x69 && x62 && x5 && x2 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y22 = 1'b1;	
							nx_state = s61;
						end
					else if( x69 && x62 && x5 && ~x2 && x4 && x1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( x69 && x62 && x5 && ~x2 && x4 && ~x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( x69 && x62 && x5 && ~x2 && ~x4 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y22 = 1'b1;	
							nx_state = s61;
						end
					else if( x69 && x62 && ~x5 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y22 = 1'b1;	
							nx_state = s61;
						end
					else if( x69 && ~x62 && x16 && x15 && x5 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x62 && x16 && x15 && ~x5 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s627;
						end
					else if( x69 && ~x62 && x16 && ~x15 && x2 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y22 = 1'b1;	
							nx_state = s61;
						end
					else if( x69 && ~x62 && x16 && ~x15 && ~x2 && x4 && x5 && x1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( x69 && ~x62 && x16 && ~x15 && ~x2 && x4 && x5 && ~x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( x69 && ~x62 && x16 && ~x15 && ~x2 && x4 && ~x5 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y22 = 1'b1;	
							nx_state = s61;
						end
					else if( x69 && ~x62 && x16 && ~x15 && ~x2 && ~x4 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y22 = 1'b1;	
							nx_state = s61;
						end
					else if( x69 && ~x62 && ~x16 && x15 && x13 && x11 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s637;
						end
					else if( x69 && ~x62 && ~x16 && x15 && x13 && ~x11 && x6 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s60;
						end
					else if( x69 && ~x62 && ~x16 && x15 && x13 && ~x11 && x6 && ~x4 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( x69 && ~x62 && ~x16 && x15 && x13 && ~x11 && ~x6 && x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( x69 && ~x62 && ~x16 && x15 && x13 && ~x11 && ~x6 && ~x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s477;
						end
					else if( x69 && ~x62 && ~x16 && x15 && ~x13 && x14 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x69 && ~x62 && ~x16 && x15 && ~x13 && ~x14 && x9 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x69 && ~x62 && ~x16 && x15 && ~x13 && ~x14 && ~x9 && x6 && x2 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x69 && ~x62 && ~x16 && x15 && ~x13 && ~x14 && ~x9 && x6 && ~x2 )
						nx_state = s478;
					else if( x69 && ~x62 && ~x16 && x15 && ~x13 && ~x14 && ~x9 && ~x6 && x8 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x69 && ~x62 && ~x16 && x15 && ~x13 && ~x14 && ~x9 && ~x6 && ~x8 )
						nx_state = s478;
					else if( x69 && ~x62 && ~x16 && ~x15 )
						nx_state = s1;
					else if( ~x69 && x28 && x64 && x43 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && x28 && x64 && ~x43 )
						nx_state = s478;
					else if( ~x69 && x28 && ~x64 && x49 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && x28 && ~x64 && ~x49 )
						nx_state = s478;
					else if( ~x69 && ~x28 && x27 && x8 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && ~x28 && x27 && ~x8 && x37 && x64 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && ~x28 && x27 && ~x8 && x37 && ~x64 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x69 && ~x28 && x27 && ~x8 && ~x37 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x69 && ~x28 && ~x27 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else nx_state = s478;
				s479 : if( x4 && x5 && x1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s477;
						end
					else if( x4 && x5 && ~x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s60;
						end
					else if( x4 && ~x5 && x1 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( x4 && ~x5 && ~x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x4 && x1 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x4 && ~x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else nx_state = s479;
				s480 : if( x69 && x62 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( x69 && ~x62 && x16 && x15 && x5 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else if( x69 && ~x62 && x16 && x15 && ~x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s634;
						end
					else if( x69 && ~x62 && x16 && ~x15 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( x69 && ~x62 && ~x16 && x15 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s634;
						end
					else if( x69 && ~x62 && ~x16 && x15 && ~x12 )
						nx_state = s480;
					else if( x69 && ~x62 && ~x16 && ~x15 && x13 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s638;
						end
					else if( x69 && ~x62 && ~x16 && ~x15 && ~x13 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s634;
						end
					else if( ~x69 && x15 && x13 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s704;
						end
					else if( ~x69 && x15 && ~x13 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s634;
						end
					else if( ~x69 && ~x15 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s634;
						end
					else if( ~x69 && ~x15 && ~x12 )
						nx_state = s480;
					else nx_state = s480;
				s481 : if( 1'b1 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s481;
				s482 : if( x17 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s1118;
						end
					else if( ~x17 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s482;
						end
					else nx_state = s482;
				s483 : if( x63 )
						nx_state = s1;
					else if( ~x63 && x64 && x11 && x10 )
						begin
							y62 = 1'b1;	
							nx_state = s1119;
						end
					else if( ~x63 && x64 && x11 && ~x10 && x4 && x5 && x3 && x12 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x63 && x64 && x11 && ~x10 && x4 && x5 && x3 && x12 && ~x8 && x7 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x63 && x64 && x11 && ~x10 && x4 && x5 && x3 && x12 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x63 && x64 && x11 && ~x10 && x4 && x5 && x3 && ~x12 )
						nx_state = s1;
					else if( ~x63 && x64 && x11 && ~x10 && x4 && x5 && ~x3 && x6 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x63 && x64 && x11 && ~x10 && x4 && x5 && ~x3 && x6 && ~x7 && x12 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x63 && x64 && x11 && ~x10 && x4 && x5 && ~x3 && x6 && ~x7 && x12 && ~x8 )
						nx_state = s1;
					else if( ~x63 && x64 && x11 && ~x10 && x4 && x5 && ~x3 && x6 && ~x7 && ~x12 )
						nx_state = s1;
					else if( ~x63 && x64 && x11 && ~x10 && x4 && x5 && ~x3 && ~x6 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x63 && x64 && x11 && ~x10 && x4 && x5 && ~x3 && ~x6 && ~x8 && x12 && x7 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x63 && x64 && x11 && ~x10 && x4 && x5 && ~x3 && ~x6 && ~x8 && x12 && ~x7 )
						nx_state = s1;
					else if( ~x63 && x64 && x11 && ~x10 && x4 && x5 && ~x3 && ~x6 && ~x8 && ~x12 )
						nx_state = s1;
					else if( ~x63 && x64 && x11 && ~x10 && x4 && ~x5 && x6 && x3 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x63 && x64 && x11 && ~x10 && x4 && ~x5 && x6 && ~x3 )
						begin
							y21 = 1'b1;	y38 = 1'b1;	
							nx_state = s412;
						end
					else if( ~x63 && x64 && x11 && ~x10 && x4 && ~x5 && ~x6 && x3 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x63 && x64 && x11 && ~x10 && x4 && ~x5 && ~x6 && ~x3 )
						begin
							y22 = 1'b1;	y29 = 1'b1;	
							nx_state = s412;
						end
					else if( ~x63 && x64 && x11 && ~x10 && ~x4 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x63 && x64 && ~x11 )
						begin
							y62 = 1'b1;	
							nx_state = s1120;
						end
					else if( ~x63 && ~x64 && x16 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x63 && ~x64 && ~x16 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x64 && ~x16 && x20 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x64 && ~x16 && x20 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x63 && ~x64 && ~x16 && ~x20 )
						nx_state = s1;
					else nx_state = s483;
				s484 : if( x69 && x70 && x62 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s1121;
						end
					else if( x69 && x70 && x62 && ~x17 )
						begin
							y1 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1122;
						end
					else if( x69 && x70 && ~x62 && x64 && x63 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x69 && x70 && ~x62 && x64 && x63 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x69 && x70 && ~x62 && x64 && x63 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && x63 && ~x10 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && x13 )
						begin
							y3 = 1'b1;	
							nx_state = s835;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && ~x13 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && ~x13 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x69 && x70 && ~x62 && x64 && ~x63 && ~x13 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && x64 && ~x63 && ~x13 && ~x14 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && x63 && x65 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && x65 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && x65 && x19 && ~x14 && ~x13 && x11 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && x65 && x19 && ~x14 && ~x13 && x11 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && x65 && x19 && ~x14 && ~x13 && ~x11 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( x69 && x70 && ~x62 && ~x64 && x63 && x65 && ~x19 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && x63 && ~x65 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && ~x63 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x63 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x69 && x70 && ~x62 && ~x64 && ~x63 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x69 && x70 && ~x62 && ~x64 && ~x63 && ~x23 )
						nx_state = s1;
					else if( x69 && ~x70 && x22 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s376;
						end
					else if( x69 && ~x70 && ~x22 )
						begin
							y3 = 1'b1;	
							nx_state = s835;
						end
					else if( ~x69 && x64 && x61 && x3 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && x64 && x61 && ~x3 && x2 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s933;
						end
					else if( ~x69 && x64 && x61 && ~x3 && ~x2 && x28 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x64 && x61 && ~x3 && ~x2 && ~x28 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x64 && ~x61 && x10 && x5 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s201;
						end
					else if( ~x69 && x64 && ~x61 && x10 && x5 && ~x3 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( ~x69 && x64 && ~x61 && x10 && x5 && ~x3 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x69 && x64 && ~x61 && x10 && ~x5 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && x64 && ~x61 && ~x10 && x11 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s759;
						end
					else if( ~x69 && x64 && ~x61 && ~x10 && x11 && ~x1 && x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && x64 && ~x61 && ~x10 && x11 && ~x1 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && x64 && ~x61 && ~x10 && ~x11 )
						nx_state = s484;
					else if( ~x69 && ~x64 && x14 && x3 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && ~x64 && x14 && ~x3 && x2 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s933;
						end
					else if( ~x69 && ~x64 && x14 && ~x3 && ~x2 && x28 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && ~x64 && x14 && ~x3 && ~x2 && ~x28 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && ~x64 && ~x14 && x10 && x5 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s201;
						end
					else if( ~x69 && ~x64 && ~x14 && x10 && x5 && ~x3 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( ~x69 && ~x64 && ~x14 && x10 && x5 && ~x3 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x69 && ~x64 && ~x14 && x10 && ~x5 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && ~x64 && ~x14 && ~x10 && x11 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s759;
						end
					else if( ~x69 && ~x64 && ~x14 && ~x10 && x11 && ~x1 && x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && ~x64 && ~x14 && ~x10 && x11 && ~x1 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x69 && ~x64 && ~x14 && ~x10 && ~x11 )
						nx_state = s484;
					else nx_state = s484;
				s485 : if( x63 && x7 )
						begin
							y69 = 1'b1;	
							nx_state = s1123;
						end
					else if( x63 && ~x7 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( ~x63 )
						nx_state = s1;
					else nx_state = s485;
				s486 : if( x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x22 && ~x17 )
						nx_state = s1;
					else if( ~x22 && x18 && x13 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x22 && x18 && x13 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x22 && x18 && ~x13 && x12 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x22 && x18 && ~x13 && x12 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x22 && ~x18 )
						nx_state = s1;
					else nx_state = s486;
				s487 : if( x60 && x61 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x60 && ~x61 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x60 && ~x61 && ~x2 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x60 && x61 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x60 && x61 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x60 && x61 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( ~x60 && x61 && x62 && ~x18 )
						nx_state = s1;
					else if( ~x60 && x61 && ~x62 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x60 && x61 && ~x62 && ~x2 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x60 && ~x61 && x62 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x60 && ~x61 && x62 && ~x7 )
						nx_state = s47;
					else if( ~x60 && ~x61 && ~x62 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else nx_state = s487;
				s488 : if( 1'b1 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s792;
						end
					else nx_state = s488;
				s489 : if( 1'b1 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else nx_state = s489;
				s490 : if( x65 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x65 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else nx_state = s490;
				s491 : if( x65 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x65 )
						begin
							y17 = 1'b1;	
							nx_state = s98;
						end
					else nx_state = s491;
				s492 : if( x21 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x21 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x21 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x21 && ~x9 )
						nx_state = s1;
					else if( ~x21 && x22 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x21 && ~x22 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s492;
				s493 : if( x66 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x66 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else nx_state = s493;
				s494 : if( x21 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x21 && x23 && x22 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x21 && x23 && ~x22 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x21 && ~x23 && x22 && x17 && x15 && x9 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( ~x21 && ~x23 && x22 && x17 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x21 && ~x23 && x22 && x17 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x23 && x22 && x17 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s495;
						end
					else if( ~x21 && ~x23 && x22 && ~x17 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x21 && ~x23 && ~x22 && x2 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x2 && x17 && x15 && x9 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x2 && x17 && x15 && ~x9 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x2 && x17 && ~x15 && x16 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x2 && x17 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s495;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x2 && ~x17 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else nx_state = s494;
				s495 : if( x21 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x21 && x22 && x23 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x21 && x22 && ~x23 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s406;
						end
					else if( ~x21 && ~x22 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s406;
						end
					else nx_state = s495;
				s496 : if( x69 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x69 && x26 && x28 && x62 && x3 && x5 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s612;
						end
					else if( ~x69 && x26 && x28 && x62 && x3 && ~x5 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s614;
						end
					else if( ~x69 && x26 && x28 && x62 && ~x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s942;
						end
					else if( ~x69 && x26 && x28 && ~x62 && x3 && x63 && x5 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s1124;
						end
					else if( ~x69 && x26 && x28 && ~x62 && x3 && x63 && ~x5 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s995;
						end
					else if( ~x69 && x26 && x28 && ~x62 && x3 && ~x63 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s920;
						end
					else if( ~x69 && x26 && x28 && ~x62 && x3 && ~x63 && ~x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else if( ~x69 && x26 && x28 && ~x62 && ~x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else if( ~x69 && x26 && ~x28 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( ~x69 && ~x26 && x27 && x62 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( ~x69 && ~x26 && x27 && ~x62 && x63 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x69 && ~x26 && x27 && ~x62 && ~x63 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && ~x26 && ~x27 && x28 && x62 && x5 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s941;
						end
					else if( ~x69 && ~x26 && ~x27 && x28 && x62 && ~x5 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s614;
						end
					else if( ~x69 && ~x26 && ~x27 && x28 && ~x62 && x63 && x36 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( ~x69 && ~x26 && ~x27 && x28 && ~x62 && x63 && ~x36 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s995;
						end
					else if( ~x69 && ~x26 && ~x27 && x28 && ~x62 && ~x63 && x5 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( ~x69 && ~x26 && ~x27 && x28 && ~x62 && ~x63 && ~x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && x62 && x5 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s613;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && x62 && x5 && ~x3 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && x62 && x5 && ~x3 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s614;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && x62 && ~x5 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && ~x62 && x63 && x36 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s922;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && ~x62 && x63 && x36 && ~x3 && x4 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s994;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && ~x62 && x63 && x36 && ~x3 && ~x4 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s995;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && ~x62 && x63 && ~x36 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && ~x62 && ~x63 && x5 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s922;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && ~x62 && ~x63 && x5 && ~x3 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && ~x62 && ~x63 && x5 && ~x3 && ~x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && ~x62 && ~x63 && ~x5 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else nx_state = s496;
				s497 : if( x24 && x26 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x24 && x26 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x24 && x26 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x24 && x26 && ~x18 )
						nx_state = s1;
					else if( x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x24 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x24 && x25 && x19 && ~x14 && ~x13 && x26 )
						nx_state = s497;
					else if( ~x24 && x25 && x19 && ~x14 && ~x13 && ~x26 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && x10 && x12 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x24 && ~x25 && ~x26 && x10 && x12 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x24 && ~x25 && ~x26 && x10 && x12 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && x10 && x12 && ~x17 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && x10 && ~x12 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x10 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x10 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x10 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && ~x10 && ~x17 )
						nx_state = s1;
					else nx_state = s497;
				s498 : if( x69 )
						nx_state = s1;
					else if( ~x69 && x63 && x55 && x35 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && x63 && x55 && ~x35 && x13 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s504;
						end
					else if( ~x69 && x63 && x55 && ~x35 && ~x13 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s456;
						end
					else if( ~x69 && x63 && ~x55 && x41 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( ~x69 && x63 && ~x55 && ~x41 && x42 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s504;
						end
					else if( ~x69 && x63 && ~x55 && ~x41 && ~x42 && x38 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x69 && x63 && ~x55 && ~x41 && ~x42 && ~x38 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s818;
						end
					else if( ~x69 && ~x63 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else nx_state = s498;
				s499 : if( x63 && x55 && x50 && x41 && x19 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( x63 && x55 && x50 && x41 && ~x19 )
						nx_state = s499;
					else if( x63 && x55 && x50 && ~x41 && x19 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( x63 && x55 && x50 && ~x41 && ~x19 )
						nx_state = s499;
					else if( x63 && x55 && ~x50 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( x63 && ~x55 && x10 && x11 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x63 && ~x55 && x10 && ~x11 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( x63 && ~x55 && ~x10 && x42 && x38 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s498;
						end
					else if( x63 && ~x55 && ~x10 && x42 && ~x38 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x63 && ~x55 && ~x10 && ~x42 && x12 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s504;
						end
					else if( x63 && ~x55 && ~x10 && ~x42 && ~x12 && x1 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y33 = 1'b1;	
							nx_state = s506;
						end
					else if( x63 && ~x55 && ~x10 && ~x42 && ~x12 && ~x1 && x35 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( x63 && ~x55 && ~x10 && ~x42 && ~x12 && ~x1 && ~x35 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x63 && x40 && x50 && x19 && x10 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x63 && x40 && x50 && x19 && ~x10 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x63 && x40 && x50 && ~x19 )
						nx_state = s499;
					else if( ~x63 && x40 && ~x50 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x63 && ~x40 && x11 && x10 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x63 && ~x40 && x11 && ~x10 && x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s507;
						end
					else if( ~x63 && ~x40 && x11 && ~x10 && ~x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1106;
						end
					else if( ~x63 && ~x40 && ~x11 && x10 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x63 && ~x40 && ~x11 && ~x10 && x12 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s510;
						end
					else if( ~x63 && ~x40 && ~x11 && ~x10 && ~x12 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s449;
						end
					else if( ~x63 && ~x40 && ~x11 && ~x10 && ~x12 && ~x1 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x63 && ~x40 && ~x11 && ~x10 && ~x12 && ~x1 && ~x4 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else nx_state = s499;
				s500 : if( x63 && x50 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s503;
						end
					else if( x63 && ~x50 )
						nx_state = s500;
					else if( ~x63 && x50 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x63 && ~x50 )
						nx_state = s500;
					else nx_state = s500;
				s501 : if( x55 && x47 && x54 && x29 && x59 && x27 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s1125;
						end
					else if( x55 && x47 && x54 && x29 && x59 && ~x27 )
						nx_state = s501;
					else if( x55 && x47 && x54 && x29 && ~x59 && x27 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( x55 && x47 && x54 && x29 && ~x59 && ~x27 )
						nx_state = s501;
					else if( x55 && x47 && x54 && ~x29 && x33 && x27 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( x55 && x47 && x54 && ~x29 && x33 && ~x27 )
						nx_state = s501;
					else if( x55 && x47 && x54 && ~x29 && ~x33 && x57 && x27 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( x55 && x47 && x54 && ~x29 && ~x33 && x57 && ~x27 )
						nx_state = s501;
					else if( x55 && x47 && x54 && ~x29 && ~x33 && ~x57 && x27 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( x55 && x47 && x54 && ~x29 && ~x33 && ~x57 && ~x27 )
						nx_state = s501;
					else if( x55 && x47 && ~x54 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x55 && ~x47 && x37 && x56 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( x55 && ~x47 && x37 && x56 && ~x1 )
						nx_state = s501;
					else if( x55 && ~x47 && x37 && ~x56 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x55 && ~x47 && ~x37 && x25 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x55 && ~x47 && ~x37 && ~x25 && x36 && x35 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s456;
						end
					else if( x55 && ~x47 && ~x37 && ~x25 && x36 && ~x35 )
						nx_state = s501;
					else if( x55 && ~x47 && ~x37 && ~x25 && ~x36 && x35 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( x55 && ~x47 && ~x37 && ~x25 && ~x36 && ~x35 )
						nx_state = s501;
					else if( ~x55 && x41 && x11 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x55 && x41 && ~x11 && x12 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x55 && x41 && ~x11 && x12 && ~x2 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x55 && x41 && ~x11 && ~x12 && x32 && x3 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( ~x55 && x41 && ~x11 && ~x12 && x32 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x55 && x41 && ~x11 && ~x12 && x32 && ~x3 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x55 && x41 && ~x11 && ~x12 && ~x32 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x55 && ~x41 && x43 && x33 && x35 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x55 && ~x41 && x43 && x33 && ~x35 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x55 && ~x41 && x43 && ~x33 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x55 && ~x41 && ~x43 && x40 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y31 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s1126;
						end
					else if( ~x55 && ~x41 && ~x43 && ~x40 && x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( ~x55 && ~x41 && ~x43 && ~x40 && ~x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else nx_state = s501;
				s502 : if( x55 && x51 && x24 && x36 )
						nx_state = s502;
					else if( x55 && x51 && x24 && ~x36 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( x55 && x51 && ~x24 && x31 && x29 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s498;
						end
					else if( x55 && x51 && ~x24 && x31 && ~x29 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( x55 && x51 && ~x24 && ~x31 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s498;
						end
					else if( x55 && ~x51 && x42 && x35 && x36 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s498;
						end
					else if( x55 && ~x51 && x42 && x35 && ~x36 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( x55 && ~x51 && x42 && ~x35 && x58 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x55 && ~x51 && x42 && ~x35 && ~x58 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( x55 && ~x51 && ~x42 && x52 && x35 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y27 = 1'b1;	
							nx_state = s833;
						end
					else if( x55 && ~x51 && ~x42 && x52 && ~x35 && x58 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x55 && ~x51 && ~x42 && x52 && ~x35 && ~x58 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( x55 && ~x51 && ~x42 && ~x52 && x3 && x6 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s504;
						end
					else if( x55 && ~x51 && ~x42 && ~x52 && x3 && ~x6 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( x55 && ~x51 && ~x42 && ~x52 && ~x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( ~x55 && x10 && x11 && x34 && x35 )
						nx_state = s502;
					else if( ~x55 && x10 && x11 && x34 && ~x35 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( ~x55 && x10 && x11 && ~x34 && x4 && x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x55 && x10 && x11 && ~x34 && x4 && ~x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x55 && x10 && x11 && ~x34 && ~x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s503;
						end
					else if( ~x55 && x10 && ~x11 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x55 && x10 && ~x11 && ~x2 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x55 && ~x10 && x42 && x37 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( ~x55 && ~x10 && x42 && ~x37 && x8 && x4 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s456;
						end
					else if( ~x55 && ~x10 && x42 && ~x37 && x8 && ~x4 && x1 && x34 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x55 && ~x10 && x42 && ~x37 && x8 && ~x4 && x1 && ~x34 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x55 && ~x10 && x42 && ~x37 && x8 && ~x4 && ~x1 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x55 && ~x10 && x42 && ~x37 && ~x8 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x55 && ~x10 && ~x42 && x12 && x9 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x55 && ~x10 && ~x42 && x12 && ~x9 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y27 = 1'b1;	
							nx_state = s833;
						end
					else if( ~x55 && ~x10 && ~x42 && ~x12 && x6 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x55 && ~x10 && ~x42 && ~x12 && ~x6 && x40 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( ~x55 && ~x10 && ~x42 && ~x12 && ~x6 && ~x40 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else nx_state = s502;
				s503 : if( x55 && x44 && x23 && x51 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s498;
						end
					else if( x55 && x44 && x23 && ~x51 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( x55 && x44 && ~x23 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s498;
						end
					else if( x55 && ~x44 && x28 && x35 && x36 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s498;
						end
					else if( x55 && ~x44 && x28 && x35 && ~x36 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( x55 && ~x44 && x28 && ~x35 && x58 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x55 && ~x44 && x28 && ~x35 && ~x58 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( x55 && ~x44 && ~x28 && x37 && x35 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y27 = 1'b1;	
							nx_state = s833;
						end
					else if( x55 && ~x44 && ~x28 && x37 && ~x35 && x58 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x55 && ~x44 && ~x28 && x37 && ~x35 && ~x58 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( x55 && ~x44 && ~x28 && ~x37 && x39 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( x55 && ~x44 && ~x28 && ~x37 && ~x39 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x55 && x41 && x11 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x55 && x41 && ~x11 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( ~x55 && ~x41 && x42 && x32 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s882;
						end
					else if( ~x55 && ~x41 && x42 && ~x32 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x55 && ~x41 && x42 && ~x32 && ~x3 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x55 && ~x41 && ~x42 && x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( ~x55 && ~x41 && ~x42 && ~x5 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else nx_state = s503;
				s504 : if( x69 && x12 && x13 && x3 )
						begin
							y3 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s881;
						end
					else if( x69 && x12 && x13 && ~x3 && x14 )
						begin
							y3 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s881;
						end
					else if( x69 && x12 && x13 && ~x3 && ~x14 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s882;
						end
					else if( x69 && x12 && ~x13 )
						begin
							y3 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s883;
						end
					else if( x69 && ~x12 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							y16 = 1'b1;	y21 = 1'b1;	
							nx_state = s884;
						end
					else if( ~x69 && x63 && x55 && x8 && x53 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s818;
						end
					else if( ~x69 && x63 && x55 && x8 && ~x53 && x37 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && x63 && x55 && x8 && ~x53 && ~x37 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s818;
						end
					else if( ~x69 && x63 && x55 && ~x8 && x51 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s818;
						end
					else if( ~x69 && x63 && x55 && ~x8 && ~x51 && x37 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && x63 && x55 && ~x8 && ~x51 && ~x37 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s818;
						end
					else if( ~x69 && x63 && ~x55 && x41 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x69 && x63 && ~x55 && ~x41 && x42 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s504;
						end
					else if( ~x69 && x63 && ~x55 && ~x41 && ~x42 && x43 && x39 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s498;
						end
					else if( ~x69 && x63 && ~x55 && ~x41 && ~x42 && x43 && ~x39 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x69 && x63 && ~x55 && ~x41 && ~x42 && ~x43 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							y16 = 1'b1;	y21 = 1'b1;	
							nx_state = s884;
						end
					else if( ~x69 && ~x63 && x40 && x37 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && ~x63 && x40 && ~x37 && x9 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && ~x63 && x40 && ~x37 && ~x9 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x69 && ~x63 && ~x40 && x10 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && ~x63 && ~x40 && ~x10 && x11 && x1 )
						begin
							y3 = 1'b1;	y13 = 1'b1;	y18 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s639;
						end
					else if( ~x69 && ~x63 && ~x40 && ~x10 && x11 && ~x1 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && ~x63 && ~x40 && ~x10 && x11 && ~x1 && ~x3 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x69 && ~x63 && ~x40 && ~x10 && ~x11 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else nx_state = s504;
				s505 : if( x7 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y33 = 1'b1;	
							nx_state = s506;
						end
					else if( ~x7 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else nx_state = s505;
				s506 : if( x55 && x29 && x50 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x55 && x29 && ~x50 )
						nx_state = s506;
					else if( x55 && ~x29 && x58 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x55 && ~x29 && ~x58 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( ~x55 && x11 && x6 && x40 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( ~x55 && x11 && x6 && ~x40 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s882;
						end
					else if( ~x55 && x11 && ~x6 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s504;
						end
					else if( ~x55 && ~x11 && x39 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( ~x55 && ~x11 && ~x39 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s456;
						end
					else nx_state = s506;
				s507 : if( x40 && x35 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x40 && ~x35 && x13 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s510;
						end
					else if( x40 && ~x35 && ~x13 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else if( ~x40 && x10 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x40 && ~x10 && x11 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s510;
						end
					else if( ~x40 && ~x10 && ~x11 && x7 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x40 && ~x10 && ~x11 && ~x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else nx_state = s507;
				s508 : if( x64 && x40 && x16 && x45 && x29 && x42 && x27 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s686;
						end
					else if( x64 && x40 && x16 && x45 && x29 && x42 && ~x27 )
						nx_state = s508;
					else if( x64 && x40 && x16 && x45 && x29 && ~x42 && x27 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( x64 && x40 && x16 && x45 && x29 && ~x42 && ~x27 )
						nx_state = s508;
					else if( x64 && x40 && x16 && x45 && ~x29 && x33 && x27 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( x64 && x40 && x16 && x45 && ~x29 && x33 && ~x27 )
						nx_state = s508;
					else if( x64 && x40 && x16 && x45 && ~x29 && ~x33 && x43 && x27 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( x64 && x40 && x16 && x45 && ~x29 && ~x33 && x43 && ~x27 )
						nx_state = s508;
					else if( x64 && x40 && x16 && x45 && ~x29 && ~x33 && ~x43 && x27 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( x64 && x40 && x16 && x45 && ~x29 && ~x33 && ~x43 && ~x27 )
						nx_state = s508;
					else if( x64 && x40 && x16 && ~x45 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x64 && x40 && ~x16 && x37 && x44 && x1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( x64 && x40 && ~x16 && x37 && x44 && ~x1 )
						nx_state = s508;
					else if( x64 && x40 && ~x16 && x37 && ~x44 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x64 && x40 && ~x16 && ~x37 && x25 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x64 && x40 && ~x16 && ~x37 && ~x25 && x5 && x4 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else if( x64 && x40 && ~x16 && ~x37 && ~x25 && x5 && ~x4 )
						nx_state = s508;
					else if( x64 && x40 && ~x16 && ~x37 && ~x25 && ~x5 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( x64 && x40 && ~x16 && ~x37 && ~x25 && ~x5 && ~x4 )
						nx_state = s508;
					else if( x64 && ~x40 && x10 && x11 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( x64 && ~x40 && x10 && ~x11 && x12 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( x64 && ~x40 && x10 && ~x11 && x12 && ~x2 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x64 && ~x40 && x10 && ~x11 && ~x12 && x1 && x3 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( x64 && ~x40 && x10 && ~x11 && ~x12 && x1 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( x64 && ~x40 && x10 && ~x11 && ~x12 && x1 && ~x3 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( x64 && ~x40 && x10 && ~x11 && ~x12 && ~x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( x64 && ~x40 && ~x10 && x12 && x2 && x4 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( x64 && ~x40 && ~x10 && x12 && x2 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( x64 && ~x40 && ~x10 && x12 && ~x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( x64 && ~x40 && ~x10 && ~x12 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s1105;
						end
					else if( x64 && ~x40 && ~x10 && ~x12 && ~x9 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( x64 && ~x40 && ~x10 && ~x12 && ~x9 && ~x5 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x64 && x44 && x16 && x54 && x29 && x48 && x27 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s686;
						end
					else if( ~x64 && x44 && x16 && x54 && x29 && x48 && ~x27 )
						nx_state = s508;
					else if( ~x64 && x44 && x16 && x54 && x29 && ~x48 && x27 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x64 && x44 && x16 && x54 && x29 && ~x48 && ~x27 )
						nx_state = s508;
					else if( ~x64 && x44 && x16 && x54 && ~x29 && x33 && x27 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x64 && x44 && x16 && x54 && ~x29 && x33 && ~x27 )
						nx_state = s508;
					else if( ~x64 && x44 && x16 && x54 && ~x29 && ~x33 && x49 && x27 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x64 && x44 && x16 && x54 && ~x29 && ~x33 && x49 && ~x27 )
						nx_state = s508;
					else if( ~x64 && x44 && x16 && x54 && ~x29 && ~x33 && ~x49 && x27 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x64 && x44 && x16 && x54 && ~x29 && ~x33 && ~x49 && ~x27 )
						nx_state = s508;
					else if( ~x64 && x44 && x16 && ~x54 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x64 && x44 && ~x16 && x36 && x55 && x37 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x64 && x44 && ~x16 && x36 && x55 && ~x37 )
						nx_state = s508;
					else if( ~x64 && x44 && ~x16 && x36 && ~x55 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x64 && x44 && ~x16 && ~x36 && x25 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x64 && x44 && ~x16 && ~x36 && ~x25 && x5 && x4 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else if( ~x64 && x44 && ~x16 && ~x36 && ~x25 && x5 && ~x4 )
						nx_state = s508;
					else if( ~x64 && x44 && ~x16 && ~x36 && ~x25 && ~x5 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x64 && x44 && ~x16 && ~x36 && ~x25 && ~x5 && ~x4 )
						nx_state = s508;
					else if( ~x64 && ~x44 && x10 && x11 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else if( ~x64 && ~x44 && x10 && ~x11 && x12 && x34 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else if( ~x64 && ~x44 && x10 && ~x11 && x12 && ~x34 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x64 && ~x44 && x10 && ~x11 && ~x12 && x37 && x41 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x64 && ~x44 && x10 && ~x11 && ~x12 && x37 && ~x41 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x64 && ~x44 && x10 && ~x11 && ~x12 && x37 && ~x41 && ~x4 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s631;
						end
					else if( ~x64 && ~x44 && x10 && ~x11 && ~x12 && ~x37 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else if( ~x64 && ~x44 && ~x10 && x12 && x2 && x4 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x64 && ~x44 && ~x10 && x12 && x2 && ~x4 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s631;
						end
					else if( ~x64 && ~x44 && ~x10 && x12 && ~x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else if( ~x64 && ~x44 && ~x10 && ~x12 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s1105;
						end
					else if( ~x64 && ~x44 && ~x10 && ~x12 && ~x9 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x64 && ~x44 && ~x10 && ~x12 && ~x9 && ~x5 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else nx_state = s508;
				s509 : if( x64 && x40 && x51 && x24 && x5 && x36 )
						nx_state = s509;
					else if( x64 && x40 && x51 && x24 && x5 && ~x36 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s507;
						end
					else if( x64 && x40 && x51 && x24 && ~x5 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( x64 && x40 && x51 && ~x24 && x31 && x29 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s507;
						end
					else if( x64 && x40 && x51 && ~x24 && x31 && ~x29 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( x64 && x40 && x51 && ~x24 && ~x31 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s507;
						end
					else if( x64 && x40 && ~x51 && x11 && x35 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s507;
						end
					else if( x64 && x40 && ~x51 && x11 && x35 && ~x5 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( x64 && x40 && ~x51 && x11 && ~x35 && x41 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x64 && x40 && ~x51 && x11 && ~x35 && ~x41 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( x64 && x40 && ~x51 && ~x11 && x49 && x35 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s638;
						end
					else if( x64 && x40 && ~x51 && ~x11 && x49 && ~x35 && x41 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x64 && x40 && ~x51 && ~x11 && x49 && ~x35 && ~x41 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( x64 && x40 && ~x51 && ~x11 && ~x49 && x3 && x6 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s510;
						end
					else if( x64 && x40 && ~x51 && ~x11 && ~x49 && x3 && ~x6 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( x64 && x40 && ~x51 && ~x11 && ~x49 && ~x3 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( x64 && ~x40 && x11 && x10 && x4 && x5 && x3 )
						nx_state = s509;
					else if( x64 && ~x40 && x11 && x10 && x4 && x5 && ~x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( x64 && ~x40 && x11 && x10 && x4 && ~x5 && x3 )
						nx_state = s509;
					else if( x64 && ~x40 && x11 && x10 && x4 && ~x5 && ~x3 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( x64 && ~x40 && x11 && x10 && ~x4 && x3 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( x64 && ~x40 && x11 && x10 && ~x4 && ~x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( x64 && ~x40 && x11 && ~x10 && x6 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( x64 && ~x40 && x11 && ~x10 && ~x6 && x8 && x4 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else if( x64 && ~x40 && x11 && ~x10 && ~x6 && x8 && ~x4 && x1 && x3 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( x64 && ~x40 && x11 && ~x10 && ~x6 && x8 && ~x4 && x1 && ~x3 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( x64 && ~x40 && x11 && ~x10 && ~x6 && x8 && ~x4 && ~x1 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( x64 && ~x40 && x11 && ~x10 && ~x6 && ~x8 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x64 && ~x40 && ~x11 && x10 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( x64 && ~x40 && ~x11 && x10 && ~x2 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x64 && ~x40 && ~x11 && ~x10 && x12 && x9 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x64 && ~x40 && ~x11 && ~x10 && x12 && ~x9 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s638;
						end
					else if( x64 && ~x40 && ~x11 && ~x10 && ~x12 && x6 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( x64 && ~x40 && ~x11 && ~x10 && ~x12 && ~x6 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( x64 && ~x40 && ~x11 && ~x10 && ~x12 && ~x6 && ~x9 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x64 && x44 && x51 && x24 && x5 && x36 )
						nx_state = s509;
					else if( ~x64 && x44 && x51 && x24 && x5 && ~x36 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s511;
						end
					else if( ~x64 && x44 && x51 && x24 && ~x5 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x64 && x44 && x51 && ~x24 && x31 && x29 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s511;
						end
					else if( ~x64 && x44 && x51 && ~x24 && x31 && ~x29 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x64 && x44 && x51 && ~x24 && ~x31 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s511;
						end
					else if( ~x64 && x44 && ~x51 && x11 && x35 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s511;
						end
					else if( ~x64 && x44 && ~x51 && x11 && x35 && ~x5 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x64 && x44 && ~x51 && x11 && ~x35 && x45 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x64 && x44 && ~x51 && x11 && ~x35 && ~x45 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x64 && x44 && ~x51 && ~x11 && x52 && x35 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s638;
						end
					else if( ~x64 && x44 && ~x51 && ~x11 && x52 && ~x35 && x45 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x64 && x44 && ~x51 && ~x11 && x52 && ~x35 && ~x45 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x64 && x44 && ~x51 && ~x11 && ~x52 && x41 && x6 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s510;
						end
					else if( ~x64 && x44 && ~x51 && ~x11 && ~x52 && x41 && ~x6 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x64 && x44 && ~x51 && ~x11 && ~x52 && ~x41 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x64 && ~x44 && x10 && x11 && x4 && x5 && x3 )
						nx_state = s509;
					else if( ~x64 && ~x44 && x10 && x11 && x4 && x5 && ~x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else if( ~x64 && ~x44 && x10 && x11 && x4 && ~x5 && x3 )
						nx_state = s509;
					else if( ~x64 && ~x44 && x10 && x11 && x4 && ~x5 && ~x3 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x64 && ~x44 && x10 && x11 && ~x4 && x3 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x64 && ~x44 && x10 && x11 && ~x4 && ~x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x64 && ~x44 && x10 && ~x11 && x34 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else if( ~x64 && ~x44 && x10 && ~x11 && ~x34 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x64 && ~x44 && ~x10 && x11 && x6 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x64 && ~x44 && ~x10 && x11 && ~x6 && x8 && x4 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else if( ~x64 && ~x44 && ~x10 && x11 && ~x6 && x8 && ~x4 && x1 && x41 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x64 && ~x44 && ~x10 && x11 && ~x6 && x8 && ~x4 && x1 && ~x41 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x64 && ~x44 && ~x10 && x11 && ~x6 && x8 && ~x4 && ~x1 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s631;
						end
					else if( ~x64 && ~x44 && ~x10 && x11 && ~x6 && ~x8 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x64 && ~x44 && ~x10 && ~x11 && x12 && x9 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x64 && ~x44 && ~x10 && ~x11 && x12 && ~x9 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s638;
						end
					else if( ~x64 && ~x44 && ~x10 && ~x11 && ~x12 && x6 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x64 && ~x44 && ~x10 && ~x11 && ~x12 && ~x6 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x64 && ~x44 && ~x10 && ~x11 && ~x12 && ~x6 && ~x9 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else nx_state = s509;
				s510 : if( x64 && x40 && x8 && x48 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x64 && x40 && x8 && ~x48 && x37 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x64 && x40 && x8 && ~x48 && ~x37 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x64 && x40 && ~x8 && x51 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x64 && x40 && ~x8 && ~x51 && x37 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x64 && x40 && ~x8 && ~x51 && ~x37 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x64 && ~x40 && x10 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( x64 && ~x40 && ~x10 && x11 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s510;
						end
					else if( x64 && ~x40 && ~x10 && ~x11 && x12 && x8 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s507;
						end
					else if( x64 && ~x40 && ~x10 && ~x11 && x12 && ~x8 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1106;
						end
					else if( x64 && ~x40 && ~x10 && ~x11 && ~x12 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s504;
						end
					else if( ~x64 && x44 && x8 && x53 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x64 && x44 && x8 && ~x53 && x37 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x64 && x44 && x8 && ~x53 && ~x37 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x64 && x44 && ~x8 && x51 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x64 && x44 && ~x8 && ~x51 && x37 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x64 && x44 && ~x8 && ~x51 && ~x37 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x64 && ~x44 && x10 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s631;
						end
					else if( ~x64 && ~x44 && ~x10 && x11 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s510;
						end
					else if( ~x64 && ~x44 && ~x10 && ~x11 && x12 && x8 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s511;
						end
					else if( ~x64 && ~x44 && ~x10 && ~x11 && x12 && ~x8 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s1107;
						end
					else if( ~x64 && ~x44 && ~x10 && ~x11 && ~x12 )
						begin
							y17 = 1'b1;	y21 = 1'b1;	y32 = 1'b1;	
							nx_state = s1127;
						end
					else nx_state = s510;
				s511 : if( x44 && x35 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( x44 && ~x35 && x13 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s510;
						end
					else if( x44 && ~x35 && ~x13 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else if( ~x44 && x10 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x44 && ~x10 && x11 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s510;
						end
					else if( ~x44 && ~x10 && ~x11 && x7 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x44 && ~x10 && ~x11 && ~x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else nx_state = s511;
				s512 : if( x44 && x50 && x19 && x10 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( x44 && x50 && x19 && ~x10 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s631;
						end
					else if( x44 && x50 && ~x19 )
						nx_state = s512;
					else if( x44 && ~x50 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x44 && x10 && x11 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x44 && x10 && ~x11 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s631;
						end
					else if( ~x44 && ~x10 && x11 && x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s511;
						end
					else if( ~x44 && ~x10 && x11 && ~x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s1107;
						end
					else if( ~x44 && ~x10 && ~x11 && x12 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s510;
						end
					else if( ~x44 && ~x10 && ~x11 && ~x12 && x37 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s449;
						end
					else if( ~x44 && ~x10 && ~x11 && ~x12 && ~x37 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x44 && ~x10 && ~x11 && ~x12 && ~x37 && ~x4 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else nx_state = s512;
				s513 : if( x44 && x53 && x47 )
						nx_state = s513;
					else if( x44 && x53 && ~x47 && x48 && x51 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( x44 && x53 && ~x47 && x48 && ~x51 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( x44 && x53 && ~x47 && ~x48 && x34 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( x44 && x53 && ~x47 && ~x48 && ~x34 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( x44 && ~x53 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x44 && x11 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x44 && ~x11 && x1 && x34 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x44 && ~x11 && x1 && ~x34 && x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x44 && ~x11 && x1 && ~x34 && ~x3 )
						nx_state = s513;
					else if( ~x44 && ~x11 && ~x1 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else nx_state = s513;
				s514 : if( x7 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s449;
						end
					else if( ~x7 && x64 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x7 && ~x64 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s631;
						end
					else nx_state = s514;
				s515 : if( x24 && x26 )
						begin
							y17 = 1'b1;	
							nx_state = s1128;
						end
					else if( x24 && ~x26 && x16 && x11 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s368;
						end
					else if( x24 && ~x26 && x16 && x11 && ~x12 && x13 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( x24 && ~x26 && x16 && x11 && ~x12 && ~x13 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x24 && ~x26 && x16 && ~x11 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s300;
						end
					else if( x24 && ~x26 && ~x16 && x17 && x11 && x13 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( x24 && ~x26 && ~x16 && x17 && x11 && ~x13 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s122;
						end
					else if( x24 && ~x26 && ~x16 && x17 && ~x11 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( x24 && ~x26 && ~x16 && ~x17 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x24 && x25 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x24 && ~x25 && x26 && x16 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x24 && ~x25 && x26 && x16 && ~x11 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x24 && ~x25 && x26 && x16 && ~x11 && ~x12 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x24 && ~x25 && x26 && x16 && ~x11 && ~x12 && ~x10 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( ~x24 && ~x25 && x26 && ~x16 && x17 && x10 && x12 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x24 && ~x25 && x26 && ~x16 && x17 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x24 && ~x25 && x26 && ~x16 && x17 && ~x10 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x24 && ~x25 && x26 && ~x16 && ~x17 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x24 && ~x25 && ~x26 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s429;
						end
					else nx_state = s515;
				s516 : if( x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x6 )
						nx_state = s1;
					else nx_state = s516;
				s517 : if( x15 )
						begin
							y44 = 1'b1;	y45 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x15 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x15 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x15 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x15 && ~x6 )
						nx_state = s1;
					else nx_state = s517;
				s518 : if( x9 && x21 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1129;
						end
					else if( x9 && ~x21 && x22 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1130;
						end
					else if( x9 && ~x21 && ~x22 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1131;
						end
					else if( ~x9 && x13 && x21 && x10 )
						begin
							y62 = 1'b1;	y65 = 1'b1;	y78 = 1'b1;	
							y90 = 1'b1;	
							nx_state = s1132;
						end
					else if( ~x9 && x13 && x21 && ~x10 && x14 && x11 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1130;
						end
					else if( ~x9 && x13 && x21 && ~x10 && x14 && ~x11 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1133;
						end
					else if( ~x9 && x13 && x21 && ~x10 && ~x14 && x11 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1134;
						end
					else if( ~x9 && x13 && x21 && ~x10 && ~x14 && ~x11 )
						begin
							y3 = 1'b1;	y74 = 1'b1;	
							nx_state = s1135;
						end
					else if( ~x9 && x13 && ~x21 && x10 && x22 && x11 && x14 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1134;
						end
					else if( ~x9 && x13 && ~x21 && x10 && x22 && x11 && ~x14 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1131;
						end
					else if( ~x9 && x13 && ~x21 && x10 && x22 && ~x11 && x14 && x19 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x9 && x13 && ~x21 && x10 && x22 && ~x11 && x14 && ~x19 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x9 && x13 && ~x21 && x10 && x22 && ~x11 && x14 && ~x19 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x9 && x13 && ~x21 && x10 && x22 && ~x11 && x14 && ~x19 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x9 && x13 && ~x21 && x10 && x22 && ~x11 && x14 && ~x19 && ~x6 )
						nx_state = s1;
					else if( ~x9 && x13 && ~x21 && x10 && x22 && ~x11 && ~x14 && x18 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x9 && x13 && ~x21 && x10 && x22 && ~x11 && ~x14 && ~x18 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x9 && x13 && ~x21 && x10 && x22 && ~x11 && ~x14 && ~x18 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x9 && x13 && ~x21 && x10 && x22 && ~x11 && ~x14 && ~x18 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x9 && x13 && ~x21 && x10 && x22 && ~x11 && ~x14 && ~x18 && ~x6 )
						nx_state = s1;
					else if( ~x9 && x13 && ~x21 && x10 && ~x22 )
						begin
							y9 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y94 = 1'b1;	
							nx_state = s849;
						end
					else if( ~x9 && x13 && ~x21 && ~x10 && x22 && x14 && x11 && x17 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x9 && x13 && ~x21 && ~x10 && x22 && x14 && x11 && ~x17 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x9 && x13 && ~x21 && ~x10 && x22 && x14 && x11 && ~x17 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x9 && x13 && ~x21 && ~x10 && x22 && x14 && x11 && ~x17 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x9 && x13 && ~x21 && ~x10 && x22 && x14 && x11 && ~x17 && ~x6 )
						nx_state = s1;
					else if( ~x9 && x13 && ~x21 && ~x10 && x22 && x14 && ~x11 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x9 && x13 && ~x21 && ~x10 && x22 && ~x14 && x11 && x16 && x18 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x9 && x13 && ~x21 && ~x10 && x22 && ~x14 && x11 && x16 && ~x18 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x9 && x13 && ~x21 && ~x10 && x22 && ~x14 && x11 && x16 && ~x18 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x9 && x13 && ~x21 && ~x10 && x22 && ~x14 && x11 && x16 && ~x18 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x9 && x13 && ~x21 && ~x10 && x22 && ~x14 && x11 && x16 && ~x18 && ~x6 )
						nx_state = s1;
					else if( ~x9 && x13 && ~x21 && ~x10 && x22 && ~x14 && x11 && ~x16 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x9 && x13 && ~x21 && ~x10 && x22 && ~x14 && x11 && ~x16 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x9 && x13 && ~x21 && ~x10 && x22 && ~x14 && x11 && ~x16 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x9 && x13 && ~x21 && ~x10 && x22 && ~x14 && x11 && ~x16 && ~x6 )
						nx_state = s1;
					else if( ~x9 && x13 && ~x21 && ~x10 && x22 && ~x14 && ~x11 )
						begin
							y102 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x9 && x13 && ~x21 && ~x10 && ~x22 )
						begin
							y9 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y94 = 1'b1;	
							nx_state = s844;
						end
					else if( ~x9 && ~x13 )
						begin
							y9 = 1'b1;	y65 = 1'b1;	y84 = 1'b1;	
							y86 = 1'b1;	y91 = 1'b1;	
							nx_state = s1136;
						end
					else nx_state = s518;
				s519 : if( x69 && x17 && x13 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && x17 && ~x13 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && ~x17 && x7 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( x69 && ~x17 && ~x7 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x69 && x70 && x16 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( ~x69 && x70 && x16 && ~x6 && x8 && x19 && x62 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s320;
						end
					else if( ~x69 && x70 && x16 && ~x6 && x8 && x19 && ~x62 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( ~x69 && x70 && x16 && ~x6 && x8 && ~x19 && x26 && x62 && x5 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x69 && x70 && x16 && ~x6 && x8 && ~x19 && x26 && x62 && ~x5 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s733;
						end
					else if( ~x69 && x70 && x16 && ~x6 && x8 && ~x19 && x26 && ~x62 && x63 && x5 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x70 && x16 && ~x6 && x8 && ~x19 && x26 && ~x62 && x63 && ~x5 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x69 && x70 && x16 && ~x6 && x8 && ~x19 && x26 && ~x62 && ~x63 && x5 && x64 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s736;
						end
					else if( ~x69 && x70 && x16 && ~x6 && x8 && ~x19 && x26 && ~x62 && ~x63 && x5 && ~x64 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s737;
						end
					else if( ~x69 && x70 && x16 && ~x6 && x8 && ~x19 && x26 && ~x62 && ~x63 && ~x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( ~x69 && x70 && x16 && ~x6 && x8 && ~x19 && ~x26 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s738;
						end
					else if( ~x69 && x70 && x16 && ~x6 && ~x8 && x62 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( ~x69 && x70 && x16 && ~x6 && ~x8 && ~x62 && x63 )
						nx_state = s1;
					else if( ~x69 && x70 && x16 && ~x6 && ~x8 && ~x62 && ~x63 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x69 && x70 && ~x16 && x62 && x10 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s840;
						end
					else if( ~x69 && x70 && ~x16 && x62 && ~x10 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( ~x69 && x70 && ~x16 && ~x62 && x10 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && x70 && ~x16 && ~x62 && ~x10 && x63 )
						nx_state = s1;
					else if( ~x69 && x70 && ~x16 && ~x62 && ~x10 && ~x63 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x69 && ~x70 && x44 && x45 && x10 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x10 && x11 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s215;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x10 && ~x11 && x7 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x69 && ~x70 && x44 && x45 && ~x10 && ~x11 && ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x16 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x16 && ~x6 && x8 && x19 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x16 && ~x6 && x8 && ~x19 && x26 && x5 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x16 && ~x6 && x8 && ~x19 && x26 && ~x5 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x16 && ~x6 && x8 && ~x19 && ~x26 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s738;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && x16 && ~x6 && ~x8 )
						nx_state = s1;
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x16 && x10 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && ~x70 && x44 && ~x45 && ~x16 && ~x10 )
						nx_state = s1;
					else if( ~x69 && ~x70 && ~x44 && x10 && x7 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x69 && ~x70 && ~x44 && x10 && ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s215;
						end
					else nx_state = s519;
				s520 : if( 1'b1 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else nx_state = s520;
				s521 : if( 1'b1 )
						begin
							y10 = 1'b1;	
							nx_state = s405;
						end
					else nx_state = s521;
				s522 : if( x69 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x69 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x69 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x69 && x26 && x28 && x9 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( ~x69 && x26 && x28 && ~x9 && x23 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( ~x69 && x26 && x28 && ~x9 && ~x23 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x69 && x26 && ~x28 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else if( ~x69 && ~x26 && x27 && x35 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else if( ~x69 && ~x26 && x27 && ~x35 )
						nx_state = s1;
					else if( ~x69 && ~x26 && ~x27 && x28 && x2 && x24 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s1124;
						end
					else if( ~x69 && ~x26 && ~x27 && x28 && x2 && ~x24 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s995;
						end
					else if( ~x69 && ~x26 && ~x27 && x28 && ~x2 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && x49 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s922;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && x49 && ~x3 && x4 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s994;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && x49 && ~x3 && ~x4 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s995;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && ~x49 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else nx_state = s522;
				s523 : if( x22 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1100;
						end
					else if( ~x22 && x8 && x9 && x23 && x10 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y5 = 1'b1;	
							y22 = 1'b1;	y23 = 1'b1;	
							nx_state = s72;
						end
					else if( ~x22 && x8 && x9 && x23 && ~x10 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( ~x22 && x8 && x9 && ~x23 && x10 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y38 = 1'b1;	
							y46 = 1'b1;	
							nx_state = s741;
						end
					else if( ~x22 && x8 && x9 && ~x23 && ~x10 )
						begin
							y47 = 1'b1;	
							nx_state = s287;
						end
					else if( ~x22 && x8 && ~x9 && x23 && x10 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x22 && x8 && ~x9 && x23 && x10 && ~x13 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && x8 && ~x9 && x23 && x10 && ~x13 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && x8 && ~x9 && x23 && x10 && ~x13 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x22 && x8 && ~x9 && x23 && x10 && ~x13 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && x8 && ~x9 && x23 && x10 && ~x13 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x22 && x8 && ~x9 && x23 && ~x10 && x1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x22 && x8 && ~x9 && x23 && ~x10 && ~x1 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && x8 && ~x9 && x23 && ~x10 && ~x1 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && x8 && ~x9 && x23 && ~x10 && ~x1 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x22 && x8 && ~x9 && x23 && ~x10 && ~x1 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && x8 && ~x9 && x23 && ~x10 && ~x1 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x22 && x8 && ~x9 && ~x23 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y42 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s1042;
						end
					else if( ~x22 && ~x8 && x9 && x23 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x22 && ~x8 && x9 && ~x23 && x10 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y38 = 1'b1;	
							y40 = 1'b1;	y41 = 1'b1;	
							nx_state = s741;
						end
					else if( ~x22 && ~x8 && x9 && ~x23 && ~x10 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y38 = 1'b1;	
							y39 = 1'b1;	y41 = 1'b1;	
							nx_state = s741;
						end
					else if( ~x22 && ~x8 && ~x9 && x23 && x10 && x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x22 && ~x8 && ~x9 && x23 && x10 && ~x3 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && ~x8 && ~x9 && x23 && x10 && ~x3 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && ~x8 && ~x9 && x23 && x10 && ~x3 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x22 && ~x8 && ~x9 && x23 && x10 && ~x3 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && ~x8 && ~x9 && x23 && x10 && ~x3 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x22 && ~x8 && ~x9 && x23 && ~x10 && x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x22 && ~x8 && ~x9 && x23 && ~x10 && ~x15 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && ~x8 && ~x9 && x23 && ~x10 && ~x15 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && ~x8 && ~x9 && x23 && ~x10 && ~x15 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x22 && ~x8 && ~x9 && x23 && ~x10 && ~x15 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && ~x8 && ~x9 && x23 && ~x10 && ~x15 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x22 && ~x8 && ~x9 && ~x23 )
						begin
							y5 = 1'b1;	y35 = 1'b1;	y36 = 1'b1;	
							y38 = 1'b1;	y41 = 1'b1;	
							nx_state = s741;
						end
					else nx_state = s523;
				s524 : if( x22 )
						begin
							y10 = 1'b1;	
							nx_state = s766;
						end
					else if( ~x22 && x23 )
						begin
							y10 = 1'b1;	
							nx_state = s193;
						end
					else if( ~x22 && ~x23 )
						begin
							y10 = 1'b1;	
							nx_state = s405;
						end
					else nx_state = s524;
				s525 : if( x63 )
						begin
							y6 = 1'b1;	y11 = 1'b1;	y26 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1028;
						end
					else if( ~x63 && x66 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x66 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x66 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x63 && x66 && ~x9 )
						nx_state = s1;
					else if( ~x63 && ~x66 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else nx_state = s525;
				s526 : if( x63 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x63 && x66 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x66 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x66 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x63 && x66 && ~x9 )
						nx_state = s1;
					else if( ~x63 && ~x66 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x63 && ~x66 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x63 && ~x66 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x63 && ~x66 && ~x18 )
						nx_state = s1;
					else nx_state = s526;
				s527 : if( x13 )
						begin
							y46 = 1'b1;	
							nx_state = s531;
						end
					else if( ~x13 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x13 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x13 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x13 && ~x9 )
						nx_state = s1;
					else nx_state = s527;
				s528 : if( x63 && x65 )
						begin
							y54 = 1'b1;	
							nx_state = s772;
						end
					else if( x63 && ~x65 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x65 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x65 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x63 && ~x65 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x65 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x63 && x64 && x67 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( ~x63 && x64 && ~x67 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x64 && ~x67 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x64 && ~x67 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x63 && x64 && ~x67 && ~x9 )
						nx_state = s1;
					else if( ~x63 && ~x64 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x64 && x20 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x64 && x20 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x63 && ~x64 && ~x20 )
						nx_state = s1;
					else nx_state = s528;
				s529 : if( 1'b1 )
						begin
							y46 = 1'b1;	
							nx_state = s531;
						end
					else nx_state = s529;
				s530 : if( x70 && x63 && x9 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && x63 && ~x9 && x67 && x7 )
						nx_state = s1;
					else if( x70 && x63 && ~x9 && x67 && ~x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( x70 && x63 && ~x9 && ~x67 )
						nx_state = s530;
					else if( x70 && ~x63 && x64 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x63 && x64 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x70 && ~x63 && x64 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x63 && x64 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && x23 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && x9 && x10 && x11 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && x9 && x10 && ~x11 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && x9 && ~x10 && x13 && x14 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && x9 && ~x10 && x13 && ~x14 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && x9 && ~x10 && x13 && ~x14 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && x9 && ~x10 && x13 && ~x14 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && x9 && ~x10 && x13 && ~x14 && ~x20 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && x9 && ~x10 && ~x13 && x15 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && x9 && ~x10 && ~x13 && ~x15 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && x9 && ~x10 && ~x13 && ~x15 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && x9 && ~x10 && ~x13 && ~x15 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && x9 && ~x10 && ~x13 && ~x15 && ~x20 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && ~x9 && x16 && x17 && x18 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && ~x9 && x16 && x17 && ~x18 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && ~x9 && x16 && x17 && ~x18 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && ~x9 && x16 && x17 && ~x18 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && ~x9 && x16 && x17 && ~x18 && ~x20 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && ~x9 && x16 && ~x17 && x19 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && ~x9 && x16 && ~x17 && ~x19 && x20 && x21 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && ~x9 && x16 && ~x17 && ~x19 && x20 && ~x21 && x22 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && ~x9 && x16 && ~x17 && ~x19 && x20 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && ~x9 && x16 && ~x17 && ~x19 && ~x20 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x66 && x24 && ~x23 && ~x9 && ~x16 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x66 && ~x24 && x11 && x12 && x23 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x66 && ~x24 && x11 && x12 && ~x23 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x66 && ~x24 && x11 && ~x12 && x13 && x23 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x66 && ~x24 && x11 && ~x12 && x13 && ~x23 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x70 && ~x63 && ~x64 && x65 && x66 && ~x24 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && x66 && ~x24 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && ~x66 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && ~x63 && ~x64 && x65 && ~x66 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && ~x63 && ~x64 && x65 && ~x66 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && x65 && ~x66 && ~x15 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && ~x65 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x63 && ~x64 && ~x65 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x70 && ~x63 && ~x64 && ~x65 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( x70 && ~x63 && ~x64 && ~x65 && ~x17 )
						nx_state = s1;
					else if( ~x70 && x21 && x65 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( ~x70 && x21 && x65 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( ~x70 && x21 && x65 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x70 && x21 && x65 && ~x8 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x65 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && ~x21 && x65 && x23 && x22 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && x65 && x23 && x22 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && x65 && x23 && x22 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x65 && x23 && x22 && ~x8 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x65 && x23 && ~x22 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && x65 && x23 && ~x22 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && x65 && x23 && ~x22 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x65 && x23 && ~x22 && ~x9 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x65 && ~x23 && x8 && x22 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && x65 && ~x23 && x8 && x22 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && x65 && ~x23 && x8 && x22 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x65 && ~x23 && x8 && ~x22 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && x65 && ~x23 && x8 && ~x22 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && x65 && ~x23 && x8 && ~x22 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x65 && ~x23 && ~x8 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x65 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else nx_state = s530;
				s531 : if( x63 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x63 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x63 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x63 && ~x1 )
						nx_state = s1;
					else if( ~x63 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x63 && ~x9 )
						nx_state = s1;
					else nx_state = s531;
				s532 : if( x64 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x64 && x31 )
						begin
							y44 = 1'b1;	
							nx_state = s1138;
						end
					else if( ~x64 && ~x31 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else nx_state = s532;
				s533 : if( x63 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x63 && x65 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x65 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x65 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x63 && x65 && ~x15 )
						nx_state = s1;
					else if( ~x63 && ~x65 )
						nx_state = s1;
					else nx_state = s533;
				s534 : if( 1'b1 )
						begin
							y9 = 1'b1;	y21 = 1'b1;	y41 = 1'b1;	
							nx_state = s1139;
						end
					else nx_state = s534;
				s535 : if( x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( ~x21 )
						nx_state = s1;
					else nx_state = s535;
				s536 : if( 1'b1 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else nx_state = s536;
				s537 : if( 1'b1 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s1140;
						end
					else nx_state = s537;
				s538 : if( x17 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y22 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s722;
						end
					else if( ~x17 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x17 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x17 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x17 && ~x10 )
						nx_state = s1;
					else nx_state = s538;
				s539 : if( x9 && x21 && x20 )
						begin
							y15 = 1'b1;	
							nx_state = s1141;
						end
					else if( x9 && x21 && ~x20 )
						begin
							y15 = 1'b1;	
							nx_state = s1142;
						end
					else if( x9 && ~x21 && x20 )
						begin
							y15 = 1'b1;	
							nx_state = s1116;
						end
					else if( x9 && ~x21 && ~x20 )
						begin
							y15 = 1'b1;	
							nx_state = s356;
						end
					else if( ~x9 )
						begin
							y7 = 1'b1;	y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s467;
						end
					else nx_state = s539;
				s540 : if( x69 && x62 && x10 && x7 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x69 && x62 && x10 && ~x7 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( x69 && x62 && ~x10 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && ~x62 && x17 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && ~x62 && x17 && ~x13 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && ~x62 && ~x17 && x7 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x69 && ~x62 && ~x17 && ~x7 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( ~x69 && x16 && x15 && x37 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x16 && x15 && ~x37 && x5 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x69 && x16 && x15 && ~x37 && ~x5 && x6 && x2 && x31 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s931;
						end
					else if( ~x69 && x16 && x15 && ~x37 && ~x5 && x6 && x2 && ~x31 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x69 && x16 && x15 && ~x37 && ~x5 && x6 && ~x2 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x69 && x16 && x15 && ~x37 && ~x5 && ~x6 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s1045;
						end
					else if( ~x69 && x16 && ~x15 && x4 && x5 && x34 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && x16 && ~x15 && x4 && x5 && ~x34 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x69 && x16 && ~x15 && x4 && x5 && ~x34 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && x16 && ~x15 && x4 && ~x5 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && x16 && ~x15 && ~x4 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && ~x16 && x15 && x7 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s1045;
						end
					else if( ~x69 && ~x16 && x15 && ~x7 && x9 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s1045;
						end
					else if( ~x69 && ~x16 && x15 && ~x7 && ~x9 && x10 && x6 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s540;
						end
					else if( ~x69 && ~x16 && x15 && ~x7 && ~x9 && x10 && ~x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s446;
						end
					else if( ~x69 && ~x16 && x15 && ~x7 && ~x9 && ~x10 && x11 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && ~x16 && x15 && ~x7 && ~x9 && ~x10 && ~x11 )
						nx_state = s540;
					else if( ~x69 && ~x16 && ~x15 && x3 && x11 && x2 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s698;
						end
					else if( ~x69 && ~x16 && ~x15 && x3 && x11 && ~x2 )
						nx_state = s540;
					else if( ~x69 && ~x16 && ~x15 && x3 && ~x11 && x4 && x12 && x13 && x31 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s455;
						end
					else if( ~x69 && ~x16 && ~x15 && x3 && ~x11 && x4 && x12 && x13 && x31 && ~x2 )
						nx_state = s540;
					else if( ~x69 && ~x16 && ~x15 && x3 && ~x11 && x4 && x12 && x13 && ~x31 && x2 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && ~x16 && ~x15 && x3 && ~x11 && x4 && x12 && x13 && ~x31 && ~x2 )
						nx_state = s540;
					else if( ~x69 && ~x16 && ~x15 && x3 && ~x11 && x4 && x12 && ~x13 )
						nx_state = s540;
					else if( ~x69 && ~x16 && ~x15 && x3 && ~x11 && x4 && ~x12 )
						nx_state = s540;
					else if( ~x69 && ~x16 && ~x15 && x3 && ~x11 && ~x4 )
						nx_state = s540;
					else if( ~x69 && ~x16 && ~x15 && ~x3 && x4 && x34 && x11 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s456;
						end
					else if( ~x69 && ~x16 && ~x15 && ~x3 && x4 && x34 && ~x11 && x12 && x13 && x14 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && ~x16 && ~x15 && ~x3 && x4 && x34 && ~x11 && x12 && x13 && ~x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s326;
						end
					else if( ~x69 && ~x16 && ~x15 && ~x3 && x4 && x34 && ~x11 && x12 && ~x13 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x69 && ~x16 && ~x15 && ~x3 && x4 && x34 && ~x11 && ~x12 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x69 && ~x16 && ~x15 && ~x3 && x4 && ~x34 )
						nx_state = s540;
					else if( ~x69 && ~x16 && ~x15 && ~x3 && ~x4 && x6 && x34 && x5 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && ~x16 && ~x15 && ~x3 && ~x4 && x6 && x34 && ~x5 && x9 && x7 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && ~x16 && ~x15 && ~x3 && ~x4 && x6 && x34 && ~x5 && x9 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s931;
						end
					else if( ~x69 && ~x16 && ~x15 && ~x3 && ~x4 && x6 && x34 && ~x5 && ~x9 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s931;
						end
					else if( ~x69 && ~x16 && ~x15 && ~x3 && ~x4 && x6 && x34 && ~x5 && ~x9 && ~x7 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && ~x16 && ~x15 && ~x3 && ~x4 && x6 && ~x34 )
						nx_state = s540;
					else if( ~x69 && ~x16 && ~x15 && ~x3 && ~x4 && ~x6 && x7 && x34 && x5 && x8 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && ~x16 && ~x15 && ~x3 && ~x4 && ~x6 && x7 && x34 && x5 && ~x8 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s931;
						end
					else if( ~x69 && ~x16 && ~x15 && ~x3 && ~x4 && ~x6 && x7 && x34 && ~x5 && x10 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && ~x16 && ~x15 && ~x3 && ~x4 && ~x6 && x7 && x34 && ~x5 && ~x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s931;
						end
					else if( ~x69 && ~x16 && ~x15 && ~x3 && ~x4 && ~x6 && x7 && ~x34 )
						nx_state = s540;
					else if( ~x69 && ~x16 && ~x15 && ~x3 && ~x4 && ~x6 && ~x7 && x34 && x5 && x8 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s931;
						end
					else if( ~x69 && ~x16 && ~x15 && ~x3 && ~x4 && ~x6 && ~x7 && x34 && x5 && ~x8 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && ~x16 && ~x15 && ~x3 && ~x4 && ~x6 && ~x7 && x34 && ~x5 && x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s931;
						end
					else if( ~x69 && ~x16 && ~x15 && ~x3 && ~x4 && ~x6 && ~x7 && x34 && ~x5 && ~x10 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x69 && ~x16 && ~x15 && ~x3 && ~x4 && ~x6 && ~x7 && ~x34 )
						nx_state = s540;
					else nx_state = s540;
				s541 : if( x69 && x62 && x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( x69 && x62 && ~x6 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s542;
						end
					else if( x69 && ~x62 && x17 && x18 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x5 && x6 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x5 && ~x6 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && x17 && ~x18 && x14 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s45;
						end
					else if( x69 && ~x62 && x17 && ~x18 && ~x14 )
						nx_state = s1;
					else if( x69 && ~x62 && ~x17 && x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( x69 && ~x62 && ~x17 && ~x6 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s542;
						end
					else if( ~x69 && x17 && x18 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( ~x69 && x17 && x18 && ~x5 && x6 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x17 && x18 && ~x5 && ~x6 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x17 && ~x18 && x14 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s45;
						end
					else if( ~x69 && x17 && ~x18 && ~x14 && x15 && x16 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x69 && x17 && ~x18 && ~x14 && x15 && x16 && ~x5 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x69 && x17 && ~x18 && ~x14 && x15 && x16 && ~x5 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x69 && x17 && ~x18 && ~x14 && x15 && ~x16 && x1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && x17 && ~x18 && ~x14 && x15 && ~x16 && ~x1 )
						nx_state = s541;
					else if( ~x69 && x17 && ~x18 && ~x14 && ~x15 && x16 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && x17 && ~x18 && ~x14 && ~x15 && ~x16 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x69 && x17 && ~x18 && ~x14 && ~x15 && ~x16 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x17 && x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( ~x69 && ~x17 && ~x6 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s542;
						end
					else nx_state = s541;
				s542 : if( x69 && x62 && x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && x62 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( x69 && ~x62 && x17 && x18 && x6 && x9 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s540;
						end
					else if( x69 && ~x62 && x17 && x18 && x6 && ~x9 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s541;
						end
					else if( x69 && ~x62 && x17 && ~x18 && x10 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && ~x62 && x17 && ~x18 && ~x10 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s544;
						end
					else if( x69 && ~x62 && ~x17 && x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && ~x62 && ~x17 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( ~x69 && x63 && x40 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( ~x69 && x63 && ~x40 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s994;
						end
					else if( ~x69 && ~x63 && x64 && x9 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( ~x69 && ~x63 && x64 && ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( ~x69 && ~x63 && ~x64 && x17 && x18 && x6 && x9 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s546;
						end
					else if( ~x69 && ~x63 && ~x64 && x17 && x18 && x6 && ~x9 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( ~x69 && ~x63 && ~x64 && x17 && x18 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s541;
						end
					else if( ~x69 && ~x63 && ~x64 && x17 && ~x18 && x10 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && ~x63 && ~x64 && x17 && ~x18 && ~x10 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s544;
						end
					else if( ~x69 && ~x63 && ~x64 && ~x17 && x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( ~x69 && ~x63 && ~x64 && ~x17 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else nx_state = s542;
				s543 : if( x18 && x17 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x18 && x17 && ~x1 && x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x18 && x17 && ~x1 && ~x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x18 && ~x17 && x31 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x18 && ~x17 && ~x31 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s546;
						end
					else if( ~x18 && x17 && x7 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x18 && x17 && ~x7 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x18 && ~x17 && x19 && x15 && x16 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x18 && ~x17 && x19 && x15 && x16 && ~x5 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x18 && ~x17 && x19 && x15 && x16 && ~x5 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x18 && ~x17 && x19 && x15 && ~x16 && x1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x18 && ~x17 && x19 && x15 && ~x16 && ~x1 )
						nx_state = s543;
					else if( ~x18 && ~x17 && x19 && ~x15 && x16 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x18 && ~x17 && x19 && ~x15 && ~x16 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x18 && ~x17 && x19 && ~x15 && ~x16 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x18 && ~x17 && ~x19 && x40 && x32 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( ~x18 && ~x17 && ~x19 && x40 && ~x32 && x15 && x16 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x18 && ~x17 && ~x19 && x40 && ~x32 && x15 && x16 && ~x5 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x18 && ~x17 && ~x19 && x40 && ~x32 && x15 && x16 && ~x5 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x18 && ~x17 && ~x19 && x40 && ~x32 && x15 && ~x16 && x1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x18 && ~x17 && ~x19 && x40 && ~x32 && x15 && ~x16 && ~x1 )
						nx_state = s543;
					else if( ~x18 && ~x17 && ~x19 && x40 && ~x32 && ~x15 && x16 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x18 && ~x17 && ~x19 && x40 && ~x32 && ~x15 && ~x16 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x18 && ~x17 && ~x19 && x40 && ~x32 && ~x15 && ~x16 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x18 && ~x17 && ~x19 && ~x40 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else nx_state = s543;
				s544 : if( x69 && x62 && x9 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && x62 && ~x9 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x69 && ~x62 && x17 && x18 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x5 && x6 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x5 && ~x6 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && x17 && ~x18 && x2 )
						nx_state = s1;
					else if( x69 && ~x62 && x17 && ~x18 && ~x2 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s541;
						end
					else if( x69 && ~x62 && ~x17 && x9 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && ~x62 && ~x17 && ~x9 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x69 && x17 && x18 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( ~x69 && x17 && x18 && ~x5 && x6 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x17 && x18 && ~x5 && ~x6 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x17 && ~x18 && x39 && x15 && x16 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x69 && x17 && ~x18 && x39 && x15 && x16 && ~x5 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x69 && x17 && ~x18 && x39 && x15 && x16 && ~x5 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x69 && x17 && ~x18 && x39 && x15 && ~x16 && x1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && x17 && ~x18 && x39 && x15 && ~x16 && ~x1 )
						nx_state = s544;
					else if( ~x69 && x17 && ~x18 && x39 && ~x15 && x16 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && x17 && ~x18 && x39 && ~x15 && ~x16 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x69 && x17 && ~x18 && x39 && ~x15 && ~x16 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && x17 && ~x18 && ~x39 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s541;
						end
					else if( ~x69 && ~x17 && x9 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && ~x17 && ~x9 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else nx_state = s544;
				s545 : if( x69 && x62 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && ~x62 && x17 && x18 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x1 && x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x1 && ~x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && ~x62 && x17 && ~x18 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( x69 && ~x62 && x17 && ~x18 && ~x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s551;
						end
					else if( x69 && ~x62 && ~x17 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( ~x69 && x63 && x11 && x43 && x13 && x10 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x69 && x63 && x11 && x43 && x13 && ~x10 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x63 && x11 && x43 && x13 && ~x10 && ~x34 && x37 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x63 && x11 && x43 && x13 && ~x10 && ~x34 && ~x37 )
						nx_state = s545;
					else if( ~x69 && x63 && x11 && x43 && ~x13 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x63 && x11 && x43 && ~x13 && ~x34 && x37 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x63 && x11 && x43 && ~x13 && ~x34 && ~x37 )
						nx_state = s545;
					else if( ~x69 && x63 && x11 && ~x43 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x63 && x11 && ~x43 && ~x34 && x37 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x63 && x11 && ~x43 && ~x34 && ~x37 )
						nx_state = s545;
					else if( ~x69 && x63 && ~x11 && x12 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x63 && ~x11 && x12 && ~x34 && x37 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x63 && ~x11 && x12 && ~x34 && ~x37 )
						nx_state = s545;
					else if( ~x69 && x63 && ~x11 && ~x12 && x44 && x14 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x63 && ~x11 && ~x12 && x44 && x14 && ~x34 && x37 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x63 && ~x11 && ~x12 && x44 && x14 && ~x34 && ~x37 )
						nx_state = s545;
					else if( ~x69 && x63 && ~x11 && ~x12 && x44 && ~x14 && x41 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x63 && ~x11 && ~x12 && x44 && ~x14 && x41 && ~x32 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x63 && ~x11 && ~x12 && x44 && ~x14 && ~x41 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x63 && ~x11 && ~x12 && x44 && ~x14 && ~x41 && ~x34 && x37 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x63 && ~x11 && ~x12 && x44 && ~x14 && ~x41 && ~x34 && ~x37 )
						nx_state = s545;
					else if( ~x69 && x63 && ~x11 && ~x12 && ~x44 && x34 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x63 && ~x11 && ~x12 && ~x44 && ~x34 && x37 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x63 && ~x11 && ~x12 && ~x44 && ~x34 && ~x37 )
						nx_state = s545;
					else if( ~x69 && ~x63 && x64 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && ~x63 && ~x64 && x17 && x18 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( ~x69 && ~x63 && ~x64 && x17 && x18 && ~x1 && x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && ~x63 && ~x64 && x17 && x18 && ~x1 && ~x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x69 && ~x63 && ~x64 && x17 && ~x18 && x35 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( ~x69 && ~x63 && ~x64 && x17 && ~x18 && ~x35 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s551;
						end
					else if( ~x69 && ~x63 && ~x64 && ~x17 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else nx_state = s545;
				s546 : if( x17 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x17 && ~x13 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x17 && x7 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x17 && ~x7 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else nx_state = s546;
				s547 : if( x16 && x15 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s1143;
						end
					else if( x16 && ~x15 && x4 && x5 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s1143;
						end
					else if( x16 && ~x15 && x4 && ~x5 )
						begin
							y21 = 1'b1;	y27 = 1'b1;	
							nx_state = s930;
						end
					else if( x16 && ~x15 && ~x4 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s929;
						end
					else if( ~x16 && x15 && x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s929;
						end
					else if( ~x16 && x15 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x16 && ~x15 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s1143;
						end
					else nx_state = s547;
				s548 : if( x69 )
						begin
							y7 = 1'b1;	
							nx_state = s747;
						end
					else if( ~x69 && x16 && x15 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s929;
						end
					else if( ~x69 && x16 && ~x15 && x4 )
						begin
							y21 = 1'b1;	y27 = 1'b1;	
							nx_state = s930;
						end
					else if( ~x69 && x16 && ~x15 && ~x4 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s929;
						end
					else if( ~x69 && ~x16 && x15 && x12 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s1143;
						end
					else if( ~x69 && ~x16 && x15 && ~x12 )
						nx_state = s548;
					else if( ~x69 && ~x16 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s929;
						end
					else if( ~x69 && ~x16 && ~x15 && ~x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s326;
						end
					else nx_state = s548;
				s549 : if( x16 && x15 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( x16 && x15 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( x16 && ~x15 && x4 && x5 && x1 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( x16 && ~x15 && x4 && x5 && ~x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( x16 && ~x15 && x4 && ~x5 && x37 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s1143;
						end
					else if( x16 && ~x15 && x4 && ~x5 && ~x37 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( x16 && ~x15 && ~x4 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( x16 && ~x15 && ~x4 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x16 && x15 && x31 && x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s326;
						end
					else if( ~x16 && x15 && x31 && ~x2 )
						nx_state = s549;
					else if( ~x16 && x15 && ~x31 && x4 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x16 && x15 && ~x31 && x4 && ~x2 )
						nx_state = s549;
					else if( ~x16 && x15 && ~x31 && ~x4 && x37 && x2 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x16 && x15 && ~x31 && ~x4 && x37 && ~x2 )
						nx_state = s549;
					else if( ~x16 && x15 && ~x31 && ~x4 && ~x37 && x2 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x16 && x15 && ~x31 && ~x4 && ~x37 && ~x2 )
						nx_state = s549;
					else if( ~x16 && ~x15 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else nx_state = s549;
				s550 : if( x15 && x16 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( x15 && ~x16 && x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s931;
						end
					else if( x15 && ~x16 && ~x5 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( ~x15 && x16 && x4 && x5 && x1 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( ~x15 && x16 && x4 && x5 && ~x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x15 && x16 && x4 && ~x5 && x37 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s1143;
						end
					else if( ~x15 && x16 && x4 && ~x5 && ~x37 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x15 && x16 && ~x4 && x37 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s1143;
						end
					else if( ~x15 && x16 && ~x4 && ~x37 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x15 && ~x16 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else nx_state = s550;
				s551 : if( x69 && x62 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && ~x62 && x17 && x18 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x1 && x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x1 && ~x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && ~x62 && x17 && ~x18 && x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( x69 && ~x62 && x17 && ~x18 && ~x6 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s542;
						end
					else if( x69 && ~x62 && ~x17 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x69 && x17 && x18 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s42;
						end
					else if( ~x69 && x17 && x18 && ~x1 && x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x17 && x18 && ~x1 && ~x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x69 && x17 && ~x18 && x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( ~x69 && x17 && ~x18 && ~x6 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s542;
						end
					else if( ~x69 && ~x17 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else nx_state = s551;
				s552 : if( x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s557;
						end
					else if( ~x3 && x2 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s46;
						end
					else if( ~x3 && x2 && ~x1 )
						begin
							y3 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							nx_state = s460;
						end
					else if( ~x3 && ~x2 && x1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x3 && ~x2 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else nx_state = s552;
				s553 : if( x68 && x6 && x15 && x10 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s605;
						end
					else if( x68 && x6 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s600;
						end
					else if( x68 && x6 && x15 && x10 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s132;
						end
					else if( x68 && x6 && x15 && ~x10 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s777;
						end
					else if( x68 && x6 && x15 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	
							nx_state = s133;
						end
					else if( x68 && x6 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s132;
						end
					else if( x68 && x6 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s607;
						end
					else if( x68 && ~x6 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s132;
						end
					else if( ~x68 && x60 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s139;
						end
					else if( ~x68 && ~x60 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else nx_state = s553;
				s554 : if( x60 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s139;
						end
					else if( ~x60 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else nx_state = s554;
				s555 : if( 1'b1 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s139;
						end
					else nx_state = s555;
				s556 : if( x65 && x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x65 && x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x65 && x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x65 && x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x65 && x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x65 && x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x65 && ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x65 && ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x20 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x65 && ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x65 && ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x65 && ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x65 && ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else nx_state = s556;
				s557 : if( x3 && x2 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s46;
						end
					else if( x3 && x2 && ~x1 )
						begin
							y3 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							nx_state = s460;
						end
					else if( x3 && ~x2 && x1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s557;
						end
					else if( x3 && ~x2 && ~x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( ~x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else nx_state = s557;
				s558 : if( x22 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s592;
						end
					else if( ~x22 && x19 && x15 && x8 )
						begin
							y11 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x22 && x19 && x15 && ~x8 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s591;
						end
					else if( ~x22 && x19 && ~x15 && x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s126;
						end
					else if( ~x22 && x19 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x22 && ~x19 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s592;
						end
					else nx_state = s558;
				s559 : if( x60 && x61 && x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s117;
						end
					else if( x60 && x61 && ~x18 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( x60 && ~x61 )
						begin
							y11 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x60 && x61 )
						begin
							y11 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x60 && ~x61 && x62 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( ~x60 && ~x61 && ~x62 )
						begin
							y7 = 1'b1;	
							nx_state = s747;
						end
					else nx_state = s559;
				s560 : if( x64 && x62 )
						begin
							y1 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s1144;
						end
					else if( x64 && ~x62 && x66 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else if( x64 && ~x62 && ~x66 )
						begin
							y4 = 1'b1;	y62 = 1'b1;	y63 = 1'b1;	
							nx_state = s1145;
						end
					else if( ~x64 && x62 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y37 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s1146;
						end
					else if( ~x64 && ~x62 && x30 )
						begin
							y33 = 1'b1;	
							nx_state = s589;
						end
					else if( ~x64 && ~x62 && ~x30 && x31 )
						begin
							y47 = 1'b1;	y56 = 1'b1;	y61 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s1110;
						end
					else if( ~x64 && ~x62 && ~x30 && ~x31 )
						begin
							y47 = 1'b1;	y52 = 1'b1;	y61 = 1'b1;	
							y66 = 1'b1;	
							nx_state = s54;
						end
					else nx_state = s560;
				s561 : if( 1'b1 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else nx_state = s561;
				s562 : if( x62 && x64 )
						begin
							y1 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1122;
						end
					else if( x62 && ~x64 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y37 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s1147;
						end
					else if( ~x62 && x64 && x5 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s35;
						end
					else if( ~x62 && x64 && ~x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x62 && ~x64 && x30 )
						begin
							y47 = 1'b1;	y52 = 1'b1;	y61 = 1'b1;	
							y66 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x62 && ~x64 && ~x30 )
						begin
							y47 = 1'b1;	y50 = 1'b1;	y61 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s1148;
						end
					else nx_state = s562;
				s563 : if( x69 && x21 && x20 && x10 && x12 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x21 && x20 && x10 && x12 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x21 && x20 && x10 && x12 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && x21 && x20 && x10 && x12 && ~x17 )
						nx_state = s1;
					else if( x69 && x21 && x20 && x10 && ~x12 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x69 && x21 && x20 && ~x10 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x21 && x20 && ~x10 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x69 && x21 && x20 && ~x10 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && x21 && x20 && ~x10 && ~x17 )
						nx_state = s1;
					else if( x69 && x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x69 && x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x21 && x10 && x12 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x21 && x10 && x12 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x21 && x10 && x12 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x21 && x10 && x12 && ~x19 )
						nx_state = s1;
					else if( x69 && ~x21 && x10 && ~x12 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x69 && ~x21 && ~x10 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x21 && ~x10 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x69 && ~x21 && ~x10 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x69 && ~x21 && ~x10 && ~x19 )
						nx_state = s1;
					else if( ~x69 && x44 && x41 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && x44 && ~x41 )
						nx_state = s563;
					else if( ~x69 && ~x44 && x45 && x46 && x2 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && ~x44 && x45 && x46 && ~x2 )
						nx_state = s563;
					else if( ~x69 && ~x44 && x45 && ~x46 && x2 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x69 && ~x44 && x45 && ~x46 && ~x2 )
						nx_state = s563;
					else if( ~x69 && ~x44 && ~x45 && x2 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x69 && ~x44 && ~x45 && ~x2 )
						nx_state = s563;
					else nx_state = s563;
				s564 : if( x61 && x60 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x61 && x60 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x61 && x60 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x61 && x60 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x61 && ~x60 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x61 && ~x60 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x61 && ~x60 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x61 && ~x60 && x62 && ~x18 )
						nx_state = s1;
					else if( x61 && ~x60 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x61 && ~x60 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x61 && ~x60 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( x61 && ~x60 && ~x62 && ~x18 )
						nx_state = s118;
					else if( ~x61 && x60 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x61 && x60 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x61 && x60 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( ~x61 && x60 && ~x18 )
						nx_state = s118;
					else if( ~x61 && ~x60 && x62 && x19 && x15 && x12 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s491;
						end
					else if( ~x61 && ~x60 && x62 && x19 && x15 && x12 && ~x7 )
						begin
							y12 = 1'b1;	
							nx_state = s490;
						end
					else if( ~x61 && ~x60 && x62 && x19 && x15 && ~x12 && x7 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x61 && ~x60 && x62 && x19 && x15 && ~x12 && ~x7 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s566;
						end
					else if( ~x61 && ~x60 && x62 && x19 && ~x15 && x16 && x7 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s490;
						end
					else if( ~x61 && ~x60 && x62 && x19 && ~x15 && x16 && x7 && ~x12 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s565;
						end
					else if( ~x61 && ~x60 && x62 && x19 && ~x15 && x16 && ~x7 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s487;
						end
					else if( ~x61 && ~x60 && x62 && x19 && ~x15 && ~x16 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x61 && ~x60 && x62 && x19 && ~x15 && ~x16 && ~x7 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x61 && ~x60 && x62 && ~x19 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y23 = 1'b1;	
							nx_state = s993;
						end
					else if( ~x61 && ~x60 && ~x62 )
						nx_state = s47;
					else nx_state = s564;
				s565 : if( x65 && x61 && x60 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x65 && x61 && x60 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x65 && x61 && x60 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x65 && x61 && x60 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x65 && x61 && ~x60 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x65 && x61 && ~x60 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x65 && x61 && ~x60 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x65 && x61 && ~x60 && x62 && ~x18 )
						nx_state = s1;
					else if( x65 && x61 && ~x60 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( x65 && x61 && ~x60 && ~x62 && ~x18 )
						nx_state = s118;
					else if( x65 && ~x61 && x60 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x65 && ~x61 && x60 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x65 && ~x61 && x60 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( x65 && ~x61 && x60 && ~x18 )
						nx_state = s118;
					else if( x65 && ~x61 && ~x60 && x62 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s487;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 )
						nx_state = s47;
					else if( ~x65 && x21 && x10 && x5 && x16 && x15 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s1039;
						end
					else if( ~x65 && x21 && x10 && x5 && x16 && ~x15 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x65 && x21 && x10 && x5 && ~x16 && x17 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s680;
						end
					else if( ~x65 && x21 && x10 && x5 && ~x16 && ~x17 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s680;
						end
					else if( ~x65 && x21 && x10 && ~x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x65 && x21 && ~x10 && x16 && x5 && x15 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s680;
						end
					else if( ~x65 && x21 && ~x10 && x16 && x5 && ~x15 )
						begin
							y13 = 1'b1;	y16 = 1'b1;	
							nx_state = s335;
						end
					else if( ~x65 && x21 && ~x10 && x16 && ~x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && x14 && x13 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && x14 && ~x13 && x15 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && x14 && ~x13 && ~x15 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && x14 && ~x13 && ~x15 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && x14 && ~x13 && ~x15 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && x14 && ~x13 && ~x15 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && ~x14 && x15 && x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && ~x14 && x15 && ~x12 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && ~x14 && x15 && ~x12 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && ~x14 && x15 && ~x12 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && ~x14 && x15 && ~x12 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && ~x14 && ~x15 && x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && ~x14 && ~x15 && ~x11 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && ~x14 && ~x15 && ~x11 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && ~x14 && ~x15 && ~x11 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && ~x14 && ~x15 && ~x11 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x21 && ~x10 && ~x16 && ~x17 && x5 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && ~x17 && ~x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x65 && ~x21 && x22 && x17 && x18 && x10 && x15 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x65 && ~x21 && x22 && x17 && x18 && x10 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && x14 && x15 && x9 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s267;
						end
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && x14 && x15 && ~x9 && x7 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && x14 && x15 && ~x9 && ~x7 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && x14 && ~x15 && x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && x14 && ~x15 && ~x8 && x7 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && x14 && ~x15 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && ~x14 && x15 && x9 )
						begin
							y6 = 1'b1;	
							nx_state = s368;
						end
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && ~x14 && x15 && ~x9 && x8 && x7 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && ~x14 && x15 && ~x9 && x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && ~x14 && x15 && ~x9 && ~x8 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && ~x14 && ~x15 && x8 )
						begin
							y6 = 1'b1;	
							nx_state = s368;
						end
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && ~x14 && ~x15 && ~x8 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x65 && ~x21 && x22 && x17 && ~x18 && x14 && x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s852;
						end
					else if( ~x65 && ~x21 && x22 && x17 && ~x18 && x14 && ~x10 && x15 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s1149;
						end
					else if( ~x65 && ~x21 && x22 && x17 && ~x18 && x14 && ~x10 && ~x15 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x65 && ~x21 && x22 && x17 && ~x18 && ~x14 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x65 && ~x21 && x22 && x17 && ~x18 && ~x14 && ~x2 && x5 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s792;
						end
					else if( ~x65 && ~x21 && x22 && x17 && ~x18 && ~x14 && ~x2 && ~x5 && x15 && x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s336;
						end
					else if( ~x65 && ~x21 && x22 && x17 && ~x18 && ~x14 && ~x2 && ~x5 && x15 && ~x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s828;
						end
					else if( ~x65 && ~x21 && x22 && x17 && ~x18 && ~x14 && ~x2 && ~x5 && ~x15 && x10 )
						begin
							y2 = 1'b1;	y16 = 1'b1;	y24 = 1'b1;	
							nx_state = s270;
						end
					else if( ~x65 && ~x21 && x22 && x17 && ~x18 && ~x14 && ~x2 && ~x5 && ~x15 && ~x10 )
						begin
							y14 = 1'b1;	y16 = 1'b1;	
							nx_state = s492;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && x10 && x5 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s792;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && x10 && ~x5 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s336;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && x14 && x15 && x5 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s792;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && x14 && x15 && ~x5 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && x14 && ~x15 && x13 && x5 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s792;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && x14 && ~x15 && x13 && ~x5 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && x14 && ~x15 && ~x13 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && x14 && ~x15 && ~x13 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && x14 && ~x15 && ~x13 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && x14 && ~x15 && ~x13 && ~x7 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && x15 && x12 && x5 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s792;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && x15 && x12 && ~x5 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && x15 && ~x12 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && x15 && ~x12 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && x15 && ~x12 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && x15 && ~x12 && ~x7 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && ~x15 && x11 && x5 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s792;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && ~x15 && x11 && ~x5 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && ~x15 && ~x11 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && ~x15 && ~x11 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && ~x15 && ~x11 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && ~x15 && ~x11 && ~x7 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && ~x18 && x5 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && ~x18 && ~x5 && x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s336;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && ~x18 && ~x5 && ~x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s829;
						end
					else if( ~x65 && ~x21 && ~x22 )
						nx_state = s1;
					else nx_state = s565;
				s566 : if( x60 && x61 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x60 && ~x61 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x60 && ~x61 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x60 && ~x61 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( x60 && ~x61 && ~x18 )
						nx_state = s118;
					else if( ~x60 && x61 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x60 && x61 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x60 && x61 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( ~x60 && x61 && x62 && ~x18 )
						nx_state = s1;
					else if( ~x60 && x61 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x60 && x61 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x60 && x61 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s118;
					else if( ~x60 && x61 && ~x62 && ~x18 )
						nx_state = s118;
					else if( ~x60 && ~x61 )
						nx_state = s47;
					else nx_state = s566;
				s567 : if( x65 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s139;
						end
					else if( ~x65 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s361;
						end
					else nx_state = s567;
				s568 : if( x70 && x62 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x70 && ~x62 && x63 && x7 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x70 && ~x62 && x63 && ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x20 && x3 )
						begin
							y14 = 1'b1;	
							nx_state = s366;
						end
					else if( x70 && ~x62 && ~x63 && x64 && x20 && ~x3 )
						begin
							y11 = 1'b1;	
							nx_state = s271;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x20 && x21 && x3 )
						begin
							y33 = 1'b1;	
							nx_state = s1033;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x20 && x21 && ~x3 )
						begin
							y31 = 1'b1;	
							nx_state = s1053;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x20 && ~x21 && x3 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x20 && ~x21 && ~x3 )
						begin
							y31 = 1'b1;	
							nx_state = s1150;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && x31 )
						begin
							y47 = 1'b1;	y54 = 1'b1;	y61 = 1'b1;	
							y68 = 1'b1;	
							nx_state = s855;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 && ~x31 )
						begin
							y47 = 1'b1;	y53 = 1'b1;	y61 = 1'b1;	
							y72 = 1'b1;	
							nx_state = s856;
						end
					else if( ~x70 && x65 && x67 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s644;
						end
					else if( ~x70 && x65 && ~x67 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x70 && ~x65 && x21 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && ~x65 && x21 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && ~x65 && x21 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x70 && ~x65 && x21 && ~x3 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && x22 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && ~x22 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x70 && ~x65 && ~x21 && ~x22 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x70 && ~x65 && ~x21 && ~x22 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x70 && ~x65 && ~x21 && ~x22 && ~x8 )
						nx_state = s1;
					else nx_state = s568;
				s569 : if( x21 )
						nx_state = s1;
					else if( ~x21 && x22 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x21 && x22 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x21 && x22 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x21 && ~x22 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x21 && ~x22 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x8 )
						nx_state = s1;
					else nx_state = s569;
				s570 : if( x65 && x2 && x18 && x19 && x14 && x17 && x20 && x16 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x65 && x2 && x18 && x19 && x14 && x17 && x20 && ~x16 )
						begin
							y24 = 1'b1;	
							nx_state = s259;
						end
					else if( x65 && x2 && x18 && x19 && x14 && x17 && ~x20 && x16 )
						begin
							y13 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	y29 = 1'b1;	y30 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s859;
						end
					else if( x65 && x2 && x18 && x19 && x14 && x17 && ~x20 && ~x16 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x65 && x2 && x18 && x19 && x14 && ~x17 && x20 && x8 && x16 )
						begin
							y13 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	y29 = 1'b1;	y30 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s859;
						end
					else if( x65 && x2 && x18 && x19 && x14 && ~x17 && x20 && x8 && ~x16 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && x18 && x19 && x14 && ~x17 && x20 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && x18 && x19 && x14 && ~x17 && ~x20 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && x15 && x17 && x20 && x16 )
						begin
							y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && x15 && x17 && x20 && ~x16 )
						begin
							y4 = 1'b1;	y12 = 1'b1;	y27 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && x15 && x17 && ~x20 && x16 )
						begin
							y24 = 1'b1;	
							nx_state = s259;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && x15 && x17 && ~x20 && ~x16 )
						begin
							y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && x15 && ~x17 && x16 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && x15 && ~x17 && ~x16 && x13 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && x15 && ~x17 && ~x16 && ~x13 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && x15 && ~x17 && ~x16 && ~x13 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && x15 && ~x17 && ~x16 && ~x13 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && x18 && x19 && ~x14 && x15 && ~x17 && ~x16 && ~x13 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && x17 && x16 && x7 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && x17 && x16 && ~x7 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && x17 && x16 && ~x7 && x5 && ~x6 )
						nx_state = s1;
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && x17 && x16 && ~x7 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && x17 && ~x16 && x6 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && x17 && ~x16 && ~x6 && x5 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && x17 && ~x16 && ~x6 && x5 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && x17 && ~x16 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && ~x17 && x16 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && ~x17 && x16 && ~x12 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && ~x17 && x16 && ~x12 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && ~x17 && x16 && ~x12 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && ~x17 && x16 && ~x12 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && ~x17 && ~x16 && x11 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && ~x17 && ~x16 && ~x11 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && ~x17 && ~x16 && ~x11 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && ~x17 && ~x16 && ~x11 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && ~x17 && ~x16 && ~x11 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && x17 && x20 && x14 && x13 )
						begin
							y10 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s861;
						end
					else if( x65 && x2 && x18 && ~x19 && x17 && x20 && x14 && ~x13 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x65 && x2 && x18 && ~x19 && x17 && x20 && ~x14 && x13 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	y19 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s861;
						end
					else if( x65 && x2 && x18 && ~x19 && x17 && x20 && ~x14 && ~x13 && x6 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s168;
						end
					else if( x65 && x2 && x18 && ~x19 && x17 && x20 && ~x14 && ~x13 && ~x6 && x5 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && x18 && ~x19 && x17 && x20 && ~x14 && ~x13 && ~x6 && x5 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && x17 && x20 && ~x14 && ~x13 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && x17 && ~x20 && x15 && x14 )
						begin
							y10 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s861;
						end
					else if( x65 && x2 && x18 && ~x19 && x17 && ~x20 && x15 && ~x14 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s168;
						end
					else if( x65 && x2 && x18 && ~x19 && x17 && ~x20 && ~x15 && x14 )
						begin
							y15 = 1'b1;	y28 = 1'b1;	
							nx_state = s862;
						end
					else if( x65 && x2 && x18 && ~x19 && x17 && ~x20 && ~x15 && ~x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && x13 && x12 && x14 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && x13 && x12 && ~x14 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && x13 && x12 && ~x14 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && x13 && x12 && ~x14 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && x13 && x12 && ~x14 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && x13 && ~x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && ~x13 && x11 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && ~x13 && x11 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && ~x13 && x11 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && ~x13 && x11 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && ~x13 && ~x11 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && x15 && x12 && x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s806;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && x15 && x12 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && x15 && ~x12 && x14 && x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s806;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && x15 && ~x12 && x14 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && x15 && ~x12 && ~x14 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && x15 && ~x12 && ~x14 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && x15 && ~x12 && ~x14 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && x15 && ~x12 && ~x14 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && x14 && x13 && x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s806;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && x14 && x13 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && x14 && ~x13 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && x14 && ~x13 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && x14 && ~x13 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && x14 && ~x13 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && ~x14 && x11 && x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s806;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && ~x14 && x11 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && ~x14 && ~x11 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && ~x14 && ~x11 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && ~x14 && ~x11 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && ~x14 && ~x11 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && ~x18 && x17 && x19 && x15 && x14 && x20 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && x15 && x14 && ~x20 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && x15 && ~x14 && x16 && x20 && x13 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && x15 && ~x14 && x16 && x20 && ~x13 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	y32 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && x15 && ~x14 && x16 && ~x20 && x13 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && x15 && ~x14 && x16 && ~x20 && ~x13 )
						begin
							y4 = 1'b1;	y29 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && x15 && ~x14 && ~x16 && x20 )
						begin
							y4 = 1'b1;	y29 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && x15 && ~x14 && ~x16 && ~x20 && x4 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s860;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && x15 && ~x14 && ~x16 && ~x20 && ~x4 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && ~x15 && x14 && x16 && x20 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && ~x15 && x14 && x16 && ~x20 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && ~x15 && x14 && ~x16 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && ~x15 && ~x14 && x20 && x8 && x16 )
						begin
							y4 = 1'b1;	y18 = 1'b1;	y29 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && ~x15 && ~x14 && x20 && x8 && ~x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && ~x15 && ~x14 && x20 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && ~x15 && ~x14 && ~x20 && x8 && x16 )
						begin
							y4 = 1'b1;	y17 = 1'b1;	y29 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && ~x15 && ~x14 && ~x20 && x8 && ~x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	y21 = 1'b1;	y28 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && ~x15 && ~x14 && ~x20 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && x16 && x14 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	y21 = 1'b1;	y28 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && x16 && ~x14 && x15 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && x16 && ~x14 && x15 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && x16 && ~x14 && x15 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && x16 && ~x14 && x15 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && x16 && ~x14 && ~x15 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && ~x16 && x13 && x14 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	y21 = 1'b1;	y28 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && ~x16 && x13 && x14 && ~x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && ~x16 && x13 && ~x14 && x4 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && ~x16 && x13 && ~x14 && ~x4 )
						begin
							y4 = 1'b1;	y12 = 1'b1;	y27 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && ~x16 && ~x13 && x8 )
						begin
							y13 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	y29 = 1'b1;	y30 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s859;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && ~x16 && ~x13 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && x14 && x16 )
						begin
							y24 = 1'b1;	
							nx_state = s259;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && x14 && ~x16 && x15 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && x14 && ~x16 && x15 && ~x13 )
						begin
							y4 = 1'b1;	y12 = 1'b1;	y27 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && x14 && ~x16 && ~x15 )
						begin
							y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && ~x14 && x15 && x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && ~x14 && x15 && ~x16 && x8 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	y21 = 1'b1;	y28 = 1'b1;	
							nx_state = s863;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && ~x14 && x15 && ~x16 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && ~x14 && ~x15 && x8 && x16 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && ~x14 && ~x15 && x8 && x16 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && ~x14 && ~x15 && x8 && x16 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && ~x14 && ~x15 && x8 && x16 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && ~x14 && ~x15 && x8 && ~x16 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	y19 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s861;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && ~x14 && ~x15 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && x2 && ~x18 && ~x17 && x8 )
						begin
							y4 = 1'b1;	y18 = 1'b1;	
							nx_state = s234;
						end
					else if( x65 && x2 && ~x18 && ~x17 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s1151;
						end
					else if( x65 && ~x2 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x65 && x21 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x65 && x21 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x65 && x21 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x65 && ~x21 && x22 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x65 && ~x21 && x22 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x21 && ~x22 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x65 && ~x21 && ~x22 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x65 && ~x21 && ~x22 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x65 && ~x21 && ~x22 && ~x8 )
						nx_state = s1;
					else nx_state = s570;
				s571 : if( 1'b1 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s377;
						end
					else nx_state = s571;
				s572 : if( x70 && x10 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && ~x10 && x11 )
						begin
							y14 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s401;
						end
					else if( x70 && ~x10 && ~x11 )
						begin
							y10 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s402;
						end
					else if( ~x70 && x21 && x66 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x21 && x66 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x21 && x66 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x21 && x66 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x66 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && x21 && ~x66 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && x21 && ~x66 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x66 && ~x3 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x66 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x70 && ~x21 && x66 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x70 && ~x21 && x66 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x66 && ~x20 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x66 && x22 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x70 && ~x21 && ~x66 && x22 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x70 && ~x21 && ~x66 && x22 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x66 && x22 && ~x6 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x66 && ~x22 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x70 && ~x21 && ~x66 && ~x22 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x70 && ~x21 && ~x66 && ~x22 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x66 && ~x22 && ~x8 )
						nx_state = s1;
					else nx_state = s572;
				s573 : if( x21 )
						begin
							y18 = 1'b1;	
							nx_state = s981;
						end
					else if( ~x21 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x21 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x21 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x6 )
						nx_state = s1;
					else nx_state = s573;
				s574 : if( x21 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x21 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else nx_state = s574;
				s575 : if( x70 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x70 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x70 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x21 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && ~x21 && x22 && x5 && x18 && x17 && x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s379;
						end
					else if( ~x70 && ~x21 && x22 && x5 && x18 && x17 && ~x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s379;
						end
					else if( ~x70 && ~x21 && x22 && x5 && x18 && ~x17 && x12 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s380;
						end
					else if( ~x70 && ~x21 && x22 && x5 && x18 && ~x17 && ~x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s6;
						end
					else if( ~x70 && ~x21 && x22 && x5 && ~x18 && x19 && x12 && x17 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s379;
						end
					else if( ~x70 && ~x21 && x22 && x5 && ~x18 && x19 && x12 && ~x17 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s382;
						end
					else if( ~x70 && ~x21 && x22 && x5 && ~x18 && x19 && ~x12 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && ~x21 && x22 && x5 && ~x18 && ~x19 && x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s379;
						end
					else if( ~x70 && ~x21 && x22 && x5 && ~x18 && ~x19 && ~x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x70 && ~x21 && x22 && ~x5 )
						begin
							y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s378;
						end
					else if( ~x70 && ~x21 && ~x22 && x18 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x70 && ~x21 && ~x22 && x18 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x70 && ~x21 && ~x22 && x18 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 && x18 && ~x8 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 && ~x18 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else nx_state = s575;
				s576 : if( x21 && x19 && x18 && x17 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s574;
						end
					else if( x21 && x19 && x18 && x17 && ~x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s574;
						end
					else if( x21 && x19 && x18 && ~x17 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x21 && x19 && x18 && ~x17 && ~x12 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s377;
						end
					else if( x21 && x19 && ~x18 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s575;
						end
					else if( x21 && ~x19 && x9 && x20 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s574;
						end
					else if( x21 && ~x19 && x9 && x20 && ~x12 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s171;
						end
					else if( x21 && ~x19 && x9 && ~x20 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s573;
						end
					else if( x21 && ~x19 && x9 && ~x20 && ~x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s175;
						end
					else if( x21 && ~x19 && ~x9 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s575;
						end
					else if( ~x21 && x22 && x3 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s575;
						end
					else if( ~x21 && x22 && ~x3 && x5 && x18 && x17 && x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s379;
						end
					else if( ~x21 && x22 && ~x3 && x5 && x18 && x17 && ~x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s379;
						end
					else if( ~x21 && x22 && ~x3 && x5 && x18 && ~x17 && x12 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s380;
						end
					else if( ~x21 && x22 && ~x3 && x5 && x18 && ~x17 && ~x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s6;
						end
					else if( ~x21 && x22 && ~x3 && x5 && ~x18 && x19 && x12 && x17 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s379;
						end
					else if( ~x21 && x22 && ~x3 && x5 && ~x18 && x19 && x12 && ~x17 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s382;
						end
					else if( ~x21 && x22 && ~x3 && x5 && ~x18 && x19 && ~x12 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x21 && x22 && ~x3 && x5 && ~x18 && ~x19 && x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s379;
						end
					else if( ~x21 && x22 && ~x3 && x5 && ~x18 && ~x19 && ~x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x21 && x22 && ~x3 && ~x5 )
						begin
							y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s378;
						end
					else if( ~x21 && ~x22 && x18 && x15 )
						begin
							y8 = 1'b1;	y18 = 1'b1;	
							nx_state = s152;
						end
					else if( ~x21 && ~x22 && x18 && ~x15 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s6;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && x15 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && x15 && ~x5 )
						begin
							y3 = 1'b1;	
							nx_state = s835;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 )
						begin
							y4 = 1'b1;	y21 = 1'b1;	
							nx_state = s377;
						end
					else if( ~x21 && ~x22 && ~x18 && ~x19 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else nx_state = s576;
				s577 : if( x69 && x67 && x11 && x5 && x6 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x67 && x11 && x5 && ~x6 && x7 )
						nx_state = s1;
					else if( x69 && x67 && x11 && x5 && ~x6 && ~x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( x69 && x67 && x11 && ~x5 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x69 && x67 && x11 && ~x5 && ~x4 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s577;
						end
					else if( x69 && x67 && ~x11 && x4 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && x67 && ~x11 && ~x4 )
						nx_state = s577;
					else if( x69 && ~x67 && x10 && x4 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && ~x67 && x10 && ~x4 )
						nx_state = s577;
					else if( x69 && ~x67 && ~x10 && x5 && x6 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && ~x67 && ~x10 && x5 && ~x6 && x7 )
						nx_state = s1;
					else if( x69 && ~x67 && ~x10 && x5 && ~x6 && ~x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( x69 && ~x67 && ~x10 && ~x5 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x69 && ~x67 && ~x10 && ~x5 && ~x4 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s577;
						end
					else if( ~x69 && x5 && x6 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x69 && x5 && ~x6 && x7 )
						nx_state = s1;
					else if( ~x69 && x5 && ~x6 && ~x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( ~x69 && ~x5 && x4 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && ~x5 && ~x4 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s577;
						end
					else nx_state = s577;
				s578 : if( x45 && x46 && x12 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x45 && x46 && ~x12 )
						nx_state = s578;
					else if( x45 && ~x46 && x12 && x5 && x6 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x45 && ~x46 && x12 && x5 && ~x6 && x7 )
						nx_state = s1;
					else if( x45 && ~x46 && x12 && x5 && ~x6 && ~x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( x45 && ~x46 && x12 && ~x5 && x4 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x45 && ~x46 && x12 && ~x5 && ~x4 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s578;
						end
					else if( x45 && ~x46 && ~x12 && x4 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x45 && ~x46 && ~x12 && ~x4 )
						nx_state = s578;
					else if( ~x45 && x46 && x4 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x45 && x46 && ~x4 )
						nx_state = s578;
					else if( ~x45 && ~x46 && x10 && x4 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x45 && ~x46 && x10 && ~x4 )
						nx_state = s578;
					else if( ~x45 && ~x46 && ~x10 && x5 && x6 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x45 && ~x46 && ~x10 && x5 && ~x6 && x7 )
						nx_state = s1;
					else if( ~x45 && ~x46 && ~x10 && x5 && ~x6 && ~x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s399;
						end
					else if( ~x45 && ~x46 && ~x10 && ~x5 && x4 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x45 && ~x46 && ~x10 && ~x5 && ~x4 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s578;
						end
					else nx_state = s578;
				s579 : if( x69 && x21 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s829;
						end
					else if( x69 && ~x21 && x22 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x69 && ~x21 && ~x22 && x3 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s443;
						end
					else if( x69 && ~x21 && ~x22 && ~x3 && x8 && x16 && x15 && x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x21 && ~x22 && ~x3 && x8 && x16 && x15 && ~x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s828;
						end
					else if( x69 && ~x21 && ~x22 && ~x3 && x8 && x16 && ~x15 && x10 )
						begin
							y2 = 1'b1;	y16 = 1'b1;	y24 = 1'b1;	
							nx_state = s270;
						end
					else if( x69 && ~x21 && ~x22 && ~x3 && x8 && x16 && ~x15 && ~x10 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s267;
						end
					else if( x69 && ~x21 && ~x22 && ~x3 && x8 && ~x16 && x17 && x10 && x15 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x21 && ~x22 && ~x3 && x8 && ~x16 && x17 && x10 && ~x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s827;
						end
					else if( x69 && ~x21 && ~x22 && ~x3 && x8 && ~x16 && x17 && ~x10 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s149;
						end
					else if( x69 && ~x21 && ~x22 && ~x3 && x8 && ~x16 && ~x17 && x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s336;
						end
					else if( x69 && ~x21 && ~x22 && ~x3 && x8 && ~x16 && ~x17 && ~x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s829;
						end
					else if( x69 && ~x21 && ~x22 && ~x3 && ~x8 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s127;
						end
					else if( ~x69 && x15 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x69 && ~x15 )
						nx_state = s579;
					else nx_state = s579;
				s580 : if( 1'b1 )
						begin
							y13 = 1'b1;	
							nx_state = s763;
						end
					else nx_state = s580;
				s581 : if( 1'b1 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else nx_state = s581;
				s582 : if( 1'b1 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else nx_state = s582;
				s583 : if( 1'b1 )
						begin
							y1 = 1'b1;	y15 = 1'b1;	y37 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s1152;
						end
					else nx_state = s583;
				s584 : if( x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( ~x27 )
						nx_state = s1;
					else nx_state = s584;
				s585 : if( x36 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y26 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s1153;
						end
					else if( ~x36 && x38 && x39 && x41 && x42 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y40 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s1154;
						end
					else if( ~x36 && x38 && x39 && x41 && ~x42 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y40 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x36 && x38 && x39 && ~x41 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y37 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s939;
						end
					else if( ~x36 && x38 && ~x39 && x40 && x55 && x56 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x36 && x38 && ~x39 && x40 && x55 && ~x56 && x58 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( ~x36 && x38 && ~x39 && x40 && x55 && ~x56 && ~x58 && x59 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x36 && x38 && ~x39 && x40 && x55 && ~x56 && ~x58 && ~x59 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x36 && x38 && ~x39 && x40 && x55 && ~x56 && ~x58 && ~x59 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x36 && x38 && ~x39 && x40 && x55 && ~x56 && ~x58 && ~x59 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( ~x36 && x38 && ~x39 && x40 && x55 && ~x56 && ~x58 && ~x59 && ~x27 )
						nx_state = s1;
					else if( ~x36 && x38 && ~x39 && x40 && ~x55 && x54 && x57 && x28 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x36 && x38 && ~x39 && x40 && ~x55 && x54 && x57 && ~x28 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x36 && x38 && ~x39 && x40 && ~x55 && x54 && x57 && ~x28 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x36 && x38 && ~x39 && x40 && ~x55 && x54 && x57 && ~x28 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( ~x36 && x38 && ~x39 && x40 && ~x55 && x54 && x57 && ~x28 && ~x27 )
						nx_state = s1;
					else if( ~x36 && x38 && ~x39 && x40 && ~x55 && x54 && ~x57 && x29 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x36 && x38 && ~x39 && x40 && ~x55 && x54 && ~x57 && ~x29 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x36 && x38 && ~x39 && x40 && ~x55 && x54 && ~x57 && ~x29 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x36 && x38 && ~x39 && x40 && ~x55 && x54 && ~x57 && ~x29 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( ~x36 && x38 && ~x39 && x40 && ~x55 && x54 && ~x57 && ~x29 && ~x27 )
						nx_state = s1;
					else if( ~x36 && x38 && ~x39 && x40 && ~x55 && ~x54 && x53 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x36 && x38 && ~x39 && x40 && ~x55 && ~x54 && ~x53 )
						begin
							y30 = 1'b1;	
							nx_state = s291;
						end
					else if( ~x36 && x38 && ~x39 && ~x40 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y37 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s1155;
						end
					else if( ~x36 && ~x38 )
						begin
							y2 = 1'b1;	y35 = 1'b1;	y37 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s1156;
						end
					else nx_state = s585;
				s586 : if( x10 )
						begin
							y25 = 1'b1;	
							nx_state = s1157;
						end
					else if( ~x10 && x11 && x14 && x30 && x36 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x10 && x11 && x14 && x30 && ~x36 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x10 && x11 && x14 && ~x30 && x31 && x33 && x34 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x10 && x11 && x14 && ~x30 && x31 && x33 && ~x34 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x10 && x11 && x14 && ~x30 && x31 && x33 && ~x34 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x10 && x11 && x14 && ~x30 && x31 && x33 && ~x34 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( ~x10 && x11 && x14 && ~x30 && x31 && x33 && ~x34 && ~x27 )
						nx_state = s1;
					else if( ~x10 && x11 && x14 && ~x30 && x31 && ~x33 && x35 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x10 && x11 && x14 && ~x30 && x31 && ~x33 && ~x35 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x10 && x11 && x14 && ~x30 && x31 && ~x33 && ~x35 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x10 && x11 && x14 && ~x30 && x31 && ~x33 && ~x35 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( ~x10 && x11 && x14 && ~x30 && x31 && ~x33 && ~x35 && ~x27 )
						nx_state = s1;
					else if( ~x10 && x11 && x14 && ~x30 && ~x31 && x32 )
						begin
							y1 = 1'b1;	y22 = 1'b1;	y37 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s581;
						end
					else if( ~x10 && x11 && x14 && ~x30 && ~x31 && ~x32 )
						begin
							y1 = 1'b1;	y20 = 1'b1;	y37 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s582;
						end
					else if( ~x10 && x11 && ~x14 && x15 && x16 && x20 && x22 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x10 && x11 && ~x14 && x15 && x16 && x20 && ~x22 )
						begin
							y36 = 1'b1;	
							nx_state = s963;
						end
					else if( ~x10 && x11 && ~x14 && x15 && x16 && ~x20 && x21 )
						begin
							y38 = 1'b1;	
							nx_state = s845;
						end
					else if( ~x10 && x11 && ~x14 && x15 && x16 && ~x20 && ~x21 )
						begin
							y37 = 1'b1;	y39 = 1'b1;	y44 = 1'b1;	
							y47 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x10 && x11 && ~x14 && x15 && ~x16 && x17 && x19 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y41 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1158;
						end
					else if( ~x10 && x11 && ~x14 && x15 && ~x16 && x17 && ~x19 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y44 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x10 && x11 && ~x14 && x15 && ~x16 && ~x17 && x18 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y39 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x10 && x11 && ~x14 && x15 && ~x16 && ~x17 && ~x18 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x10 && x11 && ~x14 && ~x15 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	y37 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1159;
						end
					else if( ~x10 && ~x11 && x12 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	y37 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1159;
						end
					else if( ~x10 && ~x11 && ~x12 && x13 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	y37 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1159;
						end
					else if( ~x10 && ~x11 && ~x12 && ~x13 && x43 && x46 && x48 )
						begin
							y37 = 1'b1;	y39 = 1'b1;	y47 = 1'b1;	
							nx_state = s1160;
						end
					else if( ~x10 && ~x11 && ~x12 && ~x13 && x43 && x46 && ~x48 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y39 = 1'b1;	
							nx_state = s1161;
						end
					else if( ~x10 && ~x11 && ~x12 && ~x13 && x43 && ~x46 && x47 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y39 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s1162;
						end
					else if( ~x10 && ~x11 && ~x12 && ~x13 && x43 && ~x46 && ~x47 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y39 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s1163;
						end
					else if( ~x10 && ~x11 && ~x12 && ~x13 && ~x43 && x44 && x45 )
						begin
							y19 = 1'b1;	y37 = 1'b1;	y39 = 1'b1;	
							y43 = 1'b1;	y44 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x10 && ~x11 && ~x12 && ~x13 && ~x43 && x44 && ~x45 )
						begin
							y14 = 1'b1;	y18 = 1'b1;	y37 = 1'b1;	
							y39 = 1'b1;	y45 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x10 && ~x11 && ~x12 && ~x13 && ~x43 && ~x44 )
						begin
							y14 = 1'b1;	y31 = 1'b1;	y35 = 1'b1;	
							y37 = 1'b1;	y39 = 1'b1;	y45 = 1'b1;	
							nx_state = s584;
						end
					else nx_state = s586;
				s587 : if( 1'b1 )
						begin
							y65 = 1'b1;	y90 = 1'b1;	y92 = 1'b1;	
							y98 = 1'b1;	y99 = 1'b1;	
							nx_state = s516;
						end
					else nx_state = s587;
				s588 : if( x62 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s537;
						end
					else if( ~x62 && x63 && x14 )
						begin
							y29 = 1'b1;	
							nx_state = s1017;
						end
					else if( ~x62 && x63 && ~x14 )
						begin
							y28 = 1'b1;	y30 = 1'b1;	
							nx_state = s1164;
						end
					else if( ~x62 && ~x63 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else nx_state = s588;
				s589 : if( x63 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x63 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x63 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x63 && ~x1 )
						nx_state = s1;
					else if( ~x63 && x64 )
						begin
							y34 = 1'b1;	
							nx_state = s1165;
						end
					else if( ~x63 && ~x64 && x66 )
						begin
							y47 = 1'b1;	y51 = 1'b1;	y61 = 1'b1;	
							y68 = 1'b1;	
							nx_state = s1166;
						end
					else if( ~x63 && ~x64 && ~x66 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y45 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s672;
						end
					else nx_state = s589;
				s590 : if( x64 && x66 )
						begin
							y3 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s1167;
						end
					else if( x64 && ~x66 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s749;
						end
					else if( ~x64 )
						begin
							y47 = 1'b1;	y49 = 1'b1;	y58 = 1'b1;	
							y61 = 1'b1;	y68 = 1'b1;	
							nx_state = s831;
						end
					else nx_state = s590;
				s591 : if( x70 && x4 && x20 && x9 && x8 && x7 && x6 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x70 && x4 && x20 && x9 && x8 && x7 && ~x6 && x5 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x70 && x4 && x20 && x9 && x8 && x7 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x70 && x4 && x20 && x9 && x8 && ~x7 )
						nx_state = s1;
					else if( x70 && x4 && x20 && x9 && ~x8 && x10 )
						begin
							y21 = 1'b1;	y38 = 1'b1;	
							nx_state = s412;
						end
					else if( x70 && x4 && x20 && x9 && ~x8 && ~x10 )
						begin
							y22 = 1'b1;	y29 = 1'b1;	
							nx_state = s412;
						end
					else if( x70 && x4 && x20 && ~x9 && x8 && x10 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s415;
						end
					else if( x70 && x4 && x20 && ~x9 && x8 && ~x10 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s301;
						end
					else if( x70 && x4 && x20 && ~x9 && ~x8 && x10 && x11 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x70 && x4 && x20 && ~x9 && ~x8 && x10 && ~x11 && x7 && x6 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x70 && x4 && x20 && ~x9 && ~x8 && x10 && ~x11 && x7 && ~x6 && x5 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x70 && x4 && x20 && ~x9 && ~x8 && x10 && ~x11 && x7 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x70 && x4 && x20 && ~x9 && ~x8 && x10 && ~x11 && ~x7 )
						nx_state = s1;
					else if( x70 && x4 && x20 && ~x9 && ~x8 && ~x10 && x12 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x70 && x4 && x20 && ~x9 && ~x8 && ~x10 && ~x12 && x7 && x6 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x70 && x4 && x20 && ~x9 && ~x8 && ~x10 && ~x12 && x7 && ~x6 && x5 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x70 && x4 && x20 && ~x9 && ~x8 && ~x10 && ~x12 && x7 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x70 && x4 && x20 && ~x9 && ~x8 && ~x10 && ~x12 && ~x7 )
						nx_state = s1;
					else if( x70 && x4 && ~x20 && x21 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x70 && x4 && ~x20 && x21 && ~x5 )
						begin
							y27 = 1'b1;	
							nx_state = s1083;
						end
					else if( x70 && x4 && ~x20 && ~x21 && x10 )
						nx_state = s47;
					else if( x70 && x4 && ~x20 && ~x21 && ~x10 )
						begin
							y27 = 1'b1;	
							nx_state = s1083;
						end
					else if( x70 && ~x4 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x22 && ~x17 )
						nx_state = s1;
					else if( ~x70 && ~x22 && x18 && x13 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && ~x22 && x18 && x13 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && ~x22 && x18 && ~x13 && x12 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && ~x22 && x18 && ~x13 && x12 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x70 && ~x22 && ~x18 )
						nx_state = s1;
					else nx_state = s591;
				s592 : if( x67 && x22 && x15 && x8 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x67 && x22 && x15 && ~x8 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x67 && x22 && ~x15 && x16 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x67 && x22 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( x67 && ~x22 )
						begin
							y10 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x67 && x60 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( ~x67 && ~x60 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else nx_state = s592;
				s593 : if( x69 && x4 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s307;
						end
					else if( x69 && ~x4 && x42 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x69 && ~x4 && x42 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && ~x4 && x42 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( x69 && ~x4 && x42 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y28 = 1'b1;	
							nx_state = s299;
						end
					else if( x69 && ~x4 && ~x42 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s1040;
						end
					else if( ~x69 && x64 && x61 && x46 && x3 && x23 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s201;
						end
					else if( ~x69 && x64 && x61 && x46 && x3 && ~x23 )
						nx_state = s593;
					else if( ~x69 && x64 && x61 && x46 && ~x3 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( ~x69 && x64 && x61 && ~x46 && x2 && x23 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s201;
						end
					else if( ~x69 && x64 && x61 && ~x46 && x2 && ~x23 )
						nx_state = s593;
					else if( ~x69 && x64 && x61 && ~x46 && ~x2 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( ~x69 && x64 && ~x61 && x10 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( ~x69 && x64 && ~x61 && ~x10 && x11 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && x64 && ~x61 && ~x10 && x11 && ~x5 && x6 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x64 && ~x61 && ~x10 && x11 && ~x5 && ~x6 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && x64 && ~x61 && ~x10 && ~x11 && x1 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( ~x69 && x64 && ~x61 && ~x10 && ~x11 && ~x1 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && ~x64 && x14 && x44 && x3 && x23 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s201;
						end
					else if( ~x69 && ~x64 && x14 && x44 && x3 && ~x23 )
						nx_state = s593;
					else if( ~x69 && ~x64 && x14 && x44 && ~x3 )
						nx_state = s1;
					else if( ~x69 && ~x64 && x14 && ~x44 && x2 && x23 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s201;
						end
					else if( ~x69 && ~x64 && x14 && ~x44 && x2 && ~x23 )
						nx_state = s593;
					else if( ~x69 && ~x64 && x14 && ~x44 && ~x2 )
						nx_state = s1;
					else if( ~x69 && ~x64 && ~x14 && x10 )
						nx_state = s1;
					else if( ~x69 && ~x64 && ~x14 && ~x10 && x11 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x69 && ~x64 && ~x14 && ~x10 && x11 && ~x5 && x6 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && ~x64 && ~x14 && ~x10 && x11 && ~x5 && ~x6 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && ~x64 && ~x14 && ~x10 && ~x11 && x1 )
						nx_state = s1;
					else if( ~x69 && ~x64 && ~x14 && ~x10 && ~x11 && ~x1 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else nx_state = s593;
				s594 : if( x70 )
						nx_state = s1;
					else if( ~x70 && x66 && x16 && x17 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x66 && x16 && x17 && x8 && ~x10 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x66 && x16 && x17 && ~x8 && x9 && x10 )
						begin
							y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s572;
						end
					else if( ~x70 && x66 && x16 && x17 && ~x8 && x9 && ~x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y15 = 1'b1;	
							y18 = 1'b1;	y25 = 1'b1;	
							nx_state = s233;
						end
					else if( ~x70 && x66 && x16 && x17 && ~x8 && ~x9 && x21 && x10 && x14 )
						begin
							y6 = 1'b1;	
							nx_state = s368;
						end
					else if( ~x70 && x66 && x16 && x17 && ~x8 && ~x9 && x21 && x10 && ~x14 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x66 && x16 && x17 && ~x8 && ~x9 && x21 && x10 && ~x14 && x19 && ~x15 )
						nx_state = s1;
					else if( ~x70 && x66 && x16 && x17 && ~x8 && ~x9 && x21 && x10 && ~x14 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x66 && x16 && x17 && ~x8 && ~x9 && x21 && ~x10 && x15 )
						begin
							y6 = 1'b1;	
							nx_state = s368;
						end
					else if( ~x70 && x66 && x16 && x17 && ~x8 && ~x9 && x21 && ~x10 && ~x15 && x19 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x66 && x16 && x17 && ~x8 && ~x9 && x21 && ~x10 && ~x15 && x19 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x66 && x16 && x17 && ~x8 && ~x9 && x21 && ~x10 && ~x15 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x66 && x16 && x17 && ~x8 && ~x9 && ~x21 && x10 && x14 )
						begin
							y6 = 1'b1;	
							nx_state = s368;
						end
					else if( ~x70 && x66 && x16 && x17 && ~x8 && ~x9 && ~x21 && x10 && ~x14 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x70 && x66 && x16 && x17 && ~x8 && ~x9 && ~x21 && x10 && ~x14 && x20 && ~x15 )
						nx_state = s1;
					else if( ~x70 && x66 && x16 && x17 && ~x8 && ~x9 && ~x21 && x10 && ~x14 && ~x20 )
						nx_state = s1;
					else if( ~x70 && x66 && x16 && x17 && ~x8 && ~x9 && ~x21 && ~x10 && x15 )
						begin
							y6 = 1'b1;	
							nx_state = s368;
						end
					else if( ~x70 && x66 && x16 && x17 && ~x8 && ~x9 && ~x21 && ~x10 && ~x15 && x20 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x70 && x66 && x16 && x17 && ~x8 && ~x9 && ~x21 && ~x10 && ~x15 && x20 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x66 && x16 && x17 && ~x8 && ~x9 && ~x21 && ~x10 && ~x15 && ~x20 )
						nx_state = s1;
					else if( ~x70 && x66 && x16 && ~x17 && x9 && x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s224;
						end
					else if( ~x70 && x66 && x16 && ~x17 && x9 && ~x21 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && x66 && x16 && ~x17 && ~x9 && x8 && x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s224;
						end
					else if( ~x70 && x66 && x16 && ~x17 && ~x9 && x8 && ~x21 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x70 && x66 && x16 && ~x17 && ~x9 && ~x8 && x2 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x70 && x66 && x16 && ~x17 && ~x9 && ~x8 && ~x2 && x21 && x3 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x70 && x66 && x16 && ~x17 && ~x9 && ~x8 && ~x2 && x21 && ~x3 && x10 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && x66 && x16 && ~x17 && ~x9 && ~x8 && ~x2 && x21 && ~x3 && ~x10 )
						begin
							y4 = 1'b1;	y18 = 1'b1;	
							nx_state = s234;
						end
					else if( ~x70 && x66 && x16 && ~x17 && ~x9 && ~x8 && ~x2 && ~x21 && x3 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x66 && x16 && ~x17 && ~x9 && ~x8 && ~x2 && ~x21 && ~x3 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s233;
						end
					else if( ~x70 && x66 && x16 && ~x17 && ~x9 && ~x8 && ~x2 && ~x21 && ~x3 && ~x10 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x70 && x66 && ~x16 && x2 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && x10 && x11 )
						begin
							y7 = 1'b1;	y12 = 1'b1;	
							nx_state = s610;
						end
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && x10 && ~x11 && x9 )
						begin
							y7 = 1'b1;	y12 = 1'b1;	
							nx_state = s610;
						end
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && x10 && ~x11 && ~x9 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && x10 && ~x11 && ~x9 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && x10 && ~x11 && ~x9 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && x10 && ~x11 && ~x9 && x21 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && x10 && ~x11 && ~x9 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && x10 && ~x11 && ~x9 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && x10 && ~x11 && ~x9 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && x10 && ~x11 && ~x9 && ~x21 && ~x20 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && ~x10 && x9 && x13 )
						begin
							y7 = 1'b1;	y12 = 1'b1;	
							nx_state = s610;
						end
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && ~x10 && x9 && ~x13 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && ~x10 && x9 && ~x13 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && ~x10 && x9 && ~x13 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && ~x10 && x9 && ~x13 && x21 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && ~x10 && x9 && ~x13 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && ~x10 && x9 && ~x13 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && ~x10 && x9 && ~x13 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && ~x10 && x9 && ~x13 && ~x21 && ~x20 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && ~x10 && ~x9 && x12 )
						begin
							y7 = 1'b1;	y12 = 1'b1;	
							nx_state = s610;
						end
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && ~x10 && ~x9 && ~x12 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && ~x10 && ~x9 && ~x12 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && ~x10 && ~x9 && ~x12 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && ~x10 && ~x9 && ~x12 && x21 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && ~x10 && ~x9 && ~x12 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && ~x10 && ~x9 && ~x12 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && ~x10 && ~x9 && ~x12 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && ~x2 && x17 && ~x10 && ~x9 && ~x12 && ~x21 && ~x20 )
						nx_state = s1;
					else if( ~x70 && x66 && ~x16 && ~x2 && ~x17 && x3 && x21 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x70 && x66 && ~x16 && ~x2 && ~x17 && x3 && ~x21 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x70 && x66 && ~x16 && ~x2 && ~x17 && ~x3 )
						begin
							y17 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x70 && ~x66 && x21 && x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s384;
						end
					else if( ~x70 && ~x66 && x21 && ~x19 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s1168;
						end
					else if( ~x70 && ~x66 && ~x21 && x22 && x18 && x17 && x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s379;
						end
					else if( ~x70 && ~x66 && ~x21 && x22 && x18 && x17 && ~x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s379;
						end
					else if( ~x70 && ~x66 && ~x21 && x22 && x18 && ~x17 && x12 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s380;
						end
					else if( ~x70 && ~x66 && ~x21 && x22 && x18 && ~x17 && ~x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s6;
						end
					else if( ~x70 && ~x66 && ~x21 && x22 && ~x18 && x19 && x12 && x17 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s379;
						end
					else if( ~x70 && ~x66 && ~x21 && x22 && ~x18 && x19 && x12 && ~x17 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s382;
						end
					else if( ~x70 && ~x66 && ~x21 && x22 && ~x18 && x19 && ~x12 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && ~x66 && ~x21 && x22 && ~x18 && ~x19 && x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s379;
						end
					else if( ~x70 && ~x66 && ~x21 && x22 && ~x18 && ~x19 && ~x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x70 && ~x66 && ~x21 && ~x22 )
						nx_state = s1;
					else nx_state = s594;
				s595 : if( 1'b1 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s315;
						end
					else nx_state = s595;
				s596 : if( 1'b1 )
						begin
							y38 = 1'b1;	y40 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s596;
				s597 : if( 1'b1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y8 = 1'b1;	y9 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s1169;
						end
					else nx_state = s597;
				s598 : if( x10 )
						begin
							y62 = 1'b1;	
							nx_state = s1119;
						end
					else if( ~x10 && x11 && x4 && x5 && x3 && x12 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x10 && x11 && x4 && x5 && x3 && x12 && ~x8 && x7 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x10 && x11 && x4 && x5 && x3 && x12 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x10 && x11 && x4 && x5 && x3 && ~x12 )
						nx_state = s1;
					else if( ~x10 && x11 && x4 && x5 && ~x3 && x6 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x10 && x11 && x4 && x5 && ~x3 && x6 && ~x7 && x12 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x10 && x11 && x4 && x5 && ~x3 && x6 && ~x7 && x12 && ~x8 )
						nx_state = s1;
					else if( ~x10 && x11 && x4 && x5 && ~x3 && x6 && ~x7 && ~x12 )
						nx_state = s1;
					else if( ~x10 && x11 && x4 && x5 && ~x3 && ~x6 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x10 && x11 && x4 && x5 && ~x3 && ~x6 && ~x8 && x12 && x7 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x10 && x11 && x4 && x5 && ~x3 && ~x6 && ~x8 && x12 && ~x7 )
						nx_state = s1;
					else if( ~x10 && x11 && x4 && x5 && ~x3 && ~x6 && ~x8 && ~x12 )
						nx_state = s1;
					else if( ~x10 && x11 && x4 && ~x5 && x6 && x3 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x10 && x11 && x4 && ~x5 && x6 && ~x3 )
						begin
							y21 = 1'b1;	y38 = 1'b1;	
							nx_state = s412;
						end
					else if( ~x10 && x11 && x4 && ~x5 && ~x6 && x3 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x10 && x11 && x4 && ~x5 && ~x6 && ~x3 )
						begin
							y22 = 1'b1;	y29 = 1'b1;	
							nx_state = s412;
						end
					else if( ~x10 && x11 && ~x4 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x10 && ~x11 )
						begin
							y62 = 1'b1;	
							nx_state = s1120;
						end
					else nx_state = s598;
				s599 : if( 1'b1 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s858;
						end
					else nx_state = s599;
				s600 : if( x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x19 )
						nx_state = s1;
					else nx_state = s600;
				s601 : if( x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( ~x21 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else nx_state = s601;
				s602 : if( x70 )
						begin
							y17 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x70 && x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x21 && x20 && ~x17 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x19 )
						nx_state = s1;
					else nx_state = s602;
				s603 : if( x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x21 && ~x20 && x10 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x21 && ~x20 && ~x10 && x11 && x12 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && ~x20 && ~x10 && x11 && x12 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && ~x20 && ~x10 && x11 && x12 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x20 && ~x10 && x11 && x12 && ~x19 )
						nx_state = s1;
					else if( x21 && ~x20 && ~x10 && x11 && ~x12 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x21 && ~x20 && ~x10 && ~x11 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x19 )
						nx_state = s1;
					else nx_state = s603;
				s604 : if( x70 && x63 && x22 && x23 )
						begin
							y10 = 1'b1;	
							nx_state = s405;
						end
					else if( x70 && x63 && x22 && ~x23 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( x70 && x63 && ~x22 )
						begin
							y10 = 1'b1;	
							nx_state = s423;
						end
					else if( x70 && ~x63 )
						begin
							y48 = 1'b1;	
							nx_state = s1009;
						end
					else if( ~x70 && x20 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && ~x20 && x21 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && ~x20 && ~x21 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else nx_state = s604;
				s605 : if( x65 && x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x65 && x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x65 && x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x65 && x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x65 && x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x65 && x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x21 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x65 && x19 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s608;
						end
					else if( ~x65 && ~x19 && x20 && x15 && x10 && x11 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x65 && ~x19 && x20 && x15 && x10 && ~x11 && x12 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x65 && ~x19 && x20 && x15 && x10 && ~x11 && ~x12 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x65 && ~x19 && x20 && x15 && ~x10 && x12 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( ~x65 && ~x19 && x20 && x15 && ~x10 && x12 && ~x11 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x65 && ~x19 && x20 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( ~x65 && ~x19 && x20 && ~x15 && x16 && x10 && x12 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && ~x19 && x20 && ~x15 && x16 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s365;
						end
					else if( ~x65 && ~x19 && x20 && ~x15 && x16 && ~x10 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && ~x19 && x20 && ~x15 && ~x16 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s151;
						end
					else if( ~x65 && ~x19 && ~x20 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else nx_state = s605;
				s606 : if( x21 && x20 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s776;
						end
					else if( x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x19 )
						nx_state = s1;
					else nx_state = s606;
				s607 : if( x20 && x21 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x20 && x21 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x20 && x21 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x20 && x21 && ~x17 )
						nx_state = s1;
					else if( x20 && ~x21 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x20 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else nx_state = s607;
				s608 : if( x21 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && x20 && x15 && x10 && x11 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x21 && x20 && x15 && x10 && ~x11 && x12 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x21 && x20 && x15 && x10 && ~x11 && ~x12 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x21 && x20 && x15 && ~x10 && x12 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( ~x21 && x20 && x15 && ~x10 && x12 && ~x11 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x21 && x20 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( ~x21 && x20 && ~x15 && x16 && x10 && x12 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x21 && x20 && ~x15 && x16 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s365;
						end
					else if( ~x21 && x20 && ~x15 && x16 && ~x10 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x21 && x20 && ~x15 && ~x16 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s151;
						end
					else if( ~x21 && ~x20 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s229;
						end
					else nx_state = s608;
				s609 : if( x65 && x60 && x61 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s139;
						end
					else if( x65 && x60 && ~x61 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x65 && ~x60 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x65 && x23 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s1149;
						end
					else if( ~x65 && ~x23 && x19 )
						begin
							y14 = 1'b1;	
							nx_state = s366;
						end
					else if( ~x65 && ~x23 && ~x19 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else nx_state = s609;
				s610 : if( x66 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x66 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x66 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x66 && x21 && ~x19 )
						nx_state = s1;
					else if( x66 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( x66 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( x66 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x66 && ~x21 && ~x20 )
						nx_state = s1;
					else if( ~x66 && x20 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s668;
						end
					else if( ~x66 && ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x66 && ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x66 && ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x66 && ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x66 && ~x20 && ~x21 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else nx_state = s610;
				s611 : if( x26 && x28 && x7 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( x26 && x28 && ~x7 && x62 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s614;
						end
					else if( x26 && x28 && ~x7 && ~x62 && x63 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s995;
						end
					else if( x26 && x28 && ~x7 && ~x62 && ~x63 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else if( x26 && ~x28 )
						nx_state = s1;
					else if( ~x26 && x27 && x25 && x62 && x9 )
						nx_state = s611;
					else if( ~x26 && x27 && x25 && x62 && ~x9 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s614;
						end
					else if( ~x26 && x27 && x25 && ~x62 && x63 && x9 )
						nx_state = s611;
					else if( ~x26 && x27 && x25 && ~x62 && x63 && ~x9 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s995;
						end
					else if( ~x26 && x27 && x25 && ~x62 && ~x63 && x9 )
						nx_state = s611;
					else if( ~x26 && x27 && x25 && ~x62 && ~x63 && ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else if( ~x26 && x27 && ~x25 && x62 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( ~x26 && x27 && ~x25 && ~x62 && x63 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x26 && x27 && ~x25 && ~x62 && ~x63 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x26 && ~x27 && x62 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s942;
						end
					else if( ~x26 && ~x27 && ~x62 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else nx_state = s611;
				s612 : if( x26 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s943;
						end
					else if( ~x26 && x28 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s1170;
						end
					else if( ~x26 && x28 && ~x5 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s1171;
						end
					else if( ~x26 && ~x28 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s614;
						end
					else nx_state = s612;
				s613 : if( x28 && x7 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x28 && ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s405;
						end
					else if( ~x28 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else nx_state = s613;
				s614 : if( x26 && x21 )
						nx_state = s1;
					else if( x26 && ~x21 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s942;
						end
					else if( ~x26 && x27 )
						nx_state = s1;
					else if( ~x26 && ~x27 && x28 && x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( ~x26 && ~x27 && x28 && ~x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s613;
						end
					else if( ~x26 && ~x27 && ~x28 && x19 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s405;
						end
					else if( ~x26 && ~x27 && ~x28 && x19 && ~x24 )
						nx_state = s1;
					else if( ~x26 && ~x27 && ~x28 && ~x19 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s612;
						end
					else nx_state = s614;
				s615 : if( 1'b1 )
						begin
							y2 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s896;
						end
					else nx_state = s615;
				s616 : if( x63 && x11 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( x63 && x11 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( x63 && ~x11 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x63 && x64 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( ~x63 && ~x64 && x30 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s1172;
						end
					else if( ~x63 && ~x64 && x30 && ~x14 )
						begin
							y37 = 1'b1;	
							nx_state = s1173;
						end
					else if( ~x63 && ~x64 && ~x30 && x31 && x14 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x63 && ~x64 && ~x30 && x31 && ~x14 )
						begin
							y37 = 1'b1;	
							nx_state = s1174;
						end
					else if( ~x63 && ~x64 && ~x30 && ~x31 && x14 )
						begin
							y45 = 1'b1;	y46 = 1'b1;	y47 = 1'b1;	
							y49 = 1'b1;	y55 = 1'b1;	y58 = 1'b1;	
							y63 = 1'b1;	y70 = 1'b1;	
							nx_state = s1175;
						end
					else if( ~x63 && ~x64 && ~x30 && ~x31 && ~x14 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else nx_state = s616;
				s617 : if( x63 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1176;
						end
					else if( ~x63 && x31 && x30 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x63 && x31 && ~x30 )
						begin
							y35 = 1'b1;	
							nx_state = s718;
						end
					else if( ~x63 && ~x31 )
						begin
							y35 = 1'b1;	
							nx_state = s718;
						end
					else nx_state = s617;
				s618 : if( x19 && x18 )
						begin
							y2 = 1'b1;	
							nx_state = s708;
						end
					else if( x19 && ~x18 )
						begin
							y2 = 1'b1;	
							nx_state = s1177;
						end
					else if( ~x19 )
						begin
							y2 = 1'b1;	
							nx_state = s1111;
						end
					else nx_state = s618;
				s619 : if( 1'b1 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y23 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s619;
				s620 : if( 1'b1 )
						begin
							y3 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1178;
						end
					else nx_state = s620;
				s621 : if( x63 )
						begin
							y47 = 1'b1;	
							nx_state = s287;
						end
					else if( ~x63 && x67 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s712;
						end
					else if( ~x63 && ~x67 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1179;
						end
					else nx_state = s621;
				s622 : if( 1'b1 )
						begin
							y3 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s1180;
						end
					else nx_state = s622;
				s623 : if( 1'b1 )
						begin
							y3 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s327;
						end
					else nx_state = s623;
				s624 : if( 1'b1 )
						begin
							y3 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s223;
						end
					else nx_state = s624;
				s625 : if( x67 && x22 && x3 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x67 && x22 && x3 && x15 && ~x8 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( x67 && x22 && x3 && ~x15 && x16 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( x67 && x22 && x3 && ~x15 && ~x16 )
						begin
							y3 = 1'b1;	y11 = 1'b1;	
							nx_state = s89;
						end
					else if( x67 && x22 && ~x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( x67 && ~x22 && x23 && x18 && x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x67 && ~x22 && x23 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x67 && ~x22 && x23 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x67 && ~x22 && x23 && ~x18 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && x16 && x15 && x14 && x8 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x67 && ~x22 && ~x23 && x16 && x15 && x14 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x67 && ~x22 && ~x23 && x16 && x15 && ~x14 && x7 && x8 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x67 && ~x22 && ~x23 && x16 && x15 && ~x14 && x7 && ~x8 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s358;
						end
					else if( x67 && ~x22 && ~x23 && x16 && x15 && ~x14 && ~x7 && x8 && x12 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s426;
						end
					else if( x67 && ~x22 && ~x23 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && x18 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x67 && ~x22 && ~x23 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && x18 && ~x13 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && ~x18 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && x16 && x15 && ~x14 && ~x7 && ~x8 && x13 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s426;
						end
					else if( x67 && ~x22 && ~x23 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && x18 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x67 && ~x22 && ~x23 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && x18 && ~x12 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && ~x18 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && x8 && x9 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && x8 && x9 && ~x2 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && x8 && x9 && ~x2 && ~x3 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s486;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && x8 && ~x9 && x7 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && x8 && ~x9 && x7 && ~x2 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && x8 && ~x9 && x7 && ~x2 && ~x3 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s486;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && x8 && ~x9 && ~x7 && x18 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && x8 && ~x9 && ~x7 && x18 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && x8 && ~x9 && ~x7 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && x8 && ~x9 && ~x7 && ~x18 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && x7 && x11 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && x7 && x11 && ~x2 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && x7 && x11 && ~x2 && ~x3 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s486;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && x7 && ~x11 && x18 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && x7 && ~x11 && x18 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && x7 && ~x11 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && x7 && ~x11 && ~x18 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && ~x7 && x10 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && ~x7 && x10 && ~x2 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && ~x7 && x10 && ~x2 && ~x3 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s486;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && x18 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && x18 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x18 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && ~x16 && x15 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x67 && ~x22 && ~x23 && ~x16 && x15 && ~x7 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( x67 && ~x22 && ~x23 && ~x16 && x15 && ~x7 && ~x2 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x67 && ~x22 && ~x23 && ~x16 && x15 && ~x7 && ~x2 && ~x3 && x8 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y28 = 1'b1;	
							nx_state = s729;
						end
					else if( x67 && ~x22 && ~x23 && ~x16 && x15 && ~x7 && ~x2 && ~x3 && ~x8 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	
							nx_state = s486;
						end
					else if( x67 && ~x22 && ~x23 && ~x16 && ~x15 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else if( x67 && ~x22 && ~x23 && ~x16 && ~x15 && ~x2 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s458;
						end
					else if( x67 && ~x22 && ~x23 && ~x16 && ~x15 && ~x2 && ~x3 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s728;
						end
					else if( ~x67 && x21 && x20 && x15 && x10 && x11 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s600;
						end
					else if( ~x67 && x21 && x20 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s601;
						end
					else if( ~x67 && x21 && x20 && x15 && x10 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s776;
						end
					else if( ~x67 && x21 && x20 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( ~x67 && x21 && x20 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s602;
						end
					else if( ~x67 && x21 && x20 && ~x15 && x16 && x10 && x12 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( ~x67 && x21 && x20 && ~x15 && x16 && x10 && ~x12 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x67 && x21 && x20 && ~x15 && x16 && ~x10 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( ~x67 && x21 && x20 && ~x15 && ~x16 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x67 && x21 && ~x20 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s129;
						end
					else if( ~x67 && ~x21 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s825;
						end
					else if( ~x67 && ~x21 && ~x4 && x18 && x15 && x10 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x67 && ~x21 && ~x4 && x18 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s605;
						end
					else if( ~x67 && ~x21 && ~x4 && x18 && x15 && x10 && ~x11 && ~x12 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s606;
						end
					else if( ~x67 && ~x21 && ~x4 && x18 && x15 && ~x10 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( ~x67 && ~x21 && ~x4 && x18 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s600;
						end
					else if( ~x67 && ~x21 && ~x4 && x18 && ~x15 && x16 && x10 && x12 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( ~x67 && ~x21 && ~x4 && x18 && ~x15 && x16 && x10 && ~x12 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( ~x67 && ~x21 && ~x4 && x18 && ~x15 && x16 && ~x10 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( ~x67 && ~x21 && ~x4 && x18 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s607;
						end
					else if( ~x67 && ~x21 && ~x4 && ~x18 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s129;
						end
					else nx_state = s625;
				s626 : if( x3 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s644;
						end
					else if( ~x3 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s1181;
						end
					else nx_state = s626;
				s627 : if( x62 && x69 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( x62 && x69 && ~x2 && x1 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( x62 && x69 && ~x2 && ~x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x62 && ~x69 && x16 && x15 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s1182;
						end
					else if( x62 && ~x69 && x16 && ~x15 && x2 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else if( x62 && ~x69 && x16 && ~x15 && ~x2 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s901;
						end
					else if( x62 && ~x69 && x16 && ~x15 && ~x2 && ~x1 )
						begin
							y10 = 1'b1;	
							nx_state = s193;
						end
					else if( x62 && ~x69 && ~x16 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s1182;
						end
					else if( ~x62 && x69 && x16 && x15 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s1182;
						end
					else if( ~x62 && x69 && x16 && ~x15 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( ~x62 && x69 && x16 && ~x15 && ~x2 && x1 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x62 && x69 && x16 && ~x15 && ~x2 && ~x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x62 && x69 && ~x16 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s1182;
						end
					else if( ~x62 && ~x69 && x64 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s1182;
						end
					else if( ~x62 && ~x69 && ~x64 )
						begin
							y14 = 1'b1;	y31 = 1'b1;	
							nx_state = s1183;
						end
					else nx_state = s627;
				s628 : if( x69 && x62 && x4 )
						nx_state = s1;
					else if( x69 && x62 && ~x4 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( x69 && x62 && ~x4 && ~x2 && x1 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( x69 && x62 && ~x4 && ~x2 && ~x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x69 && ~x62 && x16 && x15 && x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s60;
						end
					else if( x69 && ~x62 && x16 && x15 && ~x5 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x69 && ~x62 && x16 && ~x15 && x4 )
						nx_state = s1;
					else if( x69 && ~x62 && x16 && ~x15 && ~x4 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( x69 && ~x62 && x16 && ~x15 && ~x4 && ~x2 && x1 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( x69 && ~x62 && x16 && ~x15 && ~x4 && ~x2 && ~x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x69 && ~x62 && ~x16 && x15 && x12 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( x69 && ~x62 && ~x16 && x15 && ~x12 )
						nx_state = s628;
					else if( x69 && ~x62 && ~x16 && ~x15 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s627;
						end
					else if( ~x69 && x64 && x40 && x46 && x3 && x23 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x69 && x64 && x40 && x46 && x3 && ~x23 )
						nx_state = s628;
					else if( ~x69 && x64 && x40 && x46 && ~x3 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && x64 && x40 && ~x46 && x2 && x23 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x69 && x64 && x40 && ~x46 && x2 && ~x23 )
						nx_state = s628;
					else if( ~x69 && x64 && x40 && ~x46 && ~x2 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && x64 && ~x40 && x10 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && x64 && ~x40 && ~x10 && x11 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x69 && x64 && ~x40 && ~x10 && x11 && ~x5 && x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && x64 && ~x40 && ~x10 && x11 && ~x5 && ~x6 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && x64 && ~x40 && ~x10 && ~x11 && x1 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && x64 && ~x40 && ~x10 && ~x11 && ~x1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && ~x64 && x44 && x46 && x42 && x23 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x69 && ~x64 && x44 && x46 && x42 && ~x23 )
						nx_state = s628;
					else if( ~x69 && ~x64 && x44 && x46 && ~x42 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x69 && ~x64 && x44 && ~x46 && x34 && x23 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x69 && ~x64 && x44 && ~x46 && x34 && ~x23 )
						nx_state = s628;
					else if( ~x69 && ~x64 && x44 && ~x46 && ~x34 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x69 && ~x64 && ~x44 && x10 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x69 && ~x64 && ~x44 && ~x10 && x11 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x69 && ~x64 && ~x44 && ~x10 && x11 && ~x5 && x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && ~x64 && ~x44 && ~x10 && x11 && ~x5 && ~x6 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else if( ~x69 && ~x64 && ~x44 && ~x10 && ~x11 && x36 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x69 && ~x64 && ~x44 && ~x10 && ~x11 && ~x36 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else nx_state = s628;
				s629 : if( x38 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x38 )
						nx_state = s629;
					else nx_state = s629;
				s630 : if( x63 && x41 && x12 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x63 && x41 && ~x12 && x32 && x2 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s818;
						end
					else if( x63 && x41 && ~x12 && x32 && ~x2 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x63 && x41 && ~x12 && ~x32 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( x63 && ~x41 && x42 && x32 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s882;
						end
					else if( x63 && ~x41 && x42 && ~x32 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( x63 && ~x41 && x42 && ~x32 && ~x3 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( x63 && ~x41 && ~x42 && x43 && x34 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s503;
						end
					else if( x63 && ~x41 && ~x42 && x43 && ~x34 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( x63 && ~x41 && ~x42 && ~x43 && x6 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x63 && ~x41 && ~x42 && ~x43 && ~x6 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x63 && x10 && x12 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x63 && x10 && ~x12 && x1 && x2 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x63 && x10 && ~x12 && x1 && ~x2 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x63 && x10 && ~x12 && ~x1 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x63 && ~x10 && x11 && x1 )
						begin
							y3 = 1'b1;	y13 = 1'b1;	y18 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s639;
						end
					else if( ~x63 && ~x10 && x11 && ~x1 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x63 && ~x10 && x11 && ~x1 && ~x3 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x63 && ~x10 && ~x11 && x12 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x63 && ~x10 && ~x11 && x12 && ~x3 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x63 && ~x10 && ~x11 && ~x12 && x6 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x63 && ~x10 && ~x11 && ~x12 && ~x6 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else nx_state = s630;
				s631 : if( x10 && x12 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( x10 && ~x12 && x1 && x34 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x10 && ~x12 && x1 && ~x34 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( x10 && ~x12 && ~x1 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x10 && x11 && x37 )
						begin
							y3 = 1'b1;	y13 = 1'b1;	y22 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s640;
						end
					else if( ~x10 && x11 && ~x37 && x41 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else if( ~x10 && x11 && ~x37 && ~x41 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x10 && ~x11 && x12 && x41 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x10 && ~x11 && x12 && ~x41 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x10 && ~x11 && ~x12 && x6 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x10 && ~x11 && ~x12 && ~x6 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else nx_state = s631;
				s632 : if( x70 && x63 && x64 && x55 && x10 && x43 && x23 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( x70 && x63 && x64 && x55 && x10 && x43 && ~x23 && x4 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( x70 && x63 && x64 && x55 && x10 && x43 && ~x23 && ~x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && x63 && x64 && x55 && x10 && ~x43 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( x70 && x63 && x64 && x55 && ~x10 && x1 && x22 )
						begin
							y10 = 1'b1;	y26 = 1'b1;	y37 = 1'b1;	
							nx_state = s1184;
						end
					else if( x70 && x63 && x64 && x55 && ~x10 && x1 && ~x22 && x2 && x3 && x42 )
						nx_state = s632;
					else if( x70 && x63 && x64 && x55 && ~x10 && x1 && ~x22 && x2 && x3 && ~x42 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( x70 && x63 && x64 && x55 && ~x10 && x1 && ~x22 && x2 && ~x3 && x11 && x5 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && x63 && x64 && x55 && ~x10 && x1 && ~x22 && x2 && ~x3 && x11 && ~x5 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( x70 && x63 && x64 && x55 && ~x10 && x1 && ~x22 && x2 && ~x3 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( x70 && x63 && x64 && x55 && ~x10 && x1 && ~x22 && ~x2 )
						begin
							y11 = 1'b1;	
							nx_state = s250;
						end
					else if( x70 && x63 && x64 && x55 && ~x10 && ~x1 && x42 && x35 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && x63 && x64 && x55 && ~x10 && ~x1 && x42 && ~x35 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( x70 && x63 && x64 && x55 && ~x10 && ~x1 && ~x42 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && x63 && x64 && ~x55 && x41 && x39 && x46 && x51 && x36 )
						nx_state = s632;
					else if( x70 && x63 && x64 && ~x55 && x41 && x39 && x46 && x51 && ~x36 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s906;
						end
					else if( x70 && x63 && x64 && ~x55 && x41 && x39 && x46 && ~x51 && x36 )
						nx_state = s632;
					else if( x70 && x63 && x64 && ~x55 && x41 && x39 && x46 && ~x51 && ~x36 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && x63 && x64 && ~x55 && x41 && x39 && ~x46 && x36 )
						nx_state = s632;
					else if( x70 && x63 && x64 && ~x55 && x41 && x39 && ~x46 && ~x36 )
						begin
							y11 = 1'b1;	
							nx_state = s250;
						end
					else if( x70 && x63 && x64 && ~x55 && x41 && ~x39 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s909;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x41 && x11 && x34 && x8 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s735;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x41 && x11 && x34 && ~x8 && x36 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s906;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x41 && x11 && x34 && ~x8 && ~x36 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x41 && x11 && ~x34 && x32 && x38 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s735;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x41 && x11 && ~x34 && x32 && ~x38 && x54 && x36 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s906;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x41 && x11 && ~x34 && x32 && ~x38 && x54 && ~x36 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x41 && x11 && ~x34 && x32 && ~x38 && ~x54 )
						begin
							y11 = 1'b1;	
							nx_state = s250;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x41 && x11 && ~x34 && ~x32 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x41 && ~x11 && x12 && x51 )
						begin
							y11 = 1'b1;	
							nx_state = s250;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x41 && ~x11 && x12 && ~x51 && x33 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x41 && ~x11 && x12 && ~x51 && ~x33 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x41 && ~x11 && ~x12 && x44 && x32 && x34 && x37 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x41 && ~x11 && ~x12 && x44 && x32 && x34 && ~x37 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x41 && ~x11 && ~x12 && x44 && x32 && ~x34 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x41 && ~x11 && ~x12 && x44 && ~x32 )
						begin
							y11 = 1'b1;	
							nx_state = s250;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x41 && ~x11 && ~x12 && ~x44 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && x63 && ~x64 && x15 && x22 && x2 && x33 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( x70 && x63 && ~x64 && x15 && x22 && x2 && ~x33 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && x63 && ~x64 && x15 && x22 && x2 && ~x33 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && x63 && ~x64 && x15 && x22 && ~x2 )
						nx_state = s1;
					else if( x70 && x63 && ~x64 && x15 && ~x22 && x31 )
						nx_state = s1;
					else if( x70 && x63 && ~x64 && x15 && ~x22 && ~x31 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && x63 && ~x64 && ~x15 && x46 && x3 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( x70 && x63 && ~x64 && ~x15 && x46 && x3 && ~x23 )
						nx_state = s632;
					else if( x70 && x63 && ~x64 && ~x15 && x46 && ~x3 )
						nx_state = s1;
					else if( x70 && x63 && ~x64 && ~x15 && ~x46 && x2 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( x70 && x63 && ~x64 && ~x15 && ~x46 && x2 && ~x23 )
						nx_state = s632;
					else if( x70 && x63 && ~x64 && ~x15 && ~x46 && ~x2 )
						nx_state = s1;
					else if( x70 && ~x63 && x10 && x40 && x12 && x23 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s93;
						end
					else if( x70 && ~x63 && x10 && x40 && x12 && ~x23 && x4 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x70 && ~x63 && x10 && x40 && x12 && ~x23 && ~x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && ~x63 && x10 && x40 && ~x12 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( x70 && ~x63 && x10 && ~x40 && x39 && x46 && x51 && x36 )
						nx_state = s632;
					else if( x70 && ~x63 && x10 && ~x40 && x39 && x46 && x51 && ~x36 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( x70 && ~x63 && x10 && ~x40 && x39 && x46 && ~x51 && x36 )
						nx_state = s632;
					else if( x70 && ~x63 && x10 && ~x40 && x39 && x46 && ~x51 && ~x36 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && ~x63 && x10 && ~x40 && x39 && ~x46 && x36 )
						nx_state = s632;
					else if( x70 && ~x63 && x10 && ~x40 && x39 && ~x46 && ~x36 )
						begin
							y11 = 1'b1;	
							nx_state = s250;
						end
					else if( x70 && ~x63 && x10 && ~x40 && ~x39 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( x70 && ~x63 && ~x10 && x40 && x1 && x22 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							nx_state = s869;
						end
					else if( x70 && ~x63 && ~x10 && x40 && x1 && ~x22 && x2 && x11 && x5 && x3 )
						nx_state = s632;
					else if( x70 && ~x63 && ~x10 && x40 && x1 && ~x22 && x2 && x11 && x5 && ~x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && ~x63 && ~x10 && x40 && x1 && ~x22 && x2 && x11 && ~x5 && x3 )
						nx_state = s632;
					else if( x70 && ~x63 && ~x10 && x40 && x1 && ~x22 && x2 && x11 && ~x5 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( x70 && ~x63 && ~x10 && x40 && x1 && ~x22 && x2 && ~x11 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && ~x10 && x40 && x1 && ~x22 && x2 && ~x11 && ~x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x70 && ~x63 && ~x10 && x40 && x1 && ~x22 && ~x2 )
						begin
							y11 = 1'b1;	
							nx_state = s250;
						end
					else if( x70 && ~x63 && ~x10 && x40 && ~x1 && x11 && x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && ~x63 && ~x10 && x40 && ~x1 && x11 && ~x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && ~x10 && x40 && ~x1 && ~x11 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && ~x63 && ~x10 && ~x40 && x11 && x34 && x8 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( x70 && ~x63 && ~x10 && ~x40 && x11 && x34 && ~x8 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( x70 && ~x63 && ~x10 && ~x40 && x11 && x34 && ~x8 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && ~x10 && ~x40 && x11 && ~x34 && x32 && x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( x70 && ~x63 && ~x10 && ~x40 && x11 && ~x34 && x32 && ~x7 && x45 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( x70 && ~x63 && ~x10 && ~x40 && x11 && ~x34 && x32 && ~x7 && x45 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && ~x10 && ~x40 && x11 && ~x34 && x32 && ~x7 && ~x45 )
						begin
							y11 = 1'b1;	
							nx_state = s250;
						end
					else if( x70 && ~x63 && ~x10 && ~x40 && x11 && ~x34 && ~x32 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( x70 && ~x63 && ~x10 && ~x40 && ~x11 && x12 && x20 )
						begin
							y11 = 1'b1;	
							nx_state = s250;
						end
					else if( x70 && ~x63 && ~x10 && ~x40 && ~x11 && x12 && ~x20 && x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && ~x63 && ~x10 && ~x40 && ~x11 && x12 && ~x20 && ~x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x70 && ~x63 && ~x10 && ~x40 && ~x11 && ~x12 && x13 && x1 && x3 && x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( x70 && ~x63 && ~x10 && ~x40 && ~x11 && ~x12 && x13 && x1 && x3 && ~x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && ~x10 && ~x40 && ~x11 && ~x12 && x13 && x1 && ~x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && ~x10 && ~x40 && ~x11 && ~x12 && x13 && ~x1 )
						begin
							y11 = 1'b1;	
							nx_state = s250;
						end
					else if( x70 && ~x63 && ~x10 && ~x40 && ~x11 && ~x12 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x70 && x22 && x2 && x20 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x70 && x22 && x2 && ~x20 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x70 && x22 && x2 && ~x20 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x70 && x22 && ~x2 )
						nx_state = s1;
					else if( ~x70 && ~x22 && x31 )
						nx_state = s1;
					else if( ~x70 && ~x22 && ~x31 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else nx_state = s632;
				s633 : if( x4 && x5 && x1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( x4 && x5 && ~x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( x4 && ~x5 && x2 && x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s634;
						end
					else if( x4 && ~x5 && x2 && ~x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( x4 && ~x5 && ~x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s477;
						end
					else if( ~x4 && x2 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s60;
						end
					else if( ~x4 && x2 && ~x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( ~x4 && ~x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s477;
						end
					else nx_state = s633;
				s634 : if( x69 && x62 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s686;
						end
					else if( x69 && x62 && ~x4 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s479;
						end
					else if( x69 && ~x62 && x15 && x16 )
						nx_state = s1;
					else if( x69 && ~x62 && x15 && ~x16 && x13 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s60;
						end
					else if( x69 && ~x62 && x15 && ~x16 && x13 && ~x4 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( x69 && ~x62 && x15 && ~x16 && ~x13 && x14 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( x69 && ~x62 && x15 && ~x16 && ~x13 && ~x14 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( x69 && ~x62 && x15 && ~x16 && ~x13 && ~x14 && ~x9 && x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( x69 && ~x62 && x15 && ~x16 && ~x13 && ~x14 && ~x9 && ~x7 && x8 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( x69 && ~x62 && x15 && ~x16 && ~x13 && ~x14 && ~x9 && ~x7 && ~x8 )
						nx_state = s634;
					else if( x69 && ~x62 && ~x15 && x16 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s686;
						end
					else if( x69 && ~x62 && ~x15 && x16 && ~x4 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( x69 && ~x62 && ~x15 && ~x16 )
						nx_state = s1;
					else if( ~x69 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s216;
						end
					else if( ~x69 && ~x15 && x13 && x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s997;
						end
					else if( ~x69 && ~x15 && x13 && ~x4 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1000;
						end
					else if( ~x69 && ~x15 && ~x13 && x14 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( ~x69 && ~x15 && ~x13 && ~x14 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( ~x69 && ~x15 && ~x13 && ~x14 && ~x9 && x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( ~x69 && ~x15 && ~x13 && ~x14 && ~x9 && ~x7 && x8 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( ~x69 && ~x15 && ~x13 && ~x14 && ~x9 && ~x7 && ~x8 )
						nx_state = s634;
					else nx_state = s634;
				s635 : if( x69 && x62 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( x69 && ~x62 && x15 && x16 && x5 && x1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( x69 && ~x62 && x15 && x16 && x5 && ~x1 && x2 && x3 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( x69 && ~x62 && x15 && x16 && x5 && ~x1 && x2 && x3 && ~x4 )
						nx_state = s1;
					else if( x69 && ~x62 && x15 && x16 && x5 && ~x1 && x2 && ~x3 )
						nx_state = s1;
					else if( x69 && ~x62 && x15 && x16 && x5 && ~x1 && ~x2 )
						nx_state = s1;
					else if( x69 && ~x62 && x15 && x16 && ~x5 && x6 )
						nx_state = s1;
					else if( x69 && ~x62 && x15 && x16 && ~x5 && ~x6 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s637;
						end
					else if( x69 && ~x62 && x15 && x16 && ~x5 && ~x6 && ~x1 && x2 && x3 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( x69 && ~x62 && x15 && x16 && ~x5 && ~x6 && ~x1 && x2 && x3 && ~x4 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x69 && ~x62 && x15 && x16 && ~x5 && ~x6 && ~x1 && x2 && ~x3 )
						nx_state = s1;
					else if( x69 && ~x62 && x15 && x16 && ~x5 && ~x6 && ~x1 && ~x2 )
						nx_state = s1;
					else if( x69 && ~x62 && x15 && ~x16 && x6 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x69 && ~x62 && x15 && ~x16 && ~x6 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s636;
						end
					else if( x69 && ~x62 && ~x15 && x16 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( x69 && ~x62 && ~x15 && ~x16 )
						nx_state = s1;
					else if( ~x69 && x26 && x8 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( ~x69 && x26 && x8 && ~x1 && x14 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( ~x69 && x26 && x8 && ~x1 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && x26 && ~x8 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s920;
						end
					else if( ~x69 && ~x26 && x28 )
						nx_state = s1;
					else if( ~x69 && ~x26 && ~x28 && x6 && x7 && x5 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s922;
						end
					else if( ~x69 && ~x26 && ~x28 && x6 && x7 && x5 && ~x3 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( ~x69 && ~x26 && ~x28 && x6 && x7 && x5 && ~x3 && ~x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else if( ~x69 && ~x26 && ~x28 && x6 && x7 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && ~x26 && ~x28 && x6 && ~x7 && x8 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s1185;
						end
					else if( ~x69 && ~x26 && ~x28 && x6 && ~x7 && ~x8 && x5 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s922;
						end
					else if( ~x69 && ~x26 && ~x28 && x6 && ~x7 && ~x8 && x5 && ~x3 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( ~x69 && ~x26 && ~x28 && x6 && ~x7 && ~x8 && x5 && ~x3 && ~x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else if( ~x69 && ~x26 && ~x28 && x6 && ~x7 && ~x8 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && ~x26 && ~x28 && ~x6 && x24 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s1185;
						end
					else if( ~x69 && ~x26 && ~x28 && ~x6 && ~x24 )
						nx_state = s1;
					else nx_state = s635;
				s636 : if( x62 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x62 && x16 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x62 && ~x16 && x15 && x8 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s638;
						end
					else if( ~x62 && ~x16 && x15 && ~x8 && x9 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s638;
						end
					else if( ~x62 && ~x16 && x15 && ~x8 && ~x9 && x10 && x6 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x62 && ~x16 && x15 && ~x8 && ~x9 && x10 && ~x6 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s636;
						end
					else if( ~x62 && ~x16 && x15 && ~x8 && ~x9 && ~x10 && x11 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s637;
						end
					else if( ~x62 && ~x16 && x15 && ~x8 && ~x9 && ~x10 && ~x11 )
						nx_state = s636;
					else if( ~x62 && ~x16 && ~x15 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else nx_state = s636;
				s637 : if( x15 && x16 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( x15 && ~x16 )
						nx_state = s1;
					else if( ~x15 && x16 && x4 && x5 && x1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( ~x15 && x16 && x4 && x5 && ~x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( ~x15 && x16 && x4 && ~x5 && x2 && x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s634;
						end
					else if( ~x15 && x16 && x4 && ~x5 && x2 && ~x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( ~x15 && x16 && x4 && ~x5 && ~x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s477;
						end
					else if( ~x15 && x16 && ~x4 && x2 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s60;
						end
					else if( ~x15 && x16 && ~x4 && x2 && ~x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( ~x15 && x16 && ~x4 && ~x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s477;
						end
					else if( ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s60;
						end
					else nx_state = s637;
				s638 : if( x69 && x16 && x15 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s686;
						end
					else if( x69 && x16 && ~x15 && x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( x69 && x16 && ~x15 && ~x3 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else if( x69 && ~x16 && x15 && x11 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s637;
						end
					else if( x69 && ~x16 && x15 && ~x11 && x10 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( x69 && ~x16 && x15 && ~x11 && ~x10 )
						nx_state = s638;
					else if( x69 && ~x16 && ~x15 )
						nx_state = s1;
					else if( ~x69 && x64 && x40 && x37 && x28 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x69 && x64 && x40 && x37 && ~x28 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && x64 && x40 && ~x37 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && x64 && ~x40 && x2 && x10 && x1 && x3 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x69 && x64 && ~x40 && x2 && x10 && x1 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x69 && x64 && ~x40 && x2 && x10 && x1 && ~x3 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x69 && x64 && ~x40 && x2 && x10 && ~x1 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s686;
						end
					else if( ~x69 && x64 && ~x40 && x2 && x10 && ~x1 && ~x9 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x69 && x64 && ~x40 && x2 && ~x10 )
						nx_state = s638;
					else if( ~x69 && x64 && ~x40 && ~x2 && x10 && x1 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && x64 && ~x40 && ~x2 && x10 && ~x1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s507;
						end
					else if( ~x69 && x64 && ~x40 && ~x2 && ~x10 )
						nx_state = s638;
					else if( ~x69 && ~x64 && x44 && x1 && x28 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x69 && ~x64 && x44 && x1 && ~x28 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && ~x64 && x44 && ~x1 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && ~x64 && ~x44 && x10 && x37 && x2 && x41 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x69 && ~x64 && ~x44 && x10 && x37 && x2 && ~x41 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x69 && ~x64 && ~x44 && x10 && x37 && x2 && ~x41 && ~x4 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s631;
						end
					else if( ~x69 && ~x64 && ~x44 && x10 && x37 && ~x2 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x69 && ~x64 && ~x44 && x10 && ~x37 && x2 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s686;
						end
					else if( ~x69 && ~x64 && ~x44 && x10 && ~x37 && x2 && ~x9 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x69 && ~x64 && ~x44 && x10 && ~x37 && ~x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s511;
						end
					else if( ~x69 && ~x64 && ~x44 && ~x10 )
						nx_state = s638;
					else nx_state = s638;
				s639 : if( x8 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s449;
						end
					else if( x8 && ~x1 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s1105;
						end
					else if( x8 && ~x1 && ~x4 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x8 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else nx_state = s639;
				s640 : if( x8 && x37 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s449;
						end
					else if( x8 && ~x37 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s1105;
						end
					else if( x8 && ~x37 && ~x4 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s508;
						end
					else if( ~x8 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else nx_state = s640;
				s641 : if( 1'b1 )
						begin
							y2 = 1'b1;	y37 = 1'b1;	y39 = 1'b1;	
							nx_state = s80;
						end
					else nx_state = s641;
				s642 : if( x64 && x3 )
						begin
							y14 = 1'b1;	
							nx_state = s5;
						end
					else if( x64 && ~x3 )
						begin
							y31 = 1'b1;	
							nx_state = s1186;
						end
					else if( ~x64 )
						begin
							y47 = 1'b1;	y56 = 1'b1;	y61 = 1'b1;	
							y72 = 1'b1;	
							nx_state = s1187;
						end
					else nx_state = s642;
				s643 : if( x21 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && x18 && x19 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && x22 && ~x23 && x18 && x19 && x15 && ~x17 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x21 && x22 && ~x23 && x18 && x19 && ~x15 && x16 && x17 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s296;
						end
					else if( ~x21 && x22 && ~x23 && x18 && x19 && ~x15 && x16 && ~x17 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y20 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s795;
						end
					else if( ~x21 && x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && x8 && x9 && x17 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && x8 && x9 && ~x17 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s724;
						end
					else if( ~x21 && x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && x8 && ~x9 && x10 && x17 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s724;
						end
					else if( ~x21 && x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && x8 && ~x9 && x10 && ~x17 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && x18 && ~x19 && x16 && x15 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( ~x21 && x22 && ~x23 && x18 && ~x19 && x16 && ~x15 && x17 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x21 && x22 && ~x23 && x18 && ~x19 && x16 && ~x15 && ~x17 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s796;
						end
					else if( ~x21 && x22 && ~x23 && x18 && ~x19 && ~x16 && x17 && x15 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( ~x21 && x22 && ~x23 && x18 && ~x19 && ~x16 && x17 && ~x15 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s797;
						end
					else if( ~x21 && x22 && ~x23 && x18 && ~x19 && ~x16 && ~x17 && x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x21 && x22 && ~x23 && x18 && ~x19 && ~x16 && ~x17 && ~x5 && x3 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s115;
						end
					else if( ~x21 && x22 && ~x23 && x18 && ~x19 && ~x16 && ~x17 && ~x5 && ~x3 && x15 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s795;
						end
					else if( ~x21 && x22 && ~x23 && x18 && ~x19 && ~x16 && ~x17 && ~x5 && ~x3 && ~x15 )
						begin
							y16 = 1'b1;	y20 = 1'b1;	
							nx_state = s795;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && x15 && x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && x15 && ~x5 && x3 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s115;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && x15 && ~x5 && ~x3 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s793;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && x16 && x14 && x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && x16 && x14 && ~x5 && x3 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s115;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && x16 && x14 && ~x5 && ~x3 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && x16 && ~x14 && x17 && x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && x16 && ~x14 && x17 && ~x5 && x3 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s115;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && x16 && ~x14 && x17 && ~x5 && ~x3 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && x16 && ~x14 && ~x17 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && ~x16 && x17 && x13 && x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && ~x16 && x17 && x13 && ~x5 && x3 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s115;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && ~x16 && x17 && x13 && ~x5 && ~x3 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && ~x16 && x17 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && ~x16 && ~x17 && x12 && x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && ~x16 && ~x17 && x12 && ~x5 && x3 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s115;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && ~x16 && ~x17 && x12 && ~x5 && ~x3 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && ~x16 && ~x17 && ~x12 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && ~x18 && ~x19 && x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && ~x19 && ~x5 && x3 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s115;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && ~x19 && ~x5 && ~x3 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( ~x21 && ~x22 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s301;
						end
					else nx_state = s643;
				s644 : if( 1'b1 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else nx_state = s644;
				s645 : if( x70 && x62 )
						begin
							y1 = 1'b1;	y12 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1188;
						end
					else if( x70 && ~x62 && x63 && x67 && x14 && x13 && x11 && x1 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x70 && ~x62 && x63 && x67 && x14 && x13 && x11 && ~x1 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && ~x62 && x63 && x67 && x14 && x13 && ~x11 && x10 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && ~x62 && x63 && x67 && x14 && x13 && ~x11 && ~x10 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && ~x62 && x63 && x67 && x14 && x13 && ~x11 && ~x10 && ~x3 && x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s65;
						end
					else if( x70 && ~x62 && x63 && x67 && x14 && x13 && ~x11 && ~x10 && ~x3 && ~x6 )
						nx_state = s645;
					else if( x70 && ~x62 && x63 && x67 && x14 && ~x13 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && ~x62 && x63 && x67 && x14 && ~x13 && ~x3 && x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s65;
						end
					else if( x70 && ~x62 && x63 && x67 && x14 && ~x13 && ~x3 && ~x6 )
						nx_state = s645;
					else if( x70 && ~x62 && x63 && x67 && ~x14 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && ~x62 && x63 && x67 && ~x14 && ~x3 && x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s65;
						end
					else if( x70 && ~x62 && x63 && x67 && ~x14 && ~x3 && ~x6 )
						nx_state = s645;
					else if( x70 && ~x62 && x63 && ~x67 && x15 && x13 && x14 && x10 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x70 && ~x62 && x63 && ~x67 && x15 && x13 && x14 && ~x10 && x1 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( x70 && ~x62 && x63 && ~x67 && x15 && x13 && x14 && ~x10 && ~x1 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && ~x62 && x63 && ~x67 && x15 && x13 && ~x14 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && ~x62 && x63 && ~x67 && x15 && x13 && ~x14 && ~x3 && x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s65;
						end
					else if( x70 && ~x62 && x63 && ~x67 && x15 && x13 && ~x14 && ~x3 && ~x6 )
						nx_state = s645;
					else if( x70 && ~x62 && x63 && ~x67 && x15 && ~x13 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && ~x62 && x63 && ~x67 && x15 && ~x13 && ~x3 && x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s65;
						end
					else if( x70 && ~x62 && x63 && ~x67 && x15 && ~x13 && ~x3 && ~x6 )
						nx_state = s645;
					else if( x70 && ~x62 && x63 && ~x67 && ~x15 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s69;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x15 && ~x3 && x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s65;
						end
					else if( x70 && ~x62 && x63 && ~x67 && ~x15 && ~x3 && ~x6 )
						nx_state = s645;
					else if( x70 && ~x62 && ~x63 && x64 && x21 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y62 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s1189;
						end
					else if( x70 && ~x62 && ~x63 && x64 && ~x21 )
						begin
							y4 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y78 = 1'b1;	
							nx_state = s1190;
						end
					else if( x70 && ~x62 && ~x63 && ~x64 )
						begin
							y47 = 1'b1;	y52 = 1'b1;	y61 = 1'b1;	
							y66 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x70 && x66 && x22 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( ~x70 && x66 && ~x22 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x70 && ~x66 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	
							nx_state = s594;
						end
					else nx_state = s645;
				s646 : if( 1'b1 )
						begin
							y46 = 1'b1;	
							nx_state = s775;
						end
					else nx_state = s646;
				s647 : if( 1'b1 )
						begin
							y13 = 1'b1;	
							nx_state = s450;
						end
					else nx_state = s647;
				s648 : if( x62 && x61 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s584;
						end
					else if( x62 && ~x61 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y37 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s989;
						end
					else if( ~x62 && x63 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s1191;
						end
					else if( ~x62 && ~x63 )
						begin
							y29 = 1'b1;	
							nx_state = s771;
						end
					else nx_state = s648;
				s649 : if( x62 && x65 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y15 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1192;
						end
					else if( x62 && ~x65 )
						begin
							y9 = 1'b1;	y21 = 1'b1;	y41 = 1'b1;	
							nx_state = s1193;
						end
					else if( ~x62 )
						begin
							y7 = 1'b1;	
							nx_state = s1194;
						end
					else nx_state = s649;
				s650 : if( x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x3 )
						nx_state = s1;
					else nx_state = s650;
				s651 : if( 1'b1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s653;
						end
					else nx_state = s651;
				s652 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s654;
						end
					else nx_state = s652;
				s653 : if( 1'b1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1195;
						end
					else nx_state = s653;
				s654 : if( x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( ~x22 )
						nx_state = s1;
					else nx_state = s654;
				s655 : if( x63 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x63 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x63 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( x63 && ~x22 )
						nx_state = s1;
					else if( ~x63 && x64 && x66 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x64 && x66 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x64 && x66 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x63 && x64 && x66 && ~x9 )
						nx_state = s1;
					else if( ~x63 && x64 && ~x66 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x63 && x64 && ~x66 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x63 && x64 && ~x66 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x63 && x64 && ~x66 && ~x18 )
						nx_state = s1;
					else if( ~x63 && ~x64 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s1196;
						end
					else nx_state = s655;
				s656 : if( x64 )
						begin
							y26 = 1'b1;	
							nx_state = s1197;
						end
					else if( ~x64 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s864;
						end
					else nx_state = s656;
				s657 : if( x22 )
						begin
							y10 = 1'b1;	
							nx_state = s1198;
						end
					else if( ~x22 )
						begin
							y10 = 1'b1;	
							nx_state = s841;
						end
					else nx_state = s657;
				s658 : if( x63 && x65 && x11 )
						begin
							y55 = 1'b1;	
							nx_state = s526;
						end
					else if( x63 && x65 && ~x11 )
						begin
							y54 = 1'b1;	
							nx_state = s772;
						end
					else if( x63 && ~x65 && x2 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x63 && ~x65 && ~x2 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x65 && ~x2 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x65 && ~x2 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x63 && ~x65 && ~x2 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x65 && ~x2 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x63 && x64 && x65 && x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x63 && x64 && x65 && x10 && ~x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x63 && x64 && x65 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x63 && x64 && x65 && ~x10 )
						nx_state = s1;
					else if( ~x63 && x64 && ~x65 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							nx_state = s1199;
						end
					else if( ~x63 && ~x64 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x64 && x20 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x64 && x20 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x63 && ~x64 && ~x20 )
						nx_state = s1;
					else nx_state = s658;
				s659 : if( x63 && x16 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s442;
						end
					else if( x63 && ~x16 )
						begin
							y3 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s520;
						end
					else if( ~x63 && x64 )
						begin
							y7 = 1'b1;	
							nx_state = s1200;
						end
					else if( ~x63 && ~x64 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else nx_state = s659;
				s660 : if( 1'b1 )
						begin
							y3 = 1'b1;	y28 = 1'b1;	y34 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s660;
				s661 : if( 1'b1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s1201;
						end
					else nx_state = s661;
				s662 : if( 1'b1 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y16 = 1'b1;	
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s1202;
						end
					else nx_state = s662;
				s663 : if( 1'b1 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else nx_state = s663;
				s664 : if( x21 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x21 && x22 && x23 && x15 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s805;
						end
					else if( ~x21 && x22 && x23 && ~x15 && x19 && x18 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s805;
						end
					else if( ~x21 && x22 && x23 && ~x15 && x19 && ~x18 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && x23 && ~x15 && x19 && ~x18 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && x23 && ~x15 && x19 && ~x18 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x15 && x19 && ~x18 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x15 && ~x19 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s805;
						end
					else if( ~x21 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 && x15 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s805;
						end
					else if( ~x21 && ~x22 && ~x23 && ~x15 && x19 && x18 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s805;
						end
					else if( ~x21 && ~x22 && ~x23 && ~x15 && x19 && ~x18 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x22 && ~x23 && ~x15 && x19 && ~x18 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x22 && ~x23 && ~x15 && x19 && ~x18 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 && ~x15 && x19 && ~x18 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 && ~x15 && ~x19 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s805;
						end
					else nx_state = s664;
				s665 : if( x70 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1203;
						end
					else if( ~x70 && x21 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( ~x70 && x21 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( ~x70 && x21 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x8 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x23 && x22 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && x23 && x22 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && x23 && x22 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x23 && x22 && ~x8 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x23 && ~x22 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && x23 && ~x22 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && x23 && ~x22 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x23 && ~x22 && ~x9 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x23 && x8 && x22 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && ~x23 && x8 && x22 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && ~x23 && x8 && x22 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x23 && x8 && ~x22 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && ~x23 && x8 && ~x22 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && ~x23 && x8 && ~x22 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x23 && ~x8 )
						nx_state = s1;
					else nx_state = s665;
				s666 : if( x70 && x5 )
						begin
							y52 = 1'b1;	y53 = 1'b1;	
							nx_state = s1204;
						end
					else if( x70 && ~x5 && x21 && x14 && x15 && x20 && x13 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1205;
						end
					else if( x70 && ~x5 && x21 && x14 && x15 && x20 && ~x13 )
						begin
							y54 = 1'b1;	
							nx_state = s281;
						end
					else if( x70 && ~x5 && x21 && x14 && x15 && ~x20 && x13 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else if( x70 && ~x5 && x21 && x14 && x15 && ~x20 && ~x13 && x18 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( x70 && ~x5 && x21 && x14 && x15 && ~x20 && ~x13 && ~x18 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x5 && x21 && x14 && x15 && ~x20 && ~x13 && ~x18 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x5 && x21 && x14 && x15 && ~x20 && ~x13 && ~x18 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x5 && x21 && x14 && x15 && ~x20 && ~x13 && ~x18 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x5 && x21 && x14 && ~x15 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s953;
						end
					else if( x70 && ~x5 && x21 && x14 && ~x15 && x20 && ~x13 )
						begin
							y29 = 1'b1;	
							nx_state = s771;
						end
					else if( x70 && ~x5 && x21 && x14 && ~x15 && ~x20 && x13 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( x70 && ~x5 && x21 && x14 && ~x15 && ~x20 && ~x13 && x19 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( x70 && ~x5 && x21 && x14 && ~x15 && ~x20 && ~x13 && ~x19 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x5 && x21 && x14 && ~x15 && ~x20 && ~x13 && ~x19 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x5 && x21 && x14 && ~x15 && ~x20 && ~x13 && ~x19 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x5 && x21 && x14 && ~x15 && ~x20 && ~x13 && ~x19 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x5 && x21 && ~x14 && x20 && x13 && x15 && x11 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else if( x70 && ~x5 && x21 && ~x14 && x20 && x13 && x15 && ~x11 && x10 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x5 && x21 && ~x14 && x20 && x13 && x15 && ~x11 && x10 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x5 && x21 && ~x14 && x20 && x13 && x15 && ~x11 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x5 && x21 && ~x14 && x20 && x13 && ~x15 && x12 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x70 && ~x5 && x21 && ~x14 && x20 && x13 && ~x15 && ~x12 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x5 && x21 && ~x14 && x20 && x13 && ~x15 && ~x12 && x10 && ~x11 )
						nx_state = s1;
					else if( x70 && ~x5 && x21 && ~x14 && x20 && x13 && ~x15 && ~x12 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x5 && x21 && ~x14 && x20 && ~x13 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x5 && x21 && ~x14 && x20 && ~x13 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x5 && x21 && ~x14 && x20 && ~x13 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x5 && x21 && ~x14 && x20 && ~x13 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x5 && x21 && ~x14 && ~x20 && x15 && x13 && x17 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( x70 && ~x5 && x21 && ~x14 && ~x20 && x15 && x13 && ~x17 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x5 && x21 && ~x14 && ~x20 && x15 && x13 && ~x17 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x5 && x21 && ~x14 && ~x20 && x15 && x13 && ~x17 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x5 && x21 && ~x14 && ~x20 && x15 && x13 && ~x17 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x5 && x21 && ~x14 && ~x20 && x15 && ~x13 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1207;
						end
					else if( x70 && ~x5 && x21 && ~x14 && ~x20 && ~x15 && x13 && x9 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( x70 && ~x5 && x21 && ~x14 && ~x20 && ~x15 && x13 && ~x9 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x5 && x21 && ~x14 && ~x20 && ~x15 && x13 && ~x9 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x70 && ~x5 && x21 && ~x14 && ~x20 && ~x15 && x13 && ~x9 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x5 && x21 && ~x14 && ~x20 && ~x15 && x13 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x5 && x21 && ~x14 && ~x20 && ~x15 && ~x13 && x7 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1208;
						end
					else if( x70 && ~x5 && x21 && ~x14 && ~x20 && ~x15 && ~x13 && ~x7 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1209;
						end
					else if( x70 && ~x5 && ~x21 && x7 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1208;
						end
					else if( x70 && ~x5 && ~x21 && ~x7 && x20 && x14 && x15 && x13 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y22 = 1'b1;	
							y32 = 1'b1;	y33 = 1'b1;	
							nx_state = s949;
						end
					else if( x70 && ~x5 && ~x21 && ~x7 && x20 && x14 && x15 && ~x13 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							nx_state = s1210;
						end
					else if( x70 && ~x5 && ~x21 && ~x7 && x20 && x14 && ~x15 && x13 )
						begin
							y6 = 1'b1;	y17 = 1'b1;	y34 = 1'b1;	
							nx_state = s226;
						end
					else if( x70 && ~x5 && ~x21 && ~x7 && x20 && x14 && ~x15 && ~x13 )
						begin
							y54 = 1'b1;	
							nx_state = s772;
						end
					else if( x70 && ~x5 && ~x21 && ~x7 && x20 && ~x14 && x15 && x13 )
						begin
							y6 = 1'b1;	y17 = 1'b1;	y34 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s1211;
						end
					else if( x70 && ~x5 && ~x21 && ~x7 && x20 && ~x14 && x15 && ~x13 )
						begin
							y6 = 1'b1;	y17 = 1'b1;	y46 = 1'b1;	
							y47 = 1'b1;	
							nx_state = s1212;
						end
					else if( x70 && ~x5 && ~x21 && ~x7 && x20 && ~x14 && ~x15 && x13 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							nx_state = s1213;
						end
					else if( x70 && ~x5 && ~x21 && ~x7 && x20 && ~x14 && ~x15 && ~x13 )
						begin
							y7 = 1'b1;	y39 = 1'b1;	y44 = 1'b1;	
							y49 = 1'b1;	
							nx_state = s1214;
						end
					else if( x70 && ~x5 && ~x21 && ~x7 && ~x20 && x13 )
						begin
							y6 = 1'b1;	y17 = 1'b1;	y34 = 1'b1;	
							nx_state = s226;
						end
					else if( x70 && ~x5 && ~x21 && ~x7 && ~x20 && ~x13 && x14 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y22 = 1'b1;	
							y32 = 1'b1;	y33 = 1'b1;	
							nx_state = s949;
						end
					else if( x70 && ~x5 && ~x21 && ~x7 && ~x20 && ~x13 && ~x14 )
						begin
							y6 = 1'b1;	y17 = 1'b1;	y34 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s1211;
						end
					else if( ~x70 && x21 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( ~x70 && ~x21 && x22 && x23 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x70 && ~x21 && x22 && x23 && ~x12 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && x22 && x23 && ~x12 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && x22 && x23 && ~x12 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x22 && x23 && ~x12 && ~x8 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x22 && ~x23 )
						begin
							y14 = 1'b1;	y19 = 1'b1;	
							nx_state = s723;
						end
					else if( ~x70 && ~x21 && ~x22 && x23 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && ~x22 && x23 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x70 && ~x21 && ~x22 && x23 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 && x23 && ~x9 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 && ~x23 )
						begin
							y6 = 1'b1;	y19 = 1'b1;	
							nx_state = s682;
						end
					else nx_state = s666;
				s667 : if( 1'b1 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else nx_state = s667;
				s668 : if( x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x20 && ~x18 )
						nx_state = s1;
					else if( ~x20 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else nx_state = s668;
				s669 : if( x69 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s670;
						end
					else if( ~x69 && x15 && x32 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s998;
						end
					else if( ~x69 && x15 && ~x32 )
						begin
							y11 = 1'b1;	
							nx_state = s248;
						end
					else if( ~x69 && ~x15 )
						begin
							y11 = 1'b1;	
							nx_state = s248;
						end
					else nx_state = s669;
				s670 : if( x69 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s691;
						end
					else if( ~x69 && x63 && x46 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x69 && x63 && ~x46 && x43 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s1182;
						end
					else if( ~x69 && x63 && ~x46 && ~x43 )
						nx_state = s670;
					else if( ~x69 && ~x63 && x64 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s691;
						end
					else if( ~x69 && ~x63 && ~x64 )
						begin
							y19 = 1'b1;	y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s1215;
						end
					else nx_state = s670;
				s671 : if( 1'b1 )
						begin
							y11 = 1'b1;	y24 = 1'b1;	
							nx_state = s1079;
						end
					else nx_state = s671;
				s672 : if( x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x20 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x20 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x20 )
						nx_state = s1;
					else nx_state = s672;
				s673 : if( x63 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x63 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x63 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x63 && ~x1 )
						nx_state = s1;
					else if( ~x63 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && x20 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && x20 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x63 && ~x20 )
						nx_state = s1;
					else nx_state = s673;
				s674 : if( x10 )
						begin
							y5 = 1'b1;	y42 = 1'b1;	y43 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s1216;
						end
					else if( ~x10 && x14 && x6 && x8 && x7 )
						begin
							y63 = 1'b1;	
							nx_state = s483;
						end
					else if( ~x10 && x14 && x6 && x8 && ~x7 && x9 && x18 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y45 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s672;
						end
					else if( ~x10 && x14 && x6 && x8 && ~x7 && x9 && ~x18 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x10 && x14 && x6 && x8 && ~x7 && x9 && ~x18 && x20 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x10 && x14 && x6 && x8 && ~x7 && x9 && ~x18 && x20 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x10 && x14 && x6 && x8 && ~x7 && x9 && ~x18 && ~x20 )
						nx_state = s1;
					else if( ~x10 && x14 && x6 && x8 && ~x7 && ~x9 && x19 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y45 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s672;
						end
					else if( ~x10 && x14 && x6 && x8 && ~x7 && ~x9 && ~x19 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x10 && x14 && x6 && x8 && ~x7 && ~x9 && ~x19 && x20 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x10 && x14 && x6 && x8 && ~x7 && ~x9 && ~x19 && x20 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x10 && x14 && x6 && x8 && ~x7 && ~x9 && ~x19 && ~x20 )
						nx_state = s1;
					else if( ~x10 && x14 && x6 && ~x8 && x9 && x7 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y5 = 1'b1;	
							y74 = 1'b1;	
							nx_state = s1217;
						end
					else if( ~x10 && x14 && x6 && ~x8 && x9 && ~x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y45 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s672;
						end
					else if( ~x10 && x14 && x6 && ~x8 && ~x9 && x7 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y45 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s672;
						end
					else if( ~x10 && x14 && x6 && ~x8 && ~x9 && x7 && ~x17 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x10 && x14 && x6 && ~x8 && ~x9 && x7 && ~x17 && x20 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x10 && x14 && x6 && ~x8 && ~x9 && x7 && ~x17 && x20 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x10 && x14 && x6 && ~x8 && ~x9 && x7 && ~x17 && ~x20 )
						nx_state = s1;
					else if( ~x10 && x14 && x6 && ~x8 && ~x9 && ~x7 )
						begin
							y65 = 1'b1;	
							nx_state = s393;
						end
					else if( ~x10 && x14 && ~x6 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x10 && ~x14 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y40 = 1'b1;	y45 = 1'b1;	
							nx_state = s1218;
						end
					else nx_state = s674;
				s675 : if( x64 && x63 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x64 && x63 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x64 && x63 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x64 && x63 && ~x11 )
						nx_state = s1;
					else if( x64 && ~x63 )
						begin
							y56 = 1'b1;	
							nx_state = s1219;
						end
					else if( ~x64 && x20 && x63 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x64 && x20 && ~x63 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x64 && x20 && ~x63 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x64 && x20 && ~x63 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x64 && ~x20 && x63 && x19 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x64 && ~x20 && x63 && ~x19 )
						begin
							y19 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x64 && ~x20 && ~x63 )
						nx_state = s1;
					else nx_state = s675;
				s676 : if( x63 && x20 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x63 && ~x20 && x19 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( x63 && ~x20 && ~x19 )
						begin
							y19 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x63 && x64 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x63 && x64 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x63 && x64 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( ~x63 && x64 && ~x14 )
						nx_state = s1;
					else if( ~x63 && ~x64 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x64 && x20 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x64 && x20 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x63 && ~x64 && ~x20 )
						nx_state = s1;
					else nx_state = s676;
				s677 : if( x64 && x6 && x8 && x27 && x7 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s1220;
						end
					else if( x64 && x6 && x8 && x27 && ~x7 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1220;
						end
					else if( x64 && x6 && x8 && ~x27 && x7 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x64 && x6 && x8 && ~x27 && ~x7 )
						begin
							y40 = 1'b1;	
							nx_state = s751;
						end
					else if( x64 && x6 && ~x8 && x27 && x7 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y47 = 1'b1;	
							nx_state = s1220;
						end
					else if( x64 && x6 && ~x8 && x27 && ~x7 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y46 = 1'b1;	
							nx_state = s1220;
						end
					else if( x64 && x6 && ~x8 && ~x27 && x7 )
						begin
							y39 = 1'b1;	
							nx_state = s277;
						end
					else if( x64 && x6 && ~x8 && ~x27 && ~x7 )
						begin
							y18 = 1'b1;	y41 = 1'b1;	y42 = 1'b1;	
							nx_state = s1221;
						end
					else if( x64 && ~x6 && x7 && x27 && x8 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y42 = 1'b1;	y44 = 1'b1;	
							nx_state = s1220;
						end
					else if( x64 && ~x6 && x7 && x27 && ~x8 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y42 = 1'b1;	y44 = 1'b1;	
							nx_state = s1220;
						end
					else if( x64 && ~x6 && x7 && ~x27 && x13 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x64 && ~x6 && x7 && ~x27 && x13 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x64 && ~x6 && x7 && ~x27 && x13 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x64 && ~x6 && x7 && ~x27 && x13 && x22 && ~x23 )
						nx_state = s1;
					else if( x64 && ~x6 && x7 && ~x27 && x13 && ~x22 )
						nx_state = s1;
					else if( x64 && ~x6 && x7 && ~x27 && ~x13 && x3 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x64 && ~x6 && x7 && ~x27 && ~x13 && x3 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x64 && ~x6 && x7 && ~x27 && ~x13 && x3 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x64 && ~x6 && x7 && ~x27 && ~x13 && x3 && x22 && ~x23 )
						nx_state = s1;
					else if( x64 && ~x6 && x7 && ~x27 && ~x13 && x3 && ~x22 )
						nx_state = s1;
					else if( x64 && ~x6 && x7 && ~x27 && ~x13 && ~x3 )
						begin
							y5 = 1'b1;	y34 = 1'b1;	y41 = 1'b1;	
							y42 = 1'b1;	
							nx_state = s1222;
						end
					else if( x64 && ~x6 && ~x7 && x27 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y42 = 1'b1;	y44 = 1'b1;	
							nx_state = s1220;
						end
					else if( x64 && ~x6 && ~x7 && ~x27 && x8 )
						begin
							y5 = 1'b1;	y17 = 1'b1;	y32 = 1'b1;	
							y42 = 1'b1;	
							nx_state = s1220;
						end
					else if( x64 && ~x6 && ~x7 && ~x27 && ~x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y32 = 1'b1;	
							nx_state = s1220;
						end
					else if( ~x64 )
						begin
							y57 = 1'b1;	
							nx_state = s1223;
						end
					else nx_state = s677;
				s678 : if( x65 && x4 )
						begin
							y67 = 1'b1;	
							nx_state = s1224;
						end
					else if( x65 && ~x4 && x6 && x5 && x7 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( x65 && ~x4 && x6 && x5 && x7 && ~x9 )
						begin
							y75 = 1'b1;	
							nx_state = s672;
						end
					else if( x65 && ~x4 && x6 && x5 && ~x7 && x8 && x9 && x12 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x65 && ~x4 && x6 && x5 && ~x7 && x8 && x9 && ~x12 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x65 && ~x4 && x6 && x5 && ~x7 && x8 && x9 && ~x12 && x20 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x4 && x6 && x5 && ~x7 && x8 && x9 && ~x12 && ~x20 )
						nx_state = s1;
					else if( x65 && ~x4 && x6 && x5 && ~x7 && x8 && ~x9 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x65 && ~x4 && x6 && x5 && ~x7 && x8 && ~x9 && ~x13 && x20 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x65 && ~x4 && x6 && x5 && ~x7 && x8 && ~x9 && ~x13 && x20 && ~x12 )
						nx_state = s1;
					else if( x65 && ~x4 && x6 && x5 && ~x7 && x8 && ~x9 && ~x13 && ~x20 )
						nx_state = s1;
					else if( x65 && ~x4 && x6 && x5 && ~x7 && ~x8 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y24 = 1'b1;	
							y25 = 1'b1;	y26 = 1'b1;	
							nx_state = s672;
						end
					else if( x65 && ~x4 && x6 && x5 && ~x7 && ~x8 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	y29 = 1'b1;	
							nx_state = s673;
						end
					else if( x65 && ~x4 && x6 && ~x5 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s674;
						end
					else if( x65 && ~x4 && x6 && ~x5 && ~x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y46 = 1'b1;	
							nx_state = s1218;
						end
					else if( x65 && ~x4 && ~x6 && x3 && x11 && x8 && x9 && x5 && x7 )
						begin
							y47 = 1'b1;	
							nx_state = s675;
						end
					else if( x65 && ~x4 && ~x6 && x3 && x11 && x8 && x9 && x5 && ~x7 )
						begin
							y51 = 1'b1;	
							nx_state = s655;
						end
					else if( x65 && ~x4 && ~x6 && x3 && x11 && x8 && x9 && ~x5 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	y16 = 1'b1;	
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s672;
						end
					else if( x65 && ~x4 && ~x6 && x3 && x11 && x8 && ~x9 && x5 && x7 )
						begin
							y48 = 1'b1;	
							nx_state = s676;
						end
					else if( x65 && ~x4 && ~x6 && x3 && x11 && x8 && ~x9 && x5 && ~x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s677;
						end
					else if( x65 && ~x4 && ~x6 && x3 && x11 && x8 && ~x9 && ~x5 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s672;
						end
					else if( x65 && ~x4 && ~x6 && x3 && x11 && ~x8 && x5 && x7 && x9 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( x65 && ~x4 && ~x6 && x3 && x11 && ~x8 && x5 && x7 && ~x9 )
						begin
							y50 = 1'b1;	
							nx_state = s658;
						end
					else if( x65 && ~x4 && ~x6 && x3 && x11 && ~x8 && x5 && ~x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y55 = 1'b1;	
							nx_state = s672;
						end
					else if( x65 && ~x4 && ~x6 && x3 && x11 && ~x8 && ~x5 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	y16 = 1'b1;	
							y18 = 1'b1;	y20 = 1'b1;	
							nx_state = s672;
						end
					else if( x65 && ~x4 && ~x6 && x3 && ~x11 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s674;
						end
					else if( x65 && ~x4 && ~x6 && ~x3 && x10 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y46 = 1'b1;	
							nx_state = s1218;
						end
					else if( x65 && ~x4 && ~x6 && ~x3 && ~x10 && x7 && x8 && x9 && x5 )
						begin
							y47 = 1'b1;	
							nx_state = s675;
						end
					else if( x65 && ~x4 && ~x6 && ~x3 && ~x10 && x7 && x8 && x9 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							nx_state = s672;
						end
					else if( x65 && ~x4 && ~x6 && ~x3 && ~x10 && x7 && x8 && ~x9 && x5 )
						begin
							y48 = 1'b1;	
							nx_state = s676;
						end
					else if( x65 && ~x4 && ~x6 && ~x3 && ~x10 && x7 && x8 && ~x9 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y34 = 1'b1;	
							y35 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							nx_state = s672;
						end
					else if( x65 && ~x4 && ~x6 && ~x3 && ~x10 && x7 && ~x8 && x9 && x5 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( x65 && ~x4 && ~x6 && ~x3 && ~x10 && x7 && ~x8 && x9 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	y38 = 1'b1;	
							nx_state = s672;
						end
					else if( x65 && ~x4 && ~x6 && ~x3 && ~x10 && x7 && ~x8 && ~x9 && x5 )
						begin
							y50 = 1'b1;	
							nx_state = s658;
						end
					else if( x65 && ~x4 && ~x6 && ~x3 && ~x10 && x7 && ~x8 && ~x9 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y34 = 1'b1;	
							y35 = 1'b1;	y39 = 1'b1;	
							nx_state = s672;
						end
					else if( x65 && ~x4 && ~x6 && ~x3 && ~x10 && ~x7 && x8 && x9 && x5 )
						begin
							y51 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x4 && ~x6 && ~x3 && ~x10 && ~x7 && x8 && x9 && ~x5 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	y40 = 1'b1;	
							nx_state = s672;
						end
					else if( x65 && ~x4 && ~x6 && ~x3 && ~x10 && ~x7 && x8 && ~x9 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y53 = 1'b1;	
							nx_state = s672;
						end
					else if( x65 && ~x4 && ~x6 && ~x3 && ~x10 && ~x7 && x8 && ~x9 && ~x5 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	y40 = 1'b1;	
							nx_state = s672;
						end
					else if( x65 && ~x4 && ~x6 && ~x3 && ~x10 && ~x7 && ~x8 && x5 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y54 = 1'b1;	
							nx_state = s672;
						end
					else if( x65 && ~x4 && ~x6 && ~x3 && ~x10 && ~x7 && ~x8 && x5 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s672;
						end
					else if( x65 && ~x4 && ~x6 && ~x3 && ~x10 && ~x7 && ~x8 && ~x5 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y40 = 1'b1;	
							nx_state = s672;
						end
					else if( ~x65 && x16 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x65 && ~x16 && x21 && x20 && x4 && x6 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( ~x65 && ~x16 && x21 && x20 && x4 && ~x6 )
						begin
							y38 = 1'b1;	
							nx_state = s845;
						end
					else if( ~x65 && ~x16 && x21 && x20 && ~x4 && x5 && x6 && x9 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x16 && x21 && x20 && ~x4 && x5 && x6 && ~x9 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && ~x16 && x21 && x20 && ~x4 && x5 && x6 && ~x9 && x17 && ~x8 )
						nx_state = s1;
					else if( ~x65 && ~x16 && x21 && x20 && ~x4 && x5 && x6 && ~x9 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x16 && x21 && x20 && ~x4 && x5 && ~x6 && x8 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x16 && x21 && x20 && ~x4 && x5 && ~x6 && ~x8 && x17 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && ~x16 && x21 && x20 && ~x4 && x5 && ~x6 && ~x8 && x17 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x16 && x21 && x20 && ~x4 && x5 && ~x6 && ~x8 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x16 && x21 && x20 && ~x4 && ~x5 && x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y39 = 1'b1;	y41 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x65 && ~x16 && x21 && x20 && ~x4 && ~x5 && ~x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y13 = 1'b1;	
							y40 = 1'b1;	y42 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x65 && ~x16 && x21 && ~x20 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1226;
						end
					else if( ~x65 && ~x16 && ~x21 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1226;
						end
					else if( ~x65 && ~x16 && ~x21 && ~x3 && x20 && x5 && x6 && x4 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x16 && ~x21 && ~x3 && x20 && x5 && x6 && ~x4 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y23 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x65 && ~x16 && ~x21 && ~x3 && x20 && x5 && ~x6 && x4 )
						begin
							y26 = 1'b1;	
							nx_state = s262;
						end
					else if( ~x65 && ~x16 && ~x21 && ~x3 && x20 && x5 && ~x6 && ~x4 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x65 && ~x16 && ~x21 && ~x3 && x20 && ~x5 && x6 && x4 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x16 && ~x21 && ~x3 && x20 && ~x5 && x6 && ~x4 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y13 = 1'b1;	
							y30 = 1'b1;	y45 = 1'b1;	
							nx_state = s1227;
						end
					else if( ~x65 && ~x16 && ~x21 && ~x3 && x20 && ~x5 && ~x6 && x4 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y13 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s1228;
						end
					else if( ~x65 && ~x16 && ~x21 && ~x3 && x20 && ~x5 && ~x6 && ~x4 )
						begin
							y3 = 1'b1;	y20 = 1'b1;	y30 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s1229;
						end
					else if( ~x65 && ~x16 && ~x21 && ~x3 && ~x20 && x4 && x5 )
						begin
							y5 = 1'b1;	y23 = 1'b1;	y24 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x65 && ~x16 && ~x21 && ~x3 && ~x20 && x4 && ~x5 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	y24 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x65 && ~x16 && ~x21 && ~x3 && ~x20 && ~x4 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	y23 = 1'b1;	
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s1225;
						end
					else nx_state = s678;
				s679 : if( x69 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x69 && x63 && x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x69 && x63 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s1230;
						end
					else if( ~x69 && ~x63 && x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x69 && ~x63 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else nx_state = s679;
				s680 : if( 1'b1 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else nx_state = s680;
				s681 : if( 1'b1 )
						begin
							y17 = 1'b1;	
							nx_state = s98;
						end
					else nx_state = s681;
				s682 : if( x21 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s301;
						end
					else if( ~x21 && x22 && x8 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && x8 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x12 && x23 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s666;
						end
					else if( ~x21 && ~x22 && x12 && ~x23 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && ~x22 && ~x12 && x23 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x22 && ~x12 && x23 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x22 && ~x12 && x23 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x12 && x23 && ~x9 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x12 && ~x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x22 && ~x12 && ~x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x22 && ~x12 && ~x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x12 && ~x23 && ~x8 )
						nx_state = s1;
					else nx_state = s682;
				s683 : if( x70 && x62 && x20 && x23 )
						begin
							y45 = 1'b1;	
							nx_state = s286;
						end
					else if( x70 && x62 && x20 && ~x23 )
						begin
							y1 = 1'b1;	y20 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	y44 = 1'b1;	
							nx_state = s535;
						end
					else if( x70 && x62 && ~x20 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s561;
						end
					else if( x70 && ~x62 && x64 )
						begin
							y7 = 1'b1;	y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s1231;
						end
					else if( x70 && ~x62 && ~x64 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x70 && x66 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else if( ~x70 && ~x66 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else nx_state = s683;
				s684 : if( 1'b1 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s315;
						end
					else nx_state = s684;
				s685 : if( x69 && x62 && x4 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x69 && x62 && x4 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y18 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1232;
						end
					else if( x69 && x62 && ~x4 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s633;
						end
					else if( x69 && ~x62 && x16 && x15 )
						nx_state = s1;
					else if( x69 && ~x62 && x16 && ~x15 && x4 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x69 && ~x62 && x16 && ~x15 && x4 && ~x5 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s638;
						end
					else if( x69 && ~x62 && x16 && ~x15 && ~x4 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s637;
						end
					else if( x69 && ~x62 && ~x16 && x15 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( x69 && ~x62 && ~x16 && ~x15 && x12 && x13 && x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s686;
						end
					else if( x69 && ~x62 && ~x16 && ~x15 && x12 && x13 && ~x3 && x14 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s686;
						end
					else if( x69 && ~x62 && ~x16 && ~x15 && x12 && x13 && ~x3 && ~x14 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( x69 && ~x62 && ~x16 && ~x15 && x12 && ~x13 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y22 = 1'b1;	
							nx_state = s61;
						end
					else if( x69 && ~x62 && ~x16 && ~x15 && ~x12 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x69 && x64 && x40 && x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s915;
						end
					else if( ~x69 && x64 && x40 && ~x10 && x25 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x69 && x64 && x40 && ~x10 && ~x25 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s910;
						end
					else if( ~x69 && x64 && ~x40 && x8 && x48 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( ~x69 && x64 && ~x40 && x8 && ~x48 && x37 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x69 && x64 && ~x40 && x8 && ~x48 && ~x37 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( ~x69 && x64 && ~x40 && ~x8 && x51 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( ~x69 && x64 && ~x40 && ~x8 && ~x51 && x37 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x69 && x64 && ~x40 && ~x8 && ~x51 && ~x37 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( ~x69 && ~x64 && x44 && x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s915;
						end
					else if( ~x69 && ~x64 && x44 && ~x10 && x25 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x69 && ~x64 && x44 && ~x10 && ~x25 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s910;
						end
					else if( ~x69 && ~x64 && ~x44 && x8 && x53 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( ~x69 && ~x64 && ~x44 && x8 && ~x53 && x36 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x69 && ~x64 && ~x44 && x8 && ~x53 && ~x36 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( ~x69 && ~x64 && ~x44 && ~x8 && x51 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( ~x69 && ~x64 && ~x44 && ~x8 && ~x51 && x36 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x69 && ~x64 && ~x44 && ~x8 && ~x51 && ~x36 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else nx_state = s685;
				s686 : if( x69 && x62 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s479;
						end
					else if( x69 && ~x62 && x15 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s60;
						end
					else if( x69 && ~x62 && ~x15 && x16 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( x69 && ~x62 && ~x15 && ~x16 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s627;
						end
					else if( ~x69 && x64 && x40 && x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x69 && x64 && x40 && ~x3 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1106;
						end
					else if( ~x69 && x64 && x40 && ~x3 && ~x2 && x28 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x69 && x64 && x40 && ~x3 && ~x2 && ~x28 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && x64 && ~x40 && x10 && x5 && x3 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x69 && x64 && ~x40 && x10 && x5 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x69 && x64 && ~x40 && x10 && x5 && ~x3 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x69 && x64 && ~x40 && x10 && ~x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x69 && x64 && ~x40 && ~x10 && x11 && x1 )
						begin
							y3 = 1'b1;	y13 = 1'b1;	y18 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s639;
						end
					else if( ~x69 && x64 && ~x40 && ~x10 && x11 && ~x1 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && x64 && ~x40 && ~x10 && x11 && ~x1 && ~x3 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x69 && x64 && ~x40 && ~x10 && ~x11 )
						nx_state = s686;
					else if( ~x69 && ~x64 && x44 && x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x69 && ~x64 && x44 && ~x3 && x34 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s1107;
						end
					else if( ~x69 && ~x64 && x44 && ~x3 && ~x34 && x28 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x69 && ~x64 && x44 && ~x3 && ~x34 && ~x28 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s509;
						end
					else if( ~x69 && ~x64 && ~x44 && x10 && x5 && x41 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( ~x69 && ~x64 && ~x44 && x10 && x5 && ~x41 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x69 && ~x64 && ~x44 && x10 && x5 && ~x41 && ~x4 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s631;
						end
					else if( ~x69 && ~x64 && ~x44 && x10 && ~x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x69 && ~x64 && ~x44 && ~x10 && x37 && x11 )
						begin
							y3 = 1'b1;	y13 = 1'b1;	y22 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s640;
						end
					else if( ~x69 && ~x64 && ~x44 && ~x10 && x37 && ~x11 )
						nx_state = s686;
					else if( ~x69 && ~x64 && ~x44 && ~x10 && ~x37 && x41 && x11 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else if( ~x69 && ~x64 && ~x44 && ~x10 && ~x37 && x41 && ~x11 )
						nx_state = s686;
					else if( ~x69 && ~x64 && ~x44 && ~x10 && ~x37 && ~x41 && x11 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x69 && ~x64 && ~x44 && ~x10 && ~x37 && ~x41 && ~x11 )
						nx_state = s686;
					else nx_state = s686;
				s687 : if( 1'b1 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y29 = 1'b1;	
							nx_state = s690;
						end
					else nx_state = s687;
				s688 : if( x12 && x63 && x46 && x13 && x3 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s689;
						end
					else if( x12 && x63 && x46 && x13 && ~x3 && x14 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s689;
						end
					else if( x12 && x63 && x46 && x13 && ~x3 && ~x14 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s691;
						end
					else if( x12 && x63 && x46 && ~x13 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s692;
						end
					else if( x12 && x63 && ~x46 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s693;
						end
					else if( x12 && ~x63 && x15 && x13 && x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s699;
						end
					else if( x12 && ~x63 && x15 && x13 && ~x3 && x14 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s699;
						end
					else if( x12 && ~x63 && x15 && x13 && ~x3 && ~x14 && x64 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( x12 && ~x63 && x15 && x13 && ~x3 && ~x14 && ~x64 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s700;
						end
					else if( x12 && ~x63 && x15 && ~x13 && x64 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s692;
						end
					else if( x12 && ~x63 && x15 && ~x13 && ~x64 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s701;
						end
					else if( x12 && ~x63 && ~x15 && x64 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s693;
						end
					else if( x12 && ~x63 && ~x15 && ~x64 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s702;
						end
					else if( ~x12 && x63 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s693;
						end
					else if( ~x12 && ~x63 && x64 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s693;
						end
					else if( ~x12 && ~x63 && ~x64 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s702;
						end
					else nx_state = s688;
				s689 : if( 1'b1 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else nx_state = s689;
				s690 : if( 1'b1 )
						begin
							y3 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s883;
						end
					else nx_state = s690;
				s691 : if( x69 )
						nx_state = s1;
					else if( ~x69 && x63 && x15 && x13 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y27 = 1'b1;	
							nx_state = s696;
						end
					else if( ~x69 && x63 && x15 && ~x13 )
						begin
							y8 = 1'b1;	
							nx_state = s783;
						end
					else if( ~x69 && x63 && ~x15 && x12 )
						begin
							y8 = 1'b1;	
							nx_state = s783;
						end
					else if( ~x69 && x63 && ~x15 && ~x12 )
						nx_state = s691;
					else if( ~x69 && ~x63 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s216;
						end
					else nx_state = s691;
				s692 : if( x15 && x63 && x45 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s670;
						end
					else if( x15 && x63 && ~x45 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s691;
						end
					else if( x15 && ~x63 && x14 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s1233;
						end
					else if( x15 && ~x63 && ~x14 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( ~x15 && x63 && x43 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s1182;
						end
					else if( ~x15 && x63 && ~x43 )
						nx_state = s692;
					else if( ~x15 && ~x63 && x12 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s1234;
						end
					else if( ~x15 && ~x63 && ~x12 )
						nx_state = s692;
					else nx_state = s692;
				s693 : if( x69 )
						begin
							y3 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1235;
						end
					else if( ~x69 && x15 && x63 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s1182;
						end
					else if( ~x69 && x15 && ~x63 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s1234;
						end
					else if( ~x69 && ~x15 && x6 && x63 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s670;
						end
					else if( ~x69 && ~x15 && x6 && ~x63 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s1233;
						end
					else if( ~x69 && ~x15 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s692;
						end
					else nx_state = s693;
				s694 : if( x15 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s997;
						end
					else if( ~x15 && x63 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y33 = 1'b1;	
							nx_state = s1236;
						end
					else if( ~x15 && ~x63 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s216;
						end
					else nx_state = s694;
				s695 : if( x15 && x63 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y33 = 1'b1;	
							nx_state = s1236;
						end
					else if( x15 && ~x63 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s216;
						end
					else if( ~x15 && x63 && x37 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x15 && x63 && ~x37 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s697;
						end
					else if( ~x15 && ~x63 && x6 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x15 && ~x63 && ~x6 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s705;
						end
					else nx_state = s695;
				s696 : if( x15 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y33 = 1'b1;	
							nx_state = s1236;
						end
					else if( ~x15 && x42 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( ~x15 && ~x42 && x41 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s688;
						end
					else if( ~x15 && ~x42 && ~x41 )
						nx_state = s696;
					else nx_state = s696;
				s697 : if( x15 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x15 && x39 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y27 = 1'b1;	
							nx_state = s696;
						end
					else if( ~x15 && ~x39 && x40 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y27 = 1'b1;	
							nx_state = s696;
						end
					else if( ~x15 && ~x39 && ~x40 && x10 && x37 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x15 && ~x39 && ~x40 && x10 && ~x37 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s697;
						end
					else if( ~x15 && ~x39 && ~x40 && ~x10 && x42 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( ~x15 && ~x39 && ~x40 && ~x10 && ~x42 )
						nx_state = s697;
					else nx_state = s697;
				s698 : if( x62 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s762;
						end
					else if( ~x62 && x64 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s670;
						end
					else if( ~x62 && ~x64 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s456;
						end
					else nx_state = s698;
				s699 : if( 1'b1 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s627;
						end
					else nx_state = s699;
				s700 : if( x15 && x13 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s704;
						end
					else if( x15 && ~x13 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s1237;
						end
					else if( ~x15 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s1237;
						end
					else if( ~x15 && ~x12 )
						nx_state = s700;
					else nx_state = s700;
				s701 : if( x15 && x14 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s1233;
						end
					else if( x15 && ~x14 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s700;
						end
					else if( ~x15 && x12 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s1234;
						end
					else if( ~x15 && ~x12 )
						nx_state = s701;
					else nx_state = s701;
				s702 : if( x15 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s1234;
						end
					else if( ~x15 && x6 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s1233;
						end
					else if( ~x15 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s701;
						end
					else nx_state = s702;
				s703 : if( x15 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s999;
						end
					else if( ~x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s216;
						end
					else nx_state = s703;
				s704 : if( x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s216;
						end
					else if( ~x15 && x11 && x64 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( ~x15 && x11 && ~x64 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s703;
						end
					else if( ~x15 && ~x11 && x10 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s688;
						end
					else if( ~x15 && ~x11 && ~x10 )
						nx_state = s704;
					else nx_state = s704;
				s705 : if( x15 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x15 && x8 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s704;
						end
					else if( ~x15 && ~x8 && x9 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s704;
						end
					else if( ~x15 && ~x8 && ~x9 && x10 && x6 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x15 && ~x8 && ~x9 && x10 && ~x6 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s705;
						end
					else if( ~x15 && ~x8 && ~x9 && ~x10 && x64 && x11 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( ~x15 && ~x8 && ~x9 && ~x10 && x64 && ~x11 )
						nx_state = s705;
					else if( ~x15 && ~x8 && ~x9 && ~x10 && ~x64 && x11 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s703;
						end
					else if( ~x15 && ~x8 && ~x9 && ~x10 && ~x64 && ~x11 )
						nx_state = s705;
					else nx_state = s705;
				s706 : if( 1'b1 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else nx_state = s706;
				s707 : if( x60 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x60 && ~x7 && x61 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x60 && ~x7 && x61 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x60 && ~x7 && x61 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x60 && ~x7 && x61 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s329;
						end
					else if( x60 && ~x7 && ~x61 )
						nx_state = s118;
					else if( ~x60 && x61 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x60 && x61 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x60 && x61 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( ~x60 && x61 && x62 && ~x18 )
						nx_state = s1;
					else if( ~x60 && x61 && ~x62 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x60 && x61 && ~x62 && ~x7 )
						nx_state = s118;
					else if( ~x60 && ~x61 && x62 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x60 && ~x61 && ~x62 )
						nx_state = s47;
					else nx_state = s707;
				s708 : if( x63 && x18 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							y17 = 1'b1;	y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1238;
						end
					else if( x63 && ~x18 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1239;
						end
					else if( ~x63 )
						begin
							y4 = 1'b1;	y31 = 1'b1;	y39 = 1'b1;	
							nx_state = s1240;
						end
					else nx_state = s708;
				s709 : if( x62 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y48 = 1'b1;	y50 = 1'b1;	
							nx_state = s1241;
						end
					else if( ~x62 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y31 = 1'b1;	
							nx_state = s1242;
						end
					else nx_state = s709;
				s710 : if( x64 )
						begin
							y15 = 1'b1;	y36 = 1'b1;	
							nx_state = s1243;
						end
					else if( ~x64 )
						begin
							y33 = 1'b1;	
							nx_state = s589;
						end
					else nx_state = s710;
				s711 : if( x64 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x64 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x64 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x64 && ~x14 )
						nx_state = s1;
					else if( ~x64 && x30 )
						begin
							y47 = 1'b1;	y50 = 1'b1;	y61 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s1148;
						end
					else if( ~x64 && ~x30 && x31 )
						begin
							y47 = 1'b1;	y50 = 1'b1;	y61 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s1244;
						end
					else if( ~x64 && ~x30 && ~x31 )
						begin
							y33 = 1'b1;	
							nx_state = s589;
						end
					else nx_state = s711;
				s712 : if( x65 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y69 = 1'b1;	
							y70 = 1'b1;	y71 = 1'b1;	
							nx_state = s1245;
						end
					else if( ~x65 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1179;
						end
					else nx_state = s712;
				s713 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s1246;
						end
					else nx_state = s713;
				s714 : if( x64 && x63 )
						nx_state = s1;
					else if( x64 && ~x63 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x64 && ~x63 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x64 && ~x63 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x64 && ~x63 && ~x18 )
						nx_state = s1;
					else if( ~x64 && x63 && x66 && x10 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x64 && x63 && x66 && ~x10 )
						begin
							y19 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x64 && x63 && ~x66 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( ~x64 && x63 && ~x66 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( ~x64 && x63 && ~x66 && x19 && ~x14 && ~x13 && x11 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( ~x64 && x63 && ~x66 && x19 && ~x14 && ~x13 && x11 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x64 && x63 && ~x66 && x19 && ~x14 && ~x13 && ~x11 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x64 && x63 && ~x66 && ~x19 )
						nx_state = s1;
					else if( ~x64 && ~x63 && x65 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x64 && ~x63 && x65 && x20 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x64 && ~x63 && x65 && x20 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x64 && ~x63 && x65 && ~x20 )
						nx_state = s1;
					else if( ~x64 && ~x63 && ~x65 && x21 && x22 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x64 && ~x63 && ~x65 && x21 && ~x22 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x64 && ~x63 && ~x65 && x21 && ~x22 && ~x23 )
						nx_state = s1;
					else if( ~x64 && ~x63 && ~x65 && ~x21 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x64 && ~x63 && ~x65 && ~x21 && ~x23 )
						nx_state = s1;
					else nx_state = s714;
				s715 : if( x2 )
						nx_state = s1;
					else if( ~x2 && x3 && x4 && x5 && x1 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x2 && x3 && x4 && x5 && ~x1 )
						begin
							y41 = 1'b1;	y45 = 1'b1;	y46 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x2 && x3 && x4 && ~x5 && x1 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x2 && x3 && x4 && ~x5 && ~x1 )
						begin
							y39 = 1'b1;	y43 = 1'b1;	y44 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x2 && x3 && ~x4 && x5 && x1 )
						begin
							y51 = 1'b1;	
							nx_state = s655;
						end
					else if( ~x2 && x3 && ~x4 && x5 && ~x1 )
						begin
							y41 = 1'b1;	y42 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x2 && x3 && ~x4 && ~x5 && x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y48 = 1'b1;	
							y50 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x2 && x3 && ~x4 && ~x5 && ~x1 )
						begin
							y39 = 1'b1;	y40 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x2 && ~x3 && x4 && x5 && x1 && x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s651;
						end
					else if( ~x2 && ~x3 && x4 && x5 && x1 && ~x6 && x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s651;
						end
					else if( ~x2 && ~x3 && x4 && x5 && x1 && ~x6 && ~x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s652;
						end
					else if( ~x2 && ~x3 && x4 && x5 && ~x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y47 = 1'b1;	y48 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x2 && ~x3 && x4 && ~x5 && x1 && x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s653;
						end
					else if( ~x2 && ~x3 && x4 && ~x5 && x1 && ~x6 && x7 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s653;
						end
					else if( ~x2 && ~x3 && x4 && ~x5 && x1 && ~x6 && ~x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x2 && ~x3 && x4 && ~x5 && ~x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y48 = 1'b1;	y49 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x2 && ~x3 && ~x4 && x1 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x2 && ~x3 && ~x4 && x1 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x2 && ~x3 && ~x4 && ~x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y32 = 1'b1;	y48 = 1'b1;	
							nx_state = s654;
						end
					else nx_state = s715;
				s716 : if( x6 )
						begin
							y30 = 1'b1;	
							nx_state = s976;
						end
					else if( ~x6 && x2 && x1 && x4 && x3 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x6 && x2 && x1 && x4 && x3 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x6 && x2 && x1 && x4 && x3 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( ~x6 && x2 && x1 && x4 && x3 && ~x22 )
						nx_state = s1;
					else if( ~x6 && x2 && x1 && x4 && ~x3 && x5 && x18 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x6 && x2 && x1 && x4 && ~x3 && x5 && ~x18 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x6 && x2 && x1 && x4 && ~x3 && x5 && ~x18 && x22 && ~x21 )
						nx_state = s1;
					else if( ~x6 && x2 && x1 && x4 && ~x3 && x5 && ~x18 && ~x22 )
						nx_state = s1;
					else if( ~x6 && x2 && x1 && x4 && ~x3 && ~x5 && x21 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x6 && x2 && x1 && x4 && ~x3 && ~x5 && ~x21 && x22 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x6 && x2 && x1 && x4 && ~x3 && ~x5 && ~x21 && x22 && ~x18 )
						nx_state = s1;
					else if( ~x6 && x2 && x1 && x4 && ~x3 && ~x5 && ~x21 && ~x22 )
						nx_state = s1;
					else if( ~x6 && x2 && x1 && ~x4 && x5 && x3 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x6 && x2 && x1 && ~x4 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	y36 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x6 && x2 && x1 && ~x4 && ~x5 && x3 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x6 && x2 && x1 && ~x4 && ~x5 && ~x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y34 = 1'b1;	y37 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x6 && x2 && ~x1 && x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s1247;
						end
					else if( ~x6 && x2 && ~x1 && ~x3 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s1247;
						end
					else if( ~x6 && x2 && ~x1 && ~x3 && ~x4 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s1247;
						end
					else if( ~x6 && x2 && ~x1 && ~x3 && ~x4 && ~x5 )
						begin
							y38 = 1'b1;	
							nx_state = s845;
						end
					else if( ~x6 && ~x2 && x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s1248;
						end
					else if( ~x6 && ~x2 && ~x7 && x3 && x4 && x5 && x1 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x6 && ~x2 && ~x7 && x3 && x4 && x5 && ~x1 )
						begin
							y41 = 1'b1;	y45 = 1'b1;	y46 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x6 && ~x2 && ~x7 && x3 && x4 && ~x5 && x1 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x6 && ~x2 && ~x7 && x3 && x4 && ~x5 && ~x1 )
						begin
							y39 = 1'b1;	y43 = 1'b1;	y44 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x6 && ~x2 && ~x7 && x3 && ~x4 && x5 && x1 )
						begin
							y51 = 1'b1;	
							nx_state = s655;
						end
					else if( ~x6 && ~x2 && ~x7 && x3 && ~x4 && x5 && ~x1 )
						begin
							y41 = 1'b1;	y42 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x6 && ~x2 && ~x7 && x3 && ~x4 && ~x5 && x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y48 = 1'b1;	
							y50 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x6 && ~x2 && ~x7 && x3 && ~x4 && ~x5 && ~x1 )
						begin
							y39 = 1'b1;	y40 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x6 && ~x2 && ~x7 && ~x3 && x1 && x5 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s328;
						end
					else if( ~x6 && ~x2 && ~x7 && ~x3 && x1 && ~x5 && x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y4 = 1'b1;	
							nx_state = s71;
						end
					else if( ~x6 && ~x2 && ~x7 && ~x3 && x1 && ~x5 && ~x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x6 && ~x2 && ~x7 && ~x3 && ~x1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s1249;
						end
					else nx_state = s716;
				s717 : if( x65 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s1250;
						end
					else if( ~x65 && x21 && x20 )
						begin
							y15 = 1'b1;	
							nx_state = s22;
						end
					else if( ~x65 && x21 && ~x20 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1251;
						end
					else if( ~x65 && ~x21 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1251;
						end
					else nx_state = s717;
				s718 : if( x63 && x65 && x17 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( x63 && x65 && ~x17 && x14 )
						begin
							y38 = 1'b1;	y39 = 1'b1;	
							nx_state = s1252;
						end
					else if( x63 && x65 && ~x17 && ~x14 )
						begin
							y36 = 1'b1;	y37 = 1'b1;	
							nx_state = s1253;
						end
					else if( x63 && ~x65 )
						begin
							y3 = 1'b1;	y18 = 1'b1;	y53 = 1'b1;	
							nx_state = s1254;
						end
					else if( ~x63 && x4 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x63 && x4 && ~x11 && x30 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s789;
						end
					else if( ~x63 && x4 && ~x11 && x30 && ~x12 && x9 && x10 && x8 )
						begin
							y11 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x63 && x4 && ~x11 && x30 && ~x12 && x9 && x10 && ~x8 )
						begin
							y8 = 1'b1;	
							nx_state = s1255;
						end
					else if( ~x63 && x4 && ~x11 && x30 && ~x12 && x9 && ~x10 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else if( ~x63 && x4 && ~x11 && x30 && ~x12 && x9 && ~x10 && ~x8 )
						begin
							y8 = 1'b1;	
							nx_state = s1256;
						end
					else if( ~x63 && x4 && ~x11 && x30 && ~x12 && ~x9 && x10 && x8 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else if( ~x63 && x4 && ~x11 && x30 && ~x12 && ~x9 && x10 && ~x8 && x27 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x63 && x4 && ~x11 && x30 && ~x12 && ~x9 && x10 && ~x8 && ~x27 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x63 && x4 && ~x11 && x30 && ~x12 && ~x9 && ~x10 && x8 )
						begin
							y8 = 1'b1;	
							nx_state = s1257;
						end
					else if( ~x63 && x4 && ~x11 && x30 && ~x12 && ~x9 && ~x10 && ~x8 && x26 )
						begin
							y17 = 1'b1;	
							nx_state = s98;
						end
					else if( ~x63 && x4 && ~x11 && x30 && ~x12 && ~x9 && ~x10 && ~x8 && ~x26 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x63 && x4 && ~x11 && ~x30 && x31 && x15 )
						begin
							y14 = 1'b1;	
							nx_state = s228;
						end
					else if( ~x63 && x4 && ~x11 && ~x30 && x31 && ~x15 )
						begin
							y3 = 1'b1;	
							nx_state = s462;
						end
					else if( ~x63 && x4 && ~x11 && ~x30 && ~x31 && x8 && x9 )
						begin
							y47 = 1'b1;	y55 = 1'b1;	y63 = 1'b1;	
							y70 = 1'b1;	
							nx_state = s1175;
						end
					else if( ~x63 && x4 && ~x11 && ~x30 && ~x31 && x8 && ~x9 )
						begin
							y47 = 1'b1;	y56 = 1'b1;	y63 = 1'b1;	
							y71 = 1'b1;	
							nx_state = s1175;
						end
					else if( ~x63 && x4 && ~x11 && ~x30 && ~x31 && ~x8 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s835;
						end
					else if( ~x63 && x4 && ~x11 && ~x30 && ~x31 && ~x8 && ~x12 )
						begin
							y45 = 1'b1;	y46 = 1'b1;	y47 = 1'b1;	
							y55 = 1'b1;	y60 = 1'b1;	y63 = 1'b1;	
							y70 = 1'b1;	
							nx_state = s1175;
						end
					else if( ~x63 && ~x4 && x30 )
						begin
							y5 = 1'b1;	
							nx_state = s562;
						end
					else if( ~x63 && ~x4 && ~x30 && x31 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( ~x63 && ~x4 && ~x30 && ~x31 )
						begin
							y5 = 1'b1;	
							nx_state = s560;
						end
					else nx_state = s718;
				s719 : if( 1'b1 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s1258;
						end
					else nx_state = s719;
				s720 : if( x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x19 && ~x14 && ~x13 && x11 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( x19 && ~x14 && ~x13 && x11 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( x19 && ~x14 && ~x13 && ~x11 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x19 )
						nx_state = s1;
					else nx_state = s720;
				s721 : if( x21 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s224;
						end
					else nx_state = s721;
				s722 : if( x20 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1259;
						end
					else if( ~x20 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x20 && ~x10 )
						nx_state = s1;
					else nx_state = s722;
				s723 : if( x21 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x21 && x22 && x8 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && x8 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x12 && x23 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s666;
						end
					else if( ~x21 && ~x22 && x12 && ~x23 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && ~x22 && ~x12 && x23 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x22 && ~x12 && x23 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x22 && ~x12 && x23 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x12 && x23 && ~x9 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x12 && ~x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x22 && ~x12 && ~x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x22 && ~x12 && ~x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x12 && ~x23 && ~x8 )
						nx_state = s1;
					else nx_state = s723;
				s724 : if( x21 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x21 && x22 && x23 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && x22 && x23 && ~x12 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && x23 && ~x12 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && x23 && ~x12 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x12 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x8 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x8 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && ~x18 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s476;
						end
					else nx_state = s724;
				s725 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1260;
						end
					else nx_state = s725;
				s726 : if( x11 )
						begin
							y20 = 1'b1;	
							nx_state = s1261;
						end
					else if( ~x11 )
						begin
							y67 = 1'b1;	
							nx_state = s1224;
						end
					else nx_state = s726;
				s727 : if( x17 )
						begin
							y24 = 1'b1;	
							nx_state = s1262;
						end
					else if( ~x17 )
						begin
							y5 = 1'b1;	y13 = 1'b1;	y30 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s727;
						end
					else nx_state = s727;
				s728 : if( x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x22 && ~x17 )
						nx_state = s1;
					else if( ~x22 && x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x22 && ~x23 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else nx_state = s728;
				s729 : if( x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x22 && ~x17 )
						nx_state = s1;
					else if( ~x22 && x23 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x22 && x23 && x15 && ~x8 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x22 && x23 && ~x15 && x16 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s486;
						end
					else if( ~x22 && x23 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( ~x22 && ~x23 && x18 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x22 && ~x23 && x18 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x22 && ~x23 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x22 && ~x23 && ~x18 )
						nx_state = s1;
					else nx_state = s729;
				s730 : if( x65 && x22 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s625;
						end
					else if( x65 && ~x22 && x23 && x15 && x16 && x14 && x8 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x65 && ~x22 && x23 && x15 && x16 && x14 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x65 && ~x22 && x23 && x15 && x16 && ~x14 && x7 && x8 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x65 && ~x22 && x23 && x15 && x16 && ~x14 && x7 && ~x8 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s358;
						end
					else if( x65 && ~x22 && x23 && x15 && x16 && ~x14 && ~x7 && x8 && x12 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x65 && ~x22 && x23 && x15 && x16 && ~x14 && ~x7 && x8 && ~x12 && x18 && x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x65 && ~x22 && x23 && x15 && x16 && ~x14 && ~x7 && x8 && ~x12 && x18 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 && x15 && x16 && ~x14 && ~x7 && x8 && ~x12 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 && x15 && x16 && ~x14 && ~x7 && ~x8 && x13 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( x65 && ~x22 && x23 && x15 && x16 && ~x14 && ~x7 && ~x8 && ~x13 && x18 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x65 && ~x22 && x23 && x15 && x16 && ~x14 && ~x7 && ~x8 && ~x13 && x18 && ~x12 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 && x15 && x16 && ~x14 && ~x7 && ~x8 && ~x13 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 && x15 && ~x16 && x7 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x65 && ~x22 && x23 && x15 && ~x16 && ~x7 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( x65 && ~x22 && x23 && x15 && ~x16 && ~x7 && ~x2 && x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y28 = 1'b1;	
							nx_state = s729;
						end
					else if( x65 && ~x22 && x23 && x15 && ~x16 && ~x7 && ~x2 && ~x3 && x8 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s625;
						end
					else if( x65 && ~x22 && x23 && x15 && ~x16 && ~x7 && ~x2 && ~x3 && ~x8 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	
							nx_state = s486;
						end
					else if( x65 && ~x22 && x23 && ~x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && x7 && x11 && x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y28 = 1'b1;	
							nx_state = s729;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && x7 && x11 && ~x3 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && x7 && ~x11 && x8 && x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y28 = 1'b1;	
							nx_state = s729;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && x7 && ~x11 && x8 && ~x3 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && x7 && ~x11 && ~x8 && x18 && x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && x7 && ~x11 && ~x8 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && x7 && ~x11 && ~x8 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && x7 && ~x11 && ~x8 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && x8 && x9 && x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y28 = 1'b1;	
							nx_state = s729;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && x8 && x9 && ~x3 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && x8 && ~x9 && x18 && x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && x8 && ~x9 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && x8 && ~x9 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && x8 && ~x9 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && x10 && x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y28 = 1'b1;	
							nx_state = s729;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && x10 && ~x3 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && ~x10 && x18 && x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && ~x10 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && ~x10 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && ~x10 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && ~x16 && x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y28 = 1'b1;	
							nx_state = s729;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && ~x16 && ~x3 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s728;
						end
					else if( x65 && ~x22 && ~x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x65 && x67 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x65 && x67 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x65 && x67 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( ~x65 && x67 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y28 = 1'b1;	
							nx_state = s299;
						end
					else if( ~x65 && ~x67 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s12;
						end
					else nx_state = s730;
				s731 : if( x70 && x6 )
						begin
							y2 = 1'b1;	
							nx_state = s1111;
						end
					else if( x70 && ~x6 && x14 && x21 && x9 )
						begin
							y44 = 1'b1;	
							nx_state = s755;
						end
					else if( x70 && ~x6 && x14 && x21 && ~x9 )
						begin
							y44 = 1'b1;	
							nx_state = s1138;
						end
					else if( x70 && ~x6 && x14 && ~x21 && x5 && x8 && x7 )
						begin
							y44 = 1'b1;	
							nx_state = s755;
						end
					else if( x70 && ~x6 && x14 && ~x21 && x5 && x8 && ~x7 && x9 && x18 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1263;
						end
					else if( x70 && ~x6 && x14 && ~x21 && x5 && x8 && ~x7 && x9 && ~x18 && x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x70 && ~x6 && x14 && ~x21 && x5 && x8 && ~x7 && x9 && ~x18 && x10 && ~x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x70 && ~x6 && x14 && ~x21 && x5 && x8 && ~x7 && x9 && ~x18 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x6 && x14 && ~x21 && x5 && x8 && ~x7 && x9 && ~x18 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x6 && x14 && ~x21 && x5 && x8 && ~x7 && ~x9 && x19 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1263;
						end
					else if( x70 && ~x6 && x14 && ~x21 && x5 && x8 && ~x7 && ~x9 && ~x19 && x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x70 && ~x6 && x14 && ~x21 && x5 && x8 && ~x7 && ~x9 && ~x19 && x10 && ~x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x70 && ~x6 && x14 && ~x21 && x5 && x8 && ~x7 && ~x9 && ~x19 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x6 && x14 && ~x21 && x5 && x8 && ~x7 && ~x9 && ~x19 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x6 && x14 && ~x21 && x5 && ~x8 && x7 && x9 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else if( x70 && ~x6 && x14 && ~x21 && x5 && ~x8 && x7 && ~x9 && x20 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1263;
						end
					else if( x70 && ~x6 && x14 && ~x21 && x5 && ~x8 && x7 && ~x9 && ~x20 && x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x70 && ~x6 && x14 && ~x21 && x5 && ~x8 && x7 && ~x9 && ~x20 && x10 && ~x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x70 && ~x6 && x14 && ~x21 && x5 && ~x8 && x7 && ~x9 && ~x20 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x70 && ~x6 && x14 && ~x21 && x5 && ~x8 && x7 && ~x9 && ~x20 && ~x10 )
						nx_state = s1;
					else if( x70 && ~x6 && x14 && ~x21 && x5 && ~x8 && ~x7 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1263;
						end
					else if( x70 && ~x6 && x14 && ~x21 && ~x5 )
						begin
							y44 = 1'b1;	
							nx_state = s755;
						end
					else if( x70 && ~x6 && ~x14 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y21 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s1264;
						end
					else if( ~x70 && x21 && x15 && x20 && x10 && x11 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s600;
						end
					else if( ~x70 && x21 && x15 && x20 && x10 && ~x11 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s601;
						end
					else if( ~x70 && x21 && x15 && x20 && ~x10 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( ~x70 && x21 && x15 && x20 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s602;
						end
					else if( ~x70 && x21 && x15 && ~x20 && x5 && x10 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s605;
						end
					else if( ~x70 && x21 && x15 && ~x20 && x5 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s600;
						end
					else if( ~x70 && x21 && x15 && ~x20 && x5 && x10 && ~x11 && ~x12 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x70 && x21 && x15 && ~x20 && x5 && ~x10 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s777;
						end
					else if( ~x70 && x21 && x15 && ~x20 && x5 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	
							nx_state = s133;
						end
					else if( ~x70 && x21 && x15 && ~x20 && ~x5 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x70 && x21 && ~x15 && x16 && x10 && x12 && x20 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y11 = 1'b1;	
							nx_state = s600;
						end
					else if( ~x70 && x21 && ~x15 && x16 && x10 && x12 && ~x20 && x8 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x70 && x21 && ~x15 && x16 && x10 && x12 && ~x20 && ~x8 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x21 && ~x15 && x16 && x10 && x12 && ~x20 && ~x8 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x21 && ~x15 && x16 && x10 && x12 && ~x20 && ~x8 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x15 && x16 && x10 && x12 && ~x20 && ~x8 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x15 && x16 && x10 && ~x12 && x20 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x70 && x21 && ~x15 && x16 && x10 && ~x12 && ~x20 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x70 && x21 && ~x15 && x16 && ~x10 && x20 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y11 = 1'b1;	
							nx_state = s600;
						end
					else if( ~x70 && x21 && ~x15 && x16 && ~x10 && ~x20 && x12 && x7 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x70 && x21 && ~x15 && x16 && ~x10 && ~x20 && x12 && ~x7 && x11 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x70 && x21 && ~x15 && x16 && ~x10 && ~x20 && x12 && ~x7 && ~x11 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x21 && ~x15 && x16 && ~x10 && ~x20 && x12 && ~x7 && ~x11 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x21 && ~x15 && x16 && ~x10 && ~x20 && x12 && ~x7 && ~x11 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x15 && x16 && ~x10 && ~x20 && x12 && ~x7 && ~x11 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x15 && x16 && ~x10 && ~x20 && ~x12 && x11 && x9 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x70 && x21 && ~x15 && x16 && ~x10 && ~x20 && ~x12 && x11 && ~x9 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x21 && ~x15 && x16 && ~x10 && ~x20 && ~x12 && x11 && ~x9 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x21 && ~x15 && x16 && ~x10 && ~x20 && ~x12 && x11 && ~x9 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x15 && x16 && ~x10 && ~x20 && ~x12 && x11 && ~x9 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x15 && x16 && ~x10 && ~x20 && ~x12 && ~x11 && x8 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x21 && ~x15 && x16 && ~x10 && ~x20 && ~x12 && ~x11 && x8 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x70 && x21 && ~x15 && x16 && ~x10 && ~x20 && ~x12 && ~x11 && x8 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x15 && x16 && ~x10 && ~x20 && ~x12 && ~x11 && x8 && ~x19 )
						nx_state = s1;
					else if( ~x70 && x21 && ~x15 && x16 && ~x10 && ~x20 && ~x12 && ~x11 && ~x8 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x70 && x21 && ~x15 && ~x16 && x20 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x70 && x21 && ~x15 && ~x16 && ~x20 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x70 && x21 && ~x15 && ~x16 && ~x20 && ~x5 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x70 && ~x21 && x3 && x15 && x10 && x11 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s600;
						end
					else if( ~x70 && ~x21 && x3 && x15 && x10 && ~x11 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s601;
						end
					else if( ~x70 && ~x21 && x3 && x15 && x10 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y13 = 1'b1;	
							nx_state = s600;
						end
					else if( ~x70 && ~x21 && x3 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( ~x70 && ~x21 && x3 && x15 && ~x10 && ~x12 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s556;
						end
					else if( ~x70 && ~x21 && x3 && ~x15 && x16 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s625;
						end
					else if( ~x70 && ~x21 && x3 && ~x15 && ~x16 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s209;
						end
					else if( ~x70 && ~x21 && ~x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s625;
						end
					else nx_state = s731;
				s732 : if( x70 && x63 && x64 && x55 && x33 && x32 && x8 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s739;
						end
					else if( x70 && x63 && x64 && x55 && x33 && x32 && ~x8 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s909;
						end
					else if( x70 && x63 && x64 && x55 && x33 && ~x32 && x8 && x35 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && x63 && x64 && x55 && x33 && ~x32 && x8 && ~x35 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( x70 && x63 && x64 && x55 && x33 && ~x32 && ~x8 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( x70 && x63 && x64 && x55 && ~x33 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( x70 && x63 && x64 && ~x55 && x37 && x28 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( x70 && x63 && x64 && ~x55 && x37 && ~x28 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && x63 && x64 && ~x55 && ~x37 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s735;
						end
					else if( x70 && x63 && ~x64 && x15 && x2 && x8 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( x70 && x63 && ~x64 && x15 && x2 && x8 && ~x1 && x35 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && x63 && ~x64 && x15 && x2 && x8 && ~x1 && ~x35 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x70 && x63 && ~x64 && x15 && x2 && ~x8 && x32 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( x70 && x63 && ~x64 && x15 && x2 && ~x8 && x32 && ~x1 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x70 && x63 && ~x64 && x15 && x2 && ~x8 && x32 && ~x1 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( x70 && x63 && ~x64 && x15 && x2 && ~x8 && ~x32 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( x70 && x63 && ~x64 && x15 && ~x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( x70 && x63 && ~x64 && ~x15 && x37 && x28 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x70 && x63 && ~x64 && ~x15 && x37 && ~x28 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && x63 && ~x64 && ~x15 && ~x37 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s192;
						end
					else if( x70 && ~x63 && x64 && x40 && x2 && x8 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( x70 && ~x63 && x64 && x40 && x2 && x8 && ~x1 && x35 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && ~x63 && x64 && x40 && x2 && x8 && ~x1 && ~x35 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( x70 && ~x63 && x64 && x40 && x2 && ~x8 && x32 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( x70 && ~x63 && x64 && x40 && x2 && ~x8 && x32 && ~x1 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s736;
						end
					else if( x70 && ~x63 && x64 && x40 && x2 && ~x8 && x32 && ~x1 && ~x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s915;
						end
					else if( x70 && ~x63 && x64 && x40 && x2 && ~x8 && ~x32 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( x70 && ~x63 && x64 && x40 && ~x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && x64 && ~x40 && x37 && x28 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x70 && ~x63 && x64 && ~x40 && x37 && ~x28 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && ~x63 && x64 && ~x40 && ~x37 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x33 && x8 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x33 && x8 && ~x1 && x35 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x33 && x8 && ~x1 && ~x35 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s870;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x33 && ~x8 && x32 && x37 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s871;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x33 && ~x8 && x32 && ~x37 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s737;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x33 && ~x8 && x32 && ~x37 && ~x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s915;
						end
					else if( x70 && ~x63 && ~x64 && x44 && x33 && ~x8 && ~x32 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s870;
						end
					else if( x70 && ~x63 && ~x64 && x44 && ~x33 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && x1 && x28 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s867;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && x1 && ~x28 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x70 && ~x63 && ~x64 && ~x44 && ~x1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( ~x70 && x2 && x8 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x70 && x2 && x8 && ~x1 && x15 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x70 && x2 && x8 && ~x1 && ~x15 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x70 && x2 && ~x8 && x21 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x70 && x2 && ~x8 && x21 && ~x1 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( ~x70 && x2 && ~x8 && x21 && ~x1 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s444;
						end
					else if( ~x70 && x2 && ~x8 && ~x21 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x70 && ~x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else nx_state = s732;
				s733 : if( x70 && x61 && x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s875;
						end
					else if( x70 && x61 && ~x10 && x25 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( x70 && x61 && ~x10 && ~x25 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s842;
						end
					else if( x70 && ~x61 && x8 && x53 )
						begin
							y10 = 1'b1;	
							nx_state = s841;
						end
					else if( x70 && ~x61 && x8 && ~x53 && x37 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( x70 && ~x61 && x8 && ~x53 && ~x37 )
						begin
							y10 = 1'b1;	
							nx_state = s841;
						end
					else if( x70 && ~x61 && ~x8 && x51 )
						begin
							y10 = 1'b1;	
							nx_state = s841;
						end
					else if( x70 && ~x61 && ~x8 && ~x51 && x37 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( x70 && ~x61 && ~x8 && ~x51 && ~x37 )
						begin
							y10 = 1'b1;	
							nx_state = s841;
						end
					else if( ~x70 && x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x70 && ~x10 && x11 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s215;
						end
					else if( ~x70 && ~x10 && ~x11 && x12 && x8 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x70 && ~x10 && ~x11 && x12 && ~x8 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s280;
						end
					else if( ~x70 && ~x10 && ~x11 && ~x12 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s935;
						end
					else nx_state = s733;
				s734 : if( x55 && x16 && x50 && x33 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s908;
						end
					else if( x55 && x16 && x50 && ~x33 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x55 && x16 && x50 && ~x33 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x55 && x16 && ~x50 && x32 && x30 && x26 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s909;
						end
					else if( x55 && x16 && ~x50 && x32 && x30 && ~x26 && x34 )
						nx_state = s734;
					else if( x55 && x16 && ~x50 && x32 && x30 && ~x26 && ~x34 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s909;
						end
					else if( x55 && x16 && ~x50 && x32 && ~x30 )
						nx_state = s734;
					else if( x55 && x16 && ~x50 && ~x32 && x30 && x26 && x4 && x1 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s734;
						end
					else if( x55 && x16 && ~x50 && ~x32 && x30 && x26 && x4 && ~x1 )
						nx_state = s734;
					else if( x55 && x16 && ~x50 && ~x32 && x30 && x26 && ~x4 && x1 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s914;
						end
					else if( x55 && x16 && ~x50 && ~x32 && x30 && x26 && ~x4 && ~x1 )
						nx_state = s734;
					else if( x55 && x16 && ~x50 && ~x32 && x30 && ~x26 && x3 )
						nx_state = s734;
					else if( x55 && x16 && ~x50 && ~x32 && x30 && ~x26 && ~x3 && x4 && x1 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s734;
						end
					else if( x55 && x16 && ~x50 && ~x32 && x30 && ~x26 && ~x3 && x4 && ~x1 )
						nx_state = s734;
					else if( x55 && x16 && ~x50 && ~x32 && x30 && ~x26 && ~x3 && ~x4 && x1 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s914;
						end
					else if( x55 && x16 && ~x50 && ~x32 && x30 && ~x26 && ~x3 && ~x4 && ~x1 )
						nx_state = s734;
					else if( x55 && x16 && ~x50 && ~x32 && ~x30 )
						nx_state = s734;
					else if( x55 && ~x16 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( ~x55 && x28 && x57 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s735;
						end
					else if( ~x55 && x28 && ~x57 )
						nx_state = s734;
					else if( ~x55 && ~x28 && x27 && x8 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s735;
						end
					else if( ~x55 && ~x28 && x27 && ~x8 && x37 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( ~x55 && ~x28 && x27 && ~x8 && ~x37 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s908;
						end
					else if( ~x55 && ~x28 && ~x27 && x50 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x55 && ~x28 && ~x27 && ~x50 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s734;
						end
					else nx_state = s734;
				s735 : if( x55 && x41 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s914;
						end
					else if( x55 && ~x41 && x25 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s906;
						end
					else if( x55 && ~x41 && ~x25 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s910;
						end
					else if( ~x55 && x39 && x53 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s908;
						end
					else if( ~x55 && x39 && ~x53 && x37 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( ~x55 && x39 && ~x53 && ~x37 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s908;
						end
					else if( ~x55 && ~x39 && x51 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s908;
						end
					else if( ~x55 && ~x39 && ~x51 && x37 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( ~x55 && ~x39 && ~x51 && ~x37 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s908;
						end
					else nx_state = s735;
				s736 : if( x40 && x16 && x19 && x33 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( x40 && x16 && x19 && ~x33 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x40 && x16 && x19 && ~x33 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x40 && x16 && ~x19 && x30 && x26 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( x40 && x16 && ~x19 && x30 && x26 && ~x1 )
						nx_state = s736;
					else if( x40 && x16 && ~x19 && x30 && ~x26 && x3 )
						nx_state = s736;
					else if( x40 && x16 && ~x19 && x30 && ~x26 && ~x3 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( x40 && x16 && ~x19 && x30 && ~x26 && ~x3 && ~x1 )
						nx_state = s736;
					else if( x40 && x16 && ~x19 && ~x30 )
						nx_state = s736;
					else if( x40 && ~x16 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x40 && x28 && x43 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( ~x40 && x28 && ~x43 )
						nx_state = s736;
					else if( ~x40 && ~x28 && x27 && x8 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( ~x40 && ~x28 && x27 && ~x8 && x37 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x40 && ~x28 && x27 && ~x8 && ~x37 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( ~x40 && ~x28 && ~x27 && x50 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x40 && ~x28 && ~x27 && ~x50 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s736;
						end
					else nx_state = s736;
				s737 : if( x44 && x16 && x19 && x33 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( x44 && x16 && x19 && ~x33 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x44 && x16 && x19 && ~x33 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x44 && x16 && ~x19 && x30 && x26 && x1 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s871;
						end
					else if( x44 && x16 && ~x19 && x30 && x26 && ~x1 && x37 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s737;
						end
					else if( x44 && x16 && ~x19 && x30 && x26 && ~x1 && x37 && ~x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s915;
						end
					else if( x44 && x16 && ~x19 && x30 && x26 && ~x1 && ~x37 )
						nx_state = s737;
					else if( x44 && x16 && ~x19 && x30 && ~x26 && x1 && x3 )
						nx_state = s737;
					else if( x44 && x16 && ~x19 && x30 && ~x26 && x1 && ~x3 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s871;
						end
					else if( x44 && x16 && ~x19 && x30 && ~x26 && ~x1 && x37 && x43 )
						nx_state = s737;
					else if( x44 && x16 && ~x19 && x30 && ~x26 && ~x1 && x37 && ~x43 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s737;
						end
					else if( x44 && x16 && ~x19 && x30 && ~x26 && ~x1 && x37 && ~x43 && ~x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s915;
						end
					else if( x44 && x16 && ~x19 && x30 && ~x26 && ~x1 && ~x37 )
						nx_state = s737;
					else if( x44 && x16 && ~x19 && ~x30 )
						nx_state = s737;
					else if( x44 && ~x16 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x44 && x28 && x49 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( ~x44 && x28 && ~x49 )
						nx_state = s737;
					else if( ~x44 && ~x28 && x27 && x8 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( ~x44 && ~x28 && x27 && ~x8 && x36 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x44 && ~x28 && x27 && ~x8 && ~x36 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( ~x44 && ~x28 && ~x27 && x50 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s867;
						end
					else if( ~x44 && ~x28 && ~x27 && ~x50 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s737;
						end
					else nx_state = s737;
				s738 : if( x69 )
						nx_state = s47;
					else if( ~x69 && x70 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && x70 && ~x1 && x62 && x35 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s840;
						end
					else if( ~x69 && x70 && ~x1 && x62 && ~x35 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( ~x69 && x70 && ~x1 && ~x62 && x35 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && x70 && ~x1 && ~x62 && ~x35 && x63 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && x70 && ~x1 && ~x62 && ~x35 && ~x63 && x64 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( ~x69 && x70 && ~x1 && ~x62 && ~x35 && ~x63 && ~x64 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s870;
						end
					else if( ~x69 && ~x70 && x44 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && ~x70 && x44 && ~x1 && x15 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && ~x70 && x44 && ~x1 && ~x15 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x70 && ~x44 && x10 && x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && ~x70 && ~x44 && x10 && ~x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 && ~x1 && x3 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( ~x69 && ~x70 && ~x44 && ~x10 && ~x1 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else nx_state = s738;
				s739 : if( x32 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s739;
						end
					else if( ~x32 && x35 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x32 && ~x35 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else nx_state = s739;
				s740 : if( x10 && x8 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( x10 && ~x8 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s280;
						end
					else if( ~x10 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s215;
						end
					else nx_state = s740;
				s741 : if( x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x6 && ~x5 )
						nx_state = s1;
					else nx_state = s741;
				s742 : if( x11 )
						begin
							y21 = 1'b1;	
							nx_state = s822;
						end
					else if( ~x11 && x22 && x9 && x8 && x23 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x11 && x22 && x9 && x8 && x23 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x11 && x22 && x9 && x8 && x23 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x11 && x22 && x9 && x8 && x23 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x11 && x22 && x9 && x8 && x23 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x11 && x22 && x9 && x8 && ~x23 && x10 )
						begin
							y62 = 1'b1;	
							nx_state = s1120;
						end
					else if( ~x11 && x22 && x9 && x8 && ~x23 && ~x10 )
						begin
							y61 = 1'b1;	
							nx_state = s1098;
						end
					else if( ~x11 && x22 && x9 && ~x8 && x23 && x10 && x5 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( ~x11 && x22 && x9 && ~x8 && x23 && x10 && ~x5 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x11 && x22 && x9 && ~x8 && x23 && x10 && ~x5 && x6 && ~x4 )
						nx_state = s1;
					else if( ~x11 && x22 && x9 && ~x8 && x23 && x10 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x11 && x22 && x9 && ~x8 && x23 && ~x10 && x4 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( ~x11 && x22 && x9 && ~x8 && x23 && ~x10 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x11 && x22 && x9 && ~x8 && x23 && ~x10 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x11 && x22 && x9 && ~x8 && ~x23 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y38 = 1'b1;	
							y63 = 1'b1;	
							nx_state = s741;
						end
					else if( ~x11 && x22 && x9 && ~x8 && ~x23 && ~x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y36 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s741;
						end
					else if( ~x11 && x22 && ~x9 && x10 && x23 && x8 )
						begin
							y33 = 1'b1;	y54 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x11 && x22 && ~x9 && x10 && x23 && ~x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y26 = 1'b1;	
							y51 = 1'b1;	y56 = 1'b1;	
							nx_state = s741;
						end
					else if( ~x11 && x22 && ~x9 && x10 && ~x23 && x8 )
						begin
							y60 = 1'b1;	
							nx_state = s424;
						end
					else if( ~x11 && x22 && ~x9 && x10 && ~x23 && ~x8 )
						begin
							y58 = 1'b1;	
							nx_state = s1265;
						end
					else if( ~x11 && x22 && ~x9 && ~x10 && x23 && x8 )
						begin
							y37 = 1'b1;	y55 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x11 && x22 && ~x9 && ~x10 && x23 && ~x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y23 = 1'b1;	
							y52 = 1'b1;	y53 = 1'b1;	
							nx_state = s741;
						end
					else if( ~x11 && x22 && ~x9 && ~x10 && ~x23 && x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y23 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1266;
						end
					else if( ~x11 && x22 && ~x9 && ~x10 && ~x23 && ~x8 )
						begin
							y56 = 1'b1;	
							nx_state = s1219;
						end
					else if( ~x11 && ~x22 && x23 && x21 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( ~x11 && ~x22 && x23 && ~x21 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s1267;
						end
					else if( ~x11 && ~x22 && ~x23 && x9 && x10 && x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y38 = 1'b1;	
							y46 = 1'b1;	
							nx_state = s741;
						end
					else if( ~x11 && ~x22 && ~x23 && x9 && x10 && ~x8 )
						begin
							y5 = 1'b1;	y34 = 1'b1;	y36 = 1'b1;	
							y38 = 1'b1;	y40 = 1'b1;	
							nx_state = s741;
						end
					else if( ~x11 && ~x22 && ~x23 && x9 && ~x10 && x8 )
						begin
							y47 = 1'b1;	
							nx_state = s287;
						end
					else if( ~x11 && ~x22 && ~x23 && x9 && ~x10 && ~x8 )
						begin
							y5 = 1'b1;	y34 = 1'b1;	y36 = 1'b1;	
							y38 = 1'b1;	y39 = 1'b1;	
							nx_state = s741;
						end
					else if( ~x11 && ~x22 && ~x23 && ~x9 && x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y42 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s1042;
						end
					else if( ~x11 && ~x22 && ~x23 && ~x9 && ~x8 )
						begin
							y5 = 1'b1;	y34 = 1'b1;	y35 = 1'b1;	
							y36 = 1'b1;	y38 = 1'b1;	
							nx_state = s741;
						end
					else nx_state = s742;
				s743 : if( x63 && x12 && x22 )
						begin
							y6 = 1'b1;	
							nx_state = s431;
						end
					else if( x63 && x12 && ~x22 && x23 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x63 && x12 && ~x22 && ~x23 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( x63 && ~x12 && x7 && x22 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1100;
						end
					else if( x63 && ~x12 && x7 && ~x22 && x8 && x9 && x23 && x10 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y5 = 1'b1;	
							y22 = 1'b1;	y23 = 1'b1;	
							nx_state = s72;
						end
					else if( x63 && ~x12 && x7 && ~x22 && x8 && x9 && x23 && ~x10 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( x63 && ~x12 && x7 && ~x22 && x8 && x9 && ~x23 && x10 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y38 = 1'b1;	
							y46 = 1'b1;	
							nx_state = s741;
						end
					else if( x63 && ~x12 && x7 && ~x22 && x8 && x9 && ~x23 && ~x10 )
						begin
							y47 = 1'b1;	
							nx_state = s287;
						end
					else if( x63 && ~x12 && x7 && ~x22 && x8 && ~x9 && x23 && x10 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( x63 && ~x12 && x7 && ~x22 && x8 && ~x9 && x23 && x10 && ~x13 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x12 && x7 && ~x22 && x8 && ~x9 && x23 && x10 && ~x13 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x12 && x7 && ~x22 && x8 && ~x9 && x23 && x10 && ~x13 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x63 && ~x12 && x7 && ~x22 && x8 && ~x9 && x23 && x10 && ~x13 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x12 && x7 && ~x22 && x8 && ~x9 && x23 && x10 && ~x13 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x63 && ~x12 && x7 && ~x22 && x8 && ~x9 && x23 && ~x10 && x1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( x63 && ~x12 && x7 && ~x22 && x8 && ~x9 && x23 && ~x10 && ~x1 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x12 && x7 && ~x22 && x8 && ~x9 && x23 && ~x10 && ~x1 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x12 && x7 && ~x22 && x8 && ~x9 && x23 && ~x10 && ~x1 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x63 && ~x12 && x7 && ~x22 && x8 && ~x9 && x23 && ~x10 && ~x1 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x12 && x7 && ~x22 && x8 && ~x9 && x23 && ~x10 && ~x1 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x63 && ~x12 && x7 && ~x22 && x8 && ~x9 && ~x23 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y42 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s1042;
						end
					else if( x63 && ~x12 && x7 && ~x22 && ~x8 && x9 && x23 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( x63 && ~x12 && x7 && ~x22 && ~x8 && x9 && ~x23 && x10 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y38 = 1'b1;	
							y40 = 1'b1;	y41 = 1'b1;	
							nx_state = s741;
						end
					else if( x63 && ~x12 && x7 && ~x22 && ~x8 && x9 && ~x23 && ~x10 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y38 = 1'b1;	
							y39 = 1'b1;	y41 = 1'b1;	
							nx_state = s741;
						end
					else if( x63 && ~x12 && x7 && ~x22 && ~x8 && ~x9 && x23 && x10 && x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( x63 && ~x12 && x7 && ~x22 && ~x8 && ~x9 && x23 && x10 && ~x3 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x12 && x7 && ~x22 && ~x8 && ~x9 && x23 && x10 && ~x3 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x12 && x7 && ~x22 && ~x8 && ~x9 && x23 && x10 && ~x3 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x63 && ~x12 && x7 && ~x22 && ~x8 && ~x9 && x23 && x10 && ~x3 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x12 && x7 && ~x22 && ~x8 && ~x9 && x23 && x10 && ~x3 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x63 && ~x12 && x7 && ~x22 && ~x8 && ~x9 && x23 && ~x10 && x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( x63 && ~x12 && x7 && ~x22 && ~x8 && ~x9 && x23 && ~x10 && ~x15 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x12 && x7 && ~x22 && ~x8 && ~x9 && x23 && ~x10 && ~x15 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x12 && x7 && ~x22 && ~x8 && ~x9 && x23 && ~x10 && ~x15 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x63 && ~x12 && x7 && ~x22 && ~x8 && ~x9 && x23 && ~x10 && ~x15 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x12 && x7 && ~x22 && ~x8 && ~x9 && x23 && ~x10 && ~x15 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x63 && ~x12 && x7 && ~x22 && ~x8 && ~x9 && ~x23 )
						begin
							y5 = 1'b1;	y35 = 1'b1;	y36 = 1'b1;	
							y38 = 1'b1;	y41 = 1'b1;	
							nx_state = s741;
						end
					else if( x63 && ~x12 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s523;
						end
					else if( ~x63 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1268;
						end
					else if( ~x63 && ~x15 && x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s1269;
						end
					else if( ~x63 && ~x15 && ~x16 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s1270;
						end
					else nx_state = s743;
				s744 : if( x64 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y62 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s425;
						end
					else if( ~x64 )
						begin
							y47 = 1'b1;	y57 = 1'b1;	y61 = 1'b1;	
							y71 = 1'b1;	
							nx_state = s1271;
						end
					else nx_state = s744;
				s745 : if( x45 && x13 )
						begin
							y3 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s883;
						end
					else if( x45 && ~x13 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s1182;
						end
					else if( ~x45 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y27 = 1'b1;	
							nx_state = s696;
						end
					else nx_state = s745;
				s746 : if( x63 && x66 && x23 && x25 )
						begin
							y57 = 1'b1;	
							nx_state = s1223;
						end
					else if( x63 && x66 && x23 && ~x25 && x5 )
						begin
							y61 = 1'b1;	
							nx_state = s1098;
						end
					else if( x63 && x66 && x23 && ~x25 && ~x5 )
						begin
							y57 = 1'b1;	
							nx_state = s1223;
						end
					else if( x63 && x66 && ~x23 && x5 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x63 && x66 && ~x23 && x5 && ~x24 )
						begin
							y60 = 1'b1;	
							nx_state = s424;
						end
					else if( x63 && x66 && ~x23 && ~x5 )
						begin
							y53 = 1'b1;	
							nx_state = s1071;
						end
					else if( x63 && ~x66 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x63 && ~x66 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x63 && ~x66 && x19 && ~x14 && ~x13 && x11 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( x63 && ~x66 && x19 && ~x14 && ~x13 && x11 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( x63 && ~x66 && x19 && ~x14 && ~x13 && ~x11 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( x63 && ~x66 && ~x19 )
						nx_state = s1;
					else if( ~x63 && x64 && x66 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x63 && x64 && x66 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x63 && x64 && x66 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x63 && x64 && x66 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x63 && x64 && x66 && ~x22 )
						nx_state = s1;
					else if( ~x63 && x64 && ~x66 )
						nx_state = s1;
					else if( ~x63 && ~x64 )
						begin
							y57 = 1'b1;	
							nx_state = s1223;
						end
					else nx_state = s746;
				s747 : if( x70 && x62 )
						begin
							y8 = 1'b1;	
							nx_state = s568;
						end
					else if( x70 && ~x62 && x65 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x70 && ~x62 && ~x65 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x70 && x65 && x66 )
						nx_state = s331;
					else if( ~x70 && x65 && ~x66 && x67 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( ~x70 && x65 && ~x66 && x67 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( ~x70 && x65 && ~x66 && x67 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && x67 && ~x8 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x19 && x18 && x14 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	y25 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x19 && x18 && ~x14 && x17 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	y25 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x19 && x18 && ~x14 && ~x17 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x19 && x18 && ~x14 && ~x17 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && x19 && x18 && ~x14 && ~x17 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x19 && x18 && ~x14 && ~x17 && ~x5 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && x19 && ~x18 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	y25 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x19 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x19 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x19 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x70 && x65 && ~x66 && ~x67 && ~x19 && ~x5 )
						nx_state = s1;
					else if( ~x70 && ~x65 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else nx_state = s747;
				s748 : if( x65 )
						begin
							y8 = 1'b1;	
							nx_state = s373;
						end
					else if( ~x65 )
						begin
							y7 = 1'b1;	
							nx_state = s1272;
						end
					else nx_state = s748;
				s749 : if( x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x18 )
						nx_state = s1;
					else nx_state = s749;
				s750 : if( x6 && x12 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s1273;
						end
					else if( x6 && ~x12 && x11 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s1008;
						end
					else if( x6 && ~x12 && ~x11 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x6 && ~x12 && ~x11 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x6 && ~x12 && ~x11 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x6 && ~x12 && ~x11 && ~x18 )
						nx_state = s1;
					else if( ~x6 && x8 && x11 && x12 && x10 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x6 && x8 && x11 && x12 && x10 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x6 && x8 && x11 && x12 && x10 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x6 && x8 && x11 && x12 && x10 && ~x18 )
						nx_state = s1;
					else if( ~x6 && x8 && x11 && x12 && ~x10 && x16 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s749;
						end
					else if( ~x6 && x8 && x11 && x12 && ~x10 && ~x16 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x6 && x8 && x11 && x12 && ~x10 && ~x16 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x6 && x8 && x11 && x12 && ~x10 && ~x16 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x6 && x8 && x11 && x12 && ~x10 && ~x16 && ~x18 )
						nx_state = s1;
					else if( ~x6 && x8 && x11 && ~x12 && x10 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s1274;
						end
					else if( ~x6 && x8 && x11 && ~x12 && ~x10 && x17 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s749;
						end
					else if( ~x6 && x8 && x11 && ~x12 && ~x10 && ~x17 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x6 && x8 && x11 && ~x12 && ~x10 && ~x17 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x6 && x8 && x11 && ~x12 && ~x10 && ~x17 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x6 && x8 && x11 && ~x12 && ~x10 && ~x17 && ~x18 )
						nx_state = s1;
					else if( ~x6 && x8 && ~x11 && x12 && x10 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y34 = 1'b1;	
							nx_state = s1275;
						end
					else if( ~x6 && x8 && ~x11 && x12 && ~x10 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s749;
						end
					else if( ~x6 && x8 && ~x11 && ~x12 && x10 && x15 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s749;
						end
					else if( ~x6 && x8 && ~x11 && ~x12 && x10 && ~x15 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x6 && x8 && ~x11 && ~x12 && x10 && ~x15 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x6 && x8 && ~x11 && ~x12 && x10 && ~x15 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x6 && x8 && ~x11 && ~x12 && x10 && ~x15 && ~x18 )
						nx_state = s1;
					else if( ~x6 && x8 && ~x11 && ~x12 && ~x10 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x6 && ~x8 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s1273;
						end
					else nx_state = s750;
				s751 : if( x62 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x62 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x62 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( x62 && ~x21 )
						nx_state = s1;
					else if( ~x62 && x63 && x16 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x62 && x63 && x16 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x62 && x63 && x16 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x62 && x63 && ~x16 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && x66 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x62 && ~x63 && x64 && x66 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x62 && ~x63 && x64 && x66 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && x66 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && x66 && ~x22 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && ~x66 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x62 && ~x63 && x64 && ~x66 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x62 && ~x63 && x64 && ~x66 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && ~x66 && ~x18 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 && x65 )
						begin
							y47 = 1'b1;	y49 = 1'b1;	y58 = 1'b1;	
							y61 = 1'b1;	y70 = 1'b1;	
							nx_state = s1276;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 && ~x65 && ~x8 )
						nx_state = s1;
					else nx_state = s751;
				s752 : if( 1'b1 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y33 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1277;
						end
					else nx_state = s752;
				s753 : if( x62 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x62 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x62 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( x62 && ~x21 )
						nx_state = s1;
					else if( ~x62 && x64 && x63 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x63 && x65 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x63 && ~x65 && x66 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && x64 && ~x63 && ~x65 && x66 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && x64 && ~x63 && ~x65 && x66 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x63 && ~x65 && x66 && ~x9 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x63 && ~x65 && ~x66 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x62 && x64 && ~x63 && ~x65 && ~x66 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x62 && x64 && ~x63 && ~x65 && ~x66 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x63 && ~x65 && ~x66 && ~x18 )
						nx_state = s1;
					else if( ~x62 && ~x64 && x63 && x16 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x62 && ~x64 && x63 && x16 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x62 && ~x64 && x63 && x16 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x62 && ~x64 && x63 && ~x16 )
						nx_state = s1;
					else if( ~x62 && ~x64 && ~x63 && x65 )
						begin
							y25 = 1'b1;	
							nx_state = s1157;
						end
					else if( ~x62 && ~x64 && ~x63 && ~x65 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x62 && ~x64 && ~x63 && ~x65 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x62 && ~x64 && ~x63 && ~x65 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x62 && ~x64 && ~x63 && ~x65 && ~x8 )
						nx_state = s1;
					else nx_state = s753;
				s754 : if( x62 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x62 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x62 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( x62 && ~x21 )
						nx_state = s1;
					else if( ~x62 && x63 && x11 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x62 && x63 && x11 && ~x18 )
						begin
							y44 = 1'b1;	y45 = 1'b1;	
							nx_state = s392;
						end
					else if( ~x62 && x63 && ~x11 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( ~x62 && ~x63 && x64 && x66 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && ~x63 && x64 && x66 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && ~x63 && x64 && x66 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && x66 && ~x9 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && ~x66 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x62 && ~x63 && x64 && ~x66 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x62 && ~x63 && x64 && ~x66 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && ~x66 && ~x18 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 && x30 && x4 && x9 && x10 && x8 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x62 && ~x63 && ~x64 && x30 && x4 && x9 && x10 && ~x8 )
						begin
							y8 = 1'b1;	
							nx_state = s784;
						end
					else if( ~x62 && ~x63 && ~x64 && x30 && x4 && x9 && ~x10 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x62 && ~x63 && ~x64 && x30 && x4 && x9 && ~x10 && ~x8 )
						begin
							y8 = 1'b1;	
							nx_state = s785;
						end
					else if( ~x62 && ~x63 && ~x64 && x30 && x4 && ~x9 && x10 && x8 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x62 && ~x63 && ~x64 && x30 && x4 && ~x9 && x10 && ~x8 && x27 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( ~x62 && ~x63 && ~x64 && x30 && x4 && ~x9 && x10 && ~x8 && ~x27 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x62 && ~x63 && ~x64 && x30 && x4 && ~x9 && ~x10 && x8 )
						begin
							y8 = 1'b1;	
							nx_state = s786;
						end
					else if( ~x62 && ~x63 && ~x64 && x30 && x4 && ~x9 && ~x10 && ~x8 && x26 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x62 && ~x63 && ~x64 && x30 && x4 && ~x9 && ~x10 && ~x8 && ~x26 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( ~x62 && ~x63 && ~x64 && x30 && ~x4 )
						begin
							y5 = 1'b1;	
							nx_state = s950;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && x9 && x10 && x8 )
						begin
							y9 = 1'b1;	
							nx_state = s790;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && x9 && x10 && ~x8 && x21 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && x9 && x10 && ~x8 && ~x21 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && x9 && x10 && ~x8 && ~x21 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && x9 && x10 && ~x8 && ~x21 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && x9 && x10 && ~x8 && ~x21 && ~x23 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && x9 && ~x10 && x8 )
						begin
							y3 = 1'b1;	
							nx_state = s789;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && x9 && ~x10 && ~x8 && x18 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && x9 && ~x10 && ~x8 && ~x18 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && x9 && ~x10 && ~x8 && ~x18 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && x9 && ~x10 && ~x8 && ~x18 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && x9 && ~x10 && ~x8 && ~x18 && ~x23 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && ~x9 && x8 && x10 && x19 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && ~x9 && x8 && x10 && ~x19 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && ~x9 && x8 && x10 && ~x19 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && ~x9 && x8 && x10 && ~x19 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && ~x9 && x8 && x10 && ~x19 && ~x23 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && ~x9 && x8 && ~x10 && x20 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && ~x9 && x8 && ~x10 && ~x20 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && ~x9 && x8 && ~x10 && ~x20 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && ~x9 && x8 && ~x10 && ~x20 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && ~x9 && x8 && ~x10 && ~x20 && ~x23 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && x31 && ~x9 && ~x8 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x30 && x4 && ~x31 )
						begin
							y9 = 1'b1;	
							nx_state = s790;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x30 && ~x4 && x31 )
						begin
							y5 = 1'b1;	
							nx_state = s560;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x30 && ~x4 && ~x31 )
						begin
							y5 = 1'b1;	
							nx_state = s791;
						end
					else nx_state = s754;
				s755 : if( x63 && x66 && x19 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( x63 && x66 && ~x19 )
						begin
							y45 = 1'b1;	
							nx_state = s286;
						end
					else if( x63 && ~x66 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1278;
						end
					else if( ~x63 && x65 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							nx_state = s1279;
						end
					else if( ~x63 && ~x65 && x66 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && ~x65 && x66 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && ~x65 && x66 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x63 && ~x65 && x66 && ~x9 )
						nx_state = s1;
					else if( ~x63 && ~x65 && ~x66 && x67 && x17 )
						begin
							y48 = 1'b1;	
							nx_state = s1009;
						end
					else if( ~x63 && ~x65 && ~x66 && x67 && ~x17 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x63 && ~x65 && ~x66 && x67 && ~x17 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x63 && ~x65 && ~x66 && x67 && ~x17 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( ~x63 && ~x65 && ~x66 && x67 && ~x17 && ~x14 )
						nx_state = s1;
					else if( ~x63 && ~x65 && ~x66 && ~x67 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x63 && ~x65 && ~x66 && ~x67 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x63 && ~x65 && ~x66 && ~x67 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x63 && ~x65 && ~x66 && ~x67 && ~x18 )
						nx_state = s1;
					else nx_state = s755;
				s756 : if( x11 && x12 && x10 )
						begin
							y47 = 1'b1;	
							nx_state = s675;
						end
					else if( x11 && x12 && ~x10 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y29 = 1'b1;	
							y35 = 1'b1;	y36 = 1'b1;	
							nx_state = s749;
						end
					else if( x11 && ~x12 && x10 )
						begin
							y48 = 1'b1;	
							nx_state = s1009;
						end
					else if( x11 && ~x12 && ~x10 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y30 = 1'b1;	
							y35 = 1'b1;	y36 = 1'b1;	
							nx_state = s749;
						end
					else if( ~x11 && x12 && x10 )
						begin
							y56 = 1'b1;	
							nx_state = s1007;
						end
					else if( ~x11 && x12 && ~x10 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y28 = 1'b1;	
							y35 = 1'b1;	y36 = 1'b1;	
							nx_state = s749;
						end
					else if( ~x11 && ~x12 && x10 )
						begin
							y54 = 1'b1;	
							nx_state = s525;
						end
					else if( ~x11 && ~x12 && ~x10 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x11 && ~x12 && ~x10 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x11 && ~x12 && ~x10 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x11 && ~x12 && ~x10 && ~x18 )
						nx_state = s1;
					else nx_state = s756;
				s757 : if( x7 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else nx_state = s757;
				s758 : if( x21 && x20 && x16 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s233;
						end
					else if( x21 && x20 && x16 && ~x10 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x21 && x20 && ~x16 && x17 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x21 && x20 && ~x16 && ~x17 )
						begin
							y5 = 1'b1;	y17 = 1'b1;	
							nx_state = s721;
						end
					else if( x21 && ~x20 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( ~x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else nx_state = s758;
				s759 : if( x69 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s131;
						end
					else if( ~x69 && x8 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s206;
						end
					else if( ~x69 && x8 && ~x1 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s934;
						end
					else if( ~x69 && x8 && ~x1 && ~x4 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && ~x8 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else nx_state = s759;
				s760 : if( x69 && x21 && x20 )
						begin
							y13 = 1'b1;	y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s1;
						end
					else if( x69 && x21 && ~x20 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x69 && x21 && ~x20 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x69 && x21 && ~x20 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x69 && x21 && ~x20 && ~x10 )
						nx_state = s1;
					else if( x69 && ~x21 )
						begin
							y13 = 1'b1;	y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x69 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x69 && ~x1 && x70 && x62 && x35 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s840;
						end
					else if( ~x69 && ~x1 && x70 && x62 && ~x35 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( ~x69 && ~x1 && x70 && ~x62 && x35 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && ~x1 && x70 && ~x62 && ~x35 && x63 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x1 && x70 && ~x62 && ~x35 && ~x63 && x64 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( ~x69 && ~x1 && x70 && ~x62 && ~x35 && ~x63 && ~x64 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s870;
						end
					else if( ~x69 && ~x1 && ~x70 && x44 && x45 && x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( ~x69 && ~x1 && ~x70 && x44 && x45 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x1 && ~x70 && x44 && ~x45 && x15 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && ~x1 && ~x70 && x44 && ~x45 && ~x15 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x69 && ~x1 && ~x70 && ~x44 && x3 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( ~x69 && ~x1 && ~x70 && ~x44 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else nx_state = s760;
				s761 : if( x69 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else if( ~x69 && x15 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s1280;
						end
					else if( ~x69 && ~x15 && x5 )
						begin
							y2 = 1'b1;	
							nx_state = s768;
						end
					else if( ~x69 && ~x15 && ~x5 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s1280;
						end
					else nx_state = s761;
				s762 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s816;
						end
					else nx_state = s762;
				s763 : if( x69 && x62 && x17 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y37 = 1'b1;	
							nx_state = s1204;
						end
					else if( x69 && x62 && ~x17 )
						begin
							y1 = 1'b1;	y21 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s580;
						end
					else if( x69 && ~x62 )
						begin
							y13 = 1'b1;	
							nx_state = s1281;
						end
					else if( ~x69 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s1233;
						end
					else nx_state = s763;
				s764 : if( x69 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x69 && x15 && x13 )
						begin
							y13 = 1'b1;	
							nx_state = s769;
						end
					else if( ~x69 && x15 && ~x13 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s1282;
						end
					else if( ~x69 && ~x15 && x12 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s1282;
						end
					else if( ~x69 && ~x15 && ~x12 )
						nx_state = s764;
					else nx_state = s764;
				s765 : if( x15 && x14 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s1283;
						end
					else if( x15 && ~x14 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s764;
						end
					else if( ~x15 && x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s817;
						end
					else if( ~x15 && ~x12 )
						nx_state = s765;
					else nx_state = s765;
				s766 : if( x69 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	y26 = 1'b1;	
							nx_state = s926;
						end
					else if( ~x69 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s817;
						end
					else if( ~x69 && ~x15 && x6 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s1283;
						end
					else if( ~x69 && ~x15 && ~x6 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s765;
						end
					else nx_state = s766;
				s767 : if( x15 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s1284;
						end
					else if( ~x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s216;
						end
					else nx_state = s767;
				s768 : if( x69 && x63 && x19 && x18 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1094;
						end
					else if( x69 && x63 && x19 && ~x18 )
						begin
							y25 = 1'b1;	y28 = 1'b1;	y48 = 1'b1;	
							nx_state = s1285;
						end
					else if( x69 && x63 && ~x19 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1286;
						end
					else if( x69 && ~x63 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y20 = 1'b1;	
							nx_state = s1287;
						end
					else if( ~x69 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s216;
						end
					else if( ~x69 && ~x15 && x6 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x69 && ~x15 && ~x6 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s770;
						end
					else nx_state = s768;
				s769 : if( x69 && x62 && x17 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y9 = 1'b1;	
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s1288;
						end
					else if( x69 && x62 && ~x17 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1018;
						end
					else if( x69 && ~x62 && x64 )
						begin
							y47 = 1'b1;	y48 = 1'b1;	
							nx_state = s1289;
						end
					else if( x69 && ~x62 && ~x64 )
						begin
							y13 = 1'b1;	
							nx_state = s897;
						end
					else if( ~x69 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s216;
						end
					else if( ~x69 && ~x15 && x11 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s767;
						end
					else if( ~x69 && ~x15 && ~x11 && x10 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s428;
						end
					else if( ~x69 && ~x15 && ~x11 && ~x10 )
						nx_state = s769;
					else nx_state = s769;
				s770 : if( x15 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x15 && x8 )
						begin
							y13 = 1'b1;	
							nx_state = s769;
						end
					else if( ~x15 && ~x8 && x9 )
						begin
							y13 = 1'b1;	
							nx_state = s769;
						end
					else if( ~x15 && ~x8 && ~x9 && x10 && x6 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x15 && ~x8 && ~x9 && x10 && ~x6 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s770;
						end
					else if( ~x15 && ~x8 && ~x9 && ~x10 && x11 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s767;
						end
					else if( ~x15 && ~x8 && ~x9 && ~x10 && ~x11 )
						nx_state = s770;
					else nx_state = s770;
				s771 : if( x64 && x62 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x64 && x62 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x64 && x62 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x64 && x62 && ~x10 )
						nx_state = s1;
					else if( x64 && ~x62 && x63 && x65 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s1290;
						end
					else if( x64 && ~x62 && x63 && ~x65 && x21 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x64 && ~x62 && x63 && ~x65 && x21 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x64 && ~x62 && x63 && ~x65 && x21 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x64 && ~x62 && x63 && ~x65 && x21 && ~x10 )
						nx_state = s1;
					else if( x64 && ~x62 && x63 && ~x65 && ~x21 )
						begin
							y13 = 1'b1;	
							nx_state = s769;
						end
					else if( x64 && ~x62 && ~x63 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x64 && ~x62 && ~x63 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x64 && ~x62 && ~x63 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x64 && ~x62 && ~x63 && ~x14 )
						nx_state = s1;
					else if( ~x64 && x62 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x64 && x62 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x64 && x62 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( ~x64 && x62 && ~x27 )
						nx_state = s1;
					else if( ~x64 && ~x62 && x63 && x66 && x14 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( ~x64 && ~x62 && x63 && x66 && x14 && ~x15 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x64 && ~x62 && x63 && x66 && ~x14 )
						begin
							y30 = 1'b1;	
							nx_state = s291;
						end
					else if( ~x64 && ~x62 && x63 && ~x66 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( ~x64 && ~x62 && x63 && ~x66 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( ~x64 && ~x62 && x63 && ~x66 && x19 && ~x14 && ~x13 && x11 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( ~x64 && ~x62 && x63 && ~x66 && x19 && ~x14 && ~x13 && x11 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x64 && ~x62 && x63 && ~x66 && x19 && ~x14 && ~x13 && ~x11 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x64 && ~x62 && x63 && ~x66 && ~x19 )
						nx_state = s1;
					else if( ~x64 && ~x62 && ~x63 && x65 && x67 )
						begin
							y30 = 1'b1;	
							nx_state = s291;
						end
					else if( ~x64 && ~x62 && ~x63 && x65 && ~x67 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x64 && ~x62 && ~x63 && x65 && ~x67 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x64 && ~x62 && ~x63 && x65 && ~x67 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x64 && ~x62 && ~x63 && x65 && ~x67 && ~x23 )
						nx_state = s1;
					else if( ~x64 && ~x62 && ~x63 && ~x65 && x21 && x22 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x64 && ~x62 && ~x63 && ~x65 && x21 && ~x22 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x64 && ~x62 && ~x63 && ~x65 && x21 && ~x22 && ~x23 )
						nx_state = s1;
					else if( ~x64 && ~x62 && ~x63 && ~x65 && ~x21 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x64 && ~x62 && ~x63 && ~x65 && ~x21 && ~x23 )
						nx_state = s1;
					else nx_state = s771;
				s772 : if( x63 && x64 )
						begin
							y13 = 1'b1;	
							nx_state = s450;
						end
					else if( x63 && ~x64 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x63 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x63 && ~x9 )
						nx_state = s1;
					else nx_state = s772;
				s773 : if( x63 )
						begin
							y6 = 1'b1;	y17 = 1'b1;	y22 = 1'b1;	
							y46 = 1'b1;	y47 = 1'b1;	
							nx_state = s1291;
						end
					else if( ~x63 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x63 && ~x9 )
						nx_state = s1;
					else nx_state = s773;
				s774 : if( x13 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x13 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x13 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x13 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x13 && ~x9 )
						nx_state = s1;
					else nx_state = s774;
				s775 : if( x63 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x63 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x63 && x19 && ~x14 && ~x13 && x11 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( x63 && x19 && ~x14 && ~x13 && x11 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( x63 && x19 && ~x14 && ~x13 && ~x11 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( x63 && ~x19 )
						nx_state = s1;
					else if( ~x63 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x63 && ~x9 )
						nx_state = s1;
					else nx_state = s775;
				s776 : if( x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x21 && ~x20 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x19 )
						nx_state = s1;
					else nx_state = s776;
				s777 : if( x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x21 && ~x20 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( ~x21 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else nx_state = s777;
				s778 : if( 1'b1 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s1292;
						end
					else nx_state = s778;
				s779 : if( x10 && x12 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( x10 && ~x12 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x10 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else nx_state = s779;
				s780 : if( x20 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x20 && ~x15 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s131;
						end
					else if( ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else nx_state = s780;
				s781 : if( x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x20 && ~x18 )
						nx_state = s1;
					else if( ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s407;
						end
					else if( ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else nx_state = s781;
				s782 : if( x1 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	
							nx_state = s813;
						end
					else if( ~x1 && x17 && x15 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s556;
						end
					else if( ~x1 && x17 && ~x15 && x16 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s131;
						end
					else if( ~x1 && x17 && ~x15 && ~x16 )
						begin
							y7 = 1'b1;	y12 = 1'b1;	
							nx_state = s610;
						end
					else if( ~x1 && ~x17 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	y22 = 1'b1;	
							nx_state = s1070;
						end
					else nx_state = s782;
				s783 : if( x69 && x64 && x3 )
						begin
							y3 = 1'b1;	
							nx_state = s1293;
						end
					else if( x69 && x64 && ~x3 && x20 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( x69 && x64 && ~x3 && ~x20 && x21 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x69 && x64 && ~x3 && ~x20 && ~x21 )
						begin
							y31 = 1'b1;	
							nx_state = s164;
						end
					else if( x69 && ~x64 && x31 )
						begin
							y47 = 1'b1;	y53 = 1'b1;	y61 = 1'b1;	
							y69 = 1'b1;	
							nx_state = s982;
						end
					else if( x69 && ~x64 && ~x31 )
						begin
							y47 = 1'b1;	y49 = 1'b1;	y58 = 1'b1;	
							y61 = 1'b1;	y68 = 1'b1;	
							nx_state = s857;
						end
					else if( ~x69 && x46 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y33 = 1'b1;	
							nx_state = s1236;
						end
					else if( ~x69 && ~x46 && x44 && x35 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s997;
						end
					else if( ~x69 && ~x46 && x44 && ~x35 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s998;
						end
					else if( ~x69 && ~x46 && ~x44 && x14 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s691;
						end
					else if( ~x69 && ~x46 && ~x44 && ~x14 && x40 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s691;
						end
					else if( ~x69 && ~x46 && ~x44 && ~x14 && ~x40 && x38 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s691;
						end
					else if( ~x69 && ~x46 && ~x44 && ~x14 && ~x40 && ~x38 && x39 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s691;
						end
					else if( ~x69 && ~x46 && ~x44 && ~x14 && ~x40 && ~x38 && ~x39 )
						nx_state = s783;
					else nx_state = s783;
				s784 : if( x64 && x3 )
						begin
							y3 = 1'b1;	
							nx_state = s710;
						end
					else if( x64 && ~x3 )
						begin
							y31 = 1'b1;	
							nx_state = s1294;
						end
					else if( ~x64 )
						begin
							y39 = 1'b1;	
							nx_state = s1295;
						end
					else nx_state = s784;
				s785 : if( x64 && x3 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x64 && ~x3 )
						begin
							y31 = 1'b1;	
							nx_state = s1243;
						end
					else if( ~x64 )
						begin
							y47 = 1'b1;	y49 = 1'b1;	y58 = 1'b1;	
							y61 = 1'b1;	y70 = 1'b1;	
							nx_state = s1276;
						end
					else nx_state = s785;
				s786 : if( x64 && x3 )
						begin
							y14 = 1'b1;	
							nx_state = s366;
						end
					else if( x64 && ~x3 )
						begin
							y31 = 1'b1;	
							nx_state = s1296;
						end
					else if( ~x64 )
						begin
							y47 = 1'b1;	y49 = 1'b1;	y58 = 1'b1;	
							y61 = 1'b1;	y68 = 1'b1;	
							nx_state = s1297;
						end
					else nx_state = s786;
				s787 : if( x30 && x9 && x10 && x8 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x30 && x9 && x10 && ~x8 )
						begin
							y8 = 1'b1;	
							nx_state = s784;
						end
					else if( x30 && x9 && ~x10 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x30 && x9 && ~x10 && ~x8 )
						begin
							y8 = 1'b1;	
							nx_state = s785;
						end
					else if( x30 && ~x9 && x10 && x8 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( x30 && ~x9 && x10 && ~x8 && x27 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( x30 && ~x9 && x10 && ~x8 && ~x27 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x30 && ~x9 && ~x10 && x8 )
						begin
							y8 = 1'b1;	
							nx_state = s786;
						end
					else if( x30 && ~x9 && ~x10 && ~x8 && x26 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x30 && ~x9 && ~x10 && ~x8 && ~x26 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( ~x30 && x31 && x9 && x10 && x8 )
						begin
							y9 = 1'b1;	
							nx_state = s790;
						end
					else if( ~x30 && x31 && x9 && x10 && ~x8 && x21 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( ~x30 && x31 && x9 && x10 && ~x8 && ~x21 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x30 && x31 && x9 && x10 && ~x8 && ~x21 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x30 && x31 && x9 && x10 && ~x8 && ~x21 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x30 && x31 && x9 && x10 && ~x8 && ~x21 && ~x23 )
						nx_state = s1;
					else if( ~x30 && x31 && x9 && ~x10 && x8 )
						begin
							y3 = 1'b1;	
							nx_state = s789;
						end
					else if( ~x30 && x31 && x9 && ~x10 && ~x8 && x18 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( ~x30 && x31 && x9 && ~x10 && ~x8 && ~x18 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x30 && x31 && x9 && ~x10 && ~x8 && ~x18 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x30 && x31 && x9 && ~x10 && ~x8 && ~x18 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x30 && x31 && x9 && ~x10 && ~x8 && ~x18 && ~x23 )
						nx_state = s1;
					else if( ~x30 && x31 && ~x9 && x8 && x10 && x19 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( ~x30 && x31 && ~x9 && x8 && x10 && ~x19 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x30 && x31 && ~x9 && x8 && x10 && ~x19 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x30 && x31 && ~x9 && x8 && x10 && ~x19 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x30 && x31 && ~x9 && x8 && x10 && ~x19 && ~x23 )
						nx_state = s1;
					else if( ~x30 && x31 && ~x9 && x8 && ~x10 && x20 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( ~x30 && x31 && ~x9 && x8 && ~x10 && ~x20 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x30 && x31 && ~x9 && x8 && ~x10 && ~x20 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x30 && x31 && ~x9 && x8 && ~x10 && ~x20 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x30 && x31 && ~x9 && x8 && ~x10 && ~x20 && ~x23 )
						nx_state = s1;
					else if( ~x30 && x31 && ~x9 && ~x8 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( ~x30 && ~x31 )
						begin
							y9 = 1'b1;	
							nx_state = s790;
						end
					else nx_state = s787;
				s788 : if( x64 )
						begin
							y15 = 1'b1;	
							nx_state = s1115;
						end
					else if( ~x64 && x30 && x31 )
						begin
							y47 = 1'b1;	y50 = 1'b1;	y61 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s1148;
						end
					else if( ~x64 && x30 && ~x31 )
						begin
							y47 = 1'b1;	y52 = 1'b1;	y61 = 1'b1;	
							y70 = 1'b1;	
							nx_state = s1298;
						end
					else if( ~x64 && ~x30 )
						begin
							y47 = 1'b1;	y49 = 1'b1;	y58 = 1'b1;	
							y61 = 1'b1;	y68 = 1'b1;	
							nx_state = s831;
						end
					else nx_state = s788;
				s789 : if( x64 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x64 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x64 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x64 && ~x14 )
						nx_state = s1;
					else if( ~x64 && x30 )
						begin
							y47 = 1'b1;	y56 = 1'b1;	y61 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s1110;
						end
					else if( ~x64 && ~x30 && x31 )
						begin
							y32 = 1'b1;	
							nx_state = s854;
						end
					else if( ~x64 && ~x30 && ~x31 )
						begin
							y47 = 1'b1;	y50 = 1'b1;	y61 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s1148;
						end
					else nx_state = s789;
				s790 : if( x65 )
						begin
							y47 = 1'b1;	y49 = 1'b1;	y58 = 1'b1;	
							y61 = 1'b1;	y68 = 1'b1;	
							nx_state = s857;
						end
					else if( ~x65 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y60 = 1'b1;	
							nx_state = s1299;
						end
					else nx_state = s790;
				s791 : if( x64 && x62 )
						begin
							y1 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1300;
						end
					else if( x64 && ~x62 && x21 )
						begin
							y4 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y93 = 1'b1;	
							nx_state = s1301;
						end
					else if( x64 && ~x62 && ~x21 && x22 )
						begin
							y4 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y78 = 1'b1;	
							nx_state = s1190;
						end
					else if( x64 && ~x62 && ~x21 && ~x22 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y62 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s1189;
						end
					else if( ~x64 && x62 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y37 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s218;
						end
					else if( ~x64 && ~x62 && x31 && x30 )
						begin
							y47 = 1'b1;	y52 = 1'b1;	y61 = 1'b1;	
							y66 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x64 && ~x62 && x31 && ~x30 )
						begin
							y47 = 1'b1;	y52 = 1'b1;	y61 = 1'b1;	
							y68 = 1'b1;	
							nx_state = s1302;
						end
					else if( ~x64 && ~x62 && ~x31 && x30 )
						begin
							y47 = 1'b1;	y52 = 1'b1;	y61 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s353;
						end
					else if( ~x64 && ~x62 && ~x31 && ~x30 )
						begin
							y47 = 1'b1;	y56 = 1'b1;	y61 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s1110;
						end
					else nx_state = s791;
				s792 : if( x21 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x21 && x22 && x17 && x10 && x15 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s334;
						end
					else if( ~x21 && x22 && x17 && x10 && ~x15 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x21 && x22 && x17 && ~x10 )
						begin
							y13 = 1'b1;	y16 = 1'b1;	
							nx_state = s335;
						end
					else if( ~x21 && x22 && ~x17 && x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s336;
						end
					else if( ~x21 && x22 && ~x17 && ~x10 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	
							nx_state = s220;
						end
					else if( ~x21 && ~x22 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s792;
				s793 : if( x21 && x18 )
						begin
							y14 = 1'b1;	y19 = 1'b1;	
							nx_state = s723;
						end
					else if( x21 && ~x18 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s724;
						end
					else if( ~x21 && x22 && x23 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && x22 && x23 && ~x12 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && x23 && ~x12 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && x23 && ~x12 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x12 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s476;
						end
					else if( ~x21 && ~x22 )
						begin
							y14 = 1'b1;	y19 = 1'b1;	
							nx_state = s723;
						end
					else nx_state = s793;
				s794 : if( x21 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && x22 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && x22 && ~x18 && x19 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && x22 && ~x18 && x19 && ~x15 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x21 && x22 && ~x18 && ~x19 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x16 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x16 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && x16 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s793;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && ~x20 )
						begin
							y12 = 1'b1;	
							nx_state = s245;
						end
					else if( ~x21 && ~x22 && ~x23 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && ~x22 && ~x23 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && ~x22 && ~x23 && ~x18 && x19 && x15 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s666;
						end
					else if( ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s664;
						end
					else if( ~x21 && ~x22 && ~x23 && ~x18 && ~x19 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s112;
						end
					else nx_state = s794;
				s795 : if( x21 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x23 && x22 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x23 && x22 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x23 && x22 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x23 && x22 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x23 && ~x22 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x23 && ~x22 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x23 && ~x22 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x23 && ~x22 && ~x9 )
						nx_state = s1;
					else if( ~x21 && ~x23 && x8 && x22 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x23 && x8 && x22 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x23 && x8 && x22 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && ~x23 && x8 && ~x22 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x23 && x8 && ~x22 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x23 && x8 && ~x22 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x23 && ~x8 )
						nx_state = s1;
					else nx_state = s795;
				s796 : if( x21 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s301;
						end
					else if( ~x21 && ~x22 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s301;
						end
					else nx_state = s796;
				s797 : if( x21 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x21 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && x22 && x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s301;
						end
					else if( ~x21 && ~x22 && x23 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s301;
						end
					else if( ~x21 && ~x22 && ~x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x22 && ~x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x22 && ~x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 && ~x8 )
						nx_state = s1;
					else nx_state = s797;
				s798 : if( 1'b1 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s107;
						end
					else nx_state = s798;
				s799 : if( x21 && x18 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && x18 && x15 && ~x17 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	
							nx_state = s807;
						end
					else if( x21 && x18 && ~x15 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x21 && ~x18 && x19 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && ~x18 && x19 && x15 && ~x17 )
						begin
							y8 = 1'b1;	
							nx_state = s568;
						end
					else if( x21 && ~x18 && x19 && ~x15 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s296;
						end
					else if( x21 && ~x18 && ~x19 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x21 && x22 && x23 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && x22 && x23 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && x22 && x23 && ~x18 && x19 && x15 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s666;
						end
					else if( ~x21 && x22 && x23 && ~x18 && x19 && ~x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x21 && x22 && x23 && ~x18 && ~x19 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x21 && x22 && ~x23 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s301;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x16 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x16 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && x16 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s793;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && x18 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x18 && x17 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x18 && ~x17 && x5 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s334;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x18 && ~x17 && ~x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && ~x20 )
						begin
							y12 = 1'b1;	
							nx_state = s245;
						end
					else if( ~x21 && ~x22 && ~x23 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && ~x22 && ~x23 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && ~x22 && ~x23 && ~x18 && x19 && x15 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s666;
						end
					else if( ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x21 && ~x22 && ~x23 && ~x18 && ~x19 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s112;
						end
					else nx_state = s799;
				s800 : if( x69 && x62 && x64 && x17 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							nx_state = s1303;
						end
					else if( x69 && x62 && x64 && ~x17 )
						begin
							y1 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s1144;
						end
					else if( x69 && x62 && ~x64 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s822;
						end
					else if( x69 && x62 && ~x64 && ~x10 && x8 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	
							nx_state = s263;
						end
					else if( x69 && x62 && ~x64 && ~x10 && ~x8 )
						begin
							y4 = 1'b1;	y18 = 1'b1;	
							nx_state = s234;
						end
					else if( x69 && ~x62 )
						begin
							y13 = 1'b1;	
							nx_state = s450;
						end
					else if( ~x69 && x64 && x61 && x37 && x28 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && x64 && x61 && x37 && ~x28 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && x64 && x61 && ~x37 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( ~x69 && x64 && ~x61 && x2 && x10 && x1 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s201;
						end
					else if( ~x69 && x64 && ~x61 && x2 && x10 && x1 && ~x3 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( ~x69 && x64 && ~x61 && x2 && x10 && x1 && ~x3 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x69 && x64 && ~x61 && x2 && x10 && ~x1 && x9 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else if( ~x69 && x64 && ~x61 && x2 && x10 && ~x1 && ~x9 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( ~x69 && x64 && ~x61 && x2 && ~x10 )
						nx_state = s800;
					else if( ~x69 && x64 && ~x61 && ~x2 && x10 && x1 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && x64 && ~x61 && ~x2 && x10 && ~x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x69 && x64 && ~x61 && ~x2 && ~x10 )
						nx_state = s800;
					else if( ~x69 && ~x64 && x14 && x37 && x28 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x69 && ~x64 && x14 && x37 && ~x28 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x69 && ~x64 && x14 && ~x37 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( ~x69 && ~x64 && ~x14 && x2 && x10 && x1 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s201;
						end
					else if( ~x69 && ~x64 && ~x14 && x2 && x10 && x1 && ~x3 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( ~x69 && ~x64 && ~x14 && x2 && x10 && x1 && ~x3 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x69 && ~x64 && ~x14 && x2 && x10 && ~x1 && x9 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else if( ~x69 && ~x64 && ~x14 && x2 && x10 && ~x1 && ~x9 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( ~x69 && ~x64 && ~x14 && x2 && ~x10 )
						nx_state = s800;
					else if( ~x69 && ~x64 && ~x14 && ~x2 && x10 && x1 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x69 && ~x64 && ~x14 && ~x2 && x10 && ~x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x69 && ~x64 && ~x14 && ~x2 && ~x10 )
						nx_state = s800;
					else nx_state = s800;
				s801 : if( x63 && x11 && x43 && x13 && x8 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x63 && x11 && x43 && x13 && ~x8 && x1 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x63 && x11 && x43 && x13 && ~x8 && ~x1 )
						nx_state = s801;
					else if( x63 && x11 && x43 && ~x13 && x10 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( x63 && x11 && x43 && ~x13 && ~x10 && x8 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x63 && x11 && x43 && ~x13 && ~x10 && ~x8 && x1 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x63 && x11 && x43 && ~x13 && ~x10 && ~x8 && ~x1 )
						nx_state = s801;
					else if( x63 && x11 && ~x43 && x8 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x63 && x11 && ~x43 && ~x8 && x1 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x63 && x11 && ~x43 && ~x8 && ~x1 )
						nx_state = s801;
					else if( x63 && ~x11 && x12 && x8 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x63 && ~x11 && x12 && ~x8 && x1 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x63 && ~x11 && x12 && ~x8 && ~x1 )
						nx_state = s801;
					else if( x63 && ~x11 && ~x12 && x44 && x45 && x8 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x63 && ~x11 && ~x12 && x44 && x45 && ~x8 && x1 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x63 && ~x11 && ~x12 && x44 && x45 && ~x8 && ~x1 )
						nx_state = s801;
					else if( x63 && ~x11 && ~x12 && x44 && ~x45 && x41 && x40 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s182;
						end
					else if( x63 && ~x11 && ~x12 && x44 && ~x45 && x41 && ~x40 && x7 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( x63 && ~x11 && ~x12 && x44 && ~x45 && x41 && ~x40 && x7 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( x63 && ~x11 && ~x12 && x44 && ~x45 && x41 && ~x40 && x7 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( x63 && ~x11 && ~x12 && x44 && ~x45 && x41 && ~x40 && x7 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x63 && ~x11 && ~x12 && x44 && ~x45 && x41 && ~x40 && x7 && x15 && ~x47 && ~x1 )
						nx_state = s801;
					else if( x63 && ~x11 && ~x12 && x44 && ~x45 && x41 && ~x40 && x7 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x63 && ~x11 && ~x12 && x44 && ~x45 && x41 && ~x40 && x7 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x63 && ~x11 && ~x12 && x44 && ~x45 && x41 && ~x40 && x7 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x63 && ~x11 && ~x12 && x44 && ~x45 && x41 && ~x40 && ~x7 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s902;
						end
					else if( x63 && ~x11 && ~x12 && x44 && ~x45 && ~x41 && x8 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x63 && ~x11 && ~x12 && x44 && ~x45 && ~x41 && ~x8 && x1 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x63 && ~x11 && ~x12 && x44 && ~x45 && ~x41 && ~x8 && ~x1 )
						nx_state = s801;
					else if( x63 && ~x11 && ~x12 && ~x44 && x8 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x63 && ~x11 && ~x12 && ~x44 && ~x8 && x1 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s454;
						end
					else if( x63 && ~x11 && ~x12 && ~x44 && ~x8 && ~x1 )
						nx_state = s801;
					else if( ~x63 && x9 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( ~x63 && ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s924;
						end
					else nx_state = s801;
				s802 : if( x64 && x40 && x14 && x8 && x10 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x64 && x40 && x14 && x8 && ~x10 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x64 && x40 && x14 && ~x8 && x30 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( x64 && x40 && x14 && ~x8 && x30 && ~x1 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s736;
						end
					else if( x64 && x40 && x14 && ~x8 && x30 && ~x1 && ~x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s915;
						end
					else if( x64 && x40 && x14 && ~x8 && ~x30 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x64 && x40 && ~x14 && x32 && x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( x64 && x40 && ~x14 && x32 && ~x3 )
						nx_state = s802;
					else if( x64 && x40 && ~x14 && ~x32 && x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x64 && x40 && ~x14 && ~x32 && ~x3 )
						nx_state = s802;
					else if( x64 && ~x40 && x16 && x45 && x29 && x42 && x27 )
						begin
							y13 = 1'b1;	
							nx_state = s450;
						end
					else if( x64 && ~x40 && x16 && x45 && x29 && x42 && ~x27 )
						nx_state = s802;
					else if( x64 && ~x40 && x16 && x45 && x29 && ~x42 && x27 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x64 && ~x40 && x16 && x45 && x29 && ~x42 && ~x27 )
						nx_state = s802;
					else if( x64 && ~x40 && x16 && x45 && ~x29 && x33 && x27 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x64 && ~x40 && x16 && x45 && ~x29 && x33 && ~x27 )
						nx_state = s802;
					else if( x64 && ~x40 && x16 && x45 && ~x29 && ~x33 && x43 && x27 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( x64 && ~x40 && x16 && x45 && ~x29 && ~x33 && x43 && ~x27 )
						nx_state = s802;
					else if( x64 && ~x40 && x16 && x45 && ~x29 && ~x33 && ~x43 && x27 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x64 && ~x40 && x16 && x45 && ~x29 && ~x33 && ~x43 && ~x27 )
						nx_state = s802;
					else if( x64 && ~x40 && x16 && ~x45 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x64 && ~x40 && ~x16 && x37 && x44 && x1 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x64 && ~x40 && ~x16 && x37 && x44 && ~x1 )
						nx_state = s802;
					else if( x64 && ~x40 && ~x16 && x37 && ~x44 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x64 && ~x40 && ~x16 && ~x37 && x25 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x64 && ~x40 && ~x16 && ~x37 && ~x25 && x5 && x4 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( x64 && ~x40 && ~x16 && ~x37 && ~x25 && x5 && ~x4 )
						nx_state = s802;
					else if( x64 && ~x40 && ~x16 && ~x37 && ~x25 && ~x5 && x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x64 && ~x40 && ~x16 && ~x37 && ~x25 && ~x5 && ~x4 )
						nx_state = s802;
					else if( ~x64 && x44 && x14 && x8 && x10 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x64 && x44 && x14 && x8 && ~x10 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x64 && x44 && x14 && ~x8 && x30 && x37 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s871;
						end
					else if( ~x64 && x44 && x14 && ~x8 && x30 && ~x37 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s737;
						end
					else if( ~x64 && x44 && x14 && ~x8 && x30 && ~x37 && ~x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s915;
						end
					else if( ~x64 && x44 && x14 && ~x8 && ~x30 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x64 && x44 && ~x14 && x32 && x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( ~x64 && x44 && ~x14 && x32 && ~x3 )
						nx_state = s802;
					else if( ~x64 && x44 && ~x14 && ~x32 && x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x64 && x44 && ~x14 && ~x32 && ~x3 )
						nx_state = s802;
					else if( ~x64 && ~x44 && x16 && x54 && x29 && x48 && x27 )
						begin
							y13 = 1'b1;	
							nx_state = s450;
						end
					else if( ~x64 && ~x44 && x16 && x54 && x29 && x48 && ~x27 )
						nx_state = s802;
					else if( ~x64 && ~x44 && x16 && x54 && x29 && ~x48 && x27 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x64 && ~x44 && x16 && x54 && x29 && ~x48 && ~x27 )
						nx_state = s802;
					else if( ~x64 && ~x44 && x16 && x54 && ~x29 && x33 && x27 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x64 && ~x44 && x16 && x54 && ~x29 && x33 && ~x27 )
						nx_state = s802;
					else if( ~x64 && ~x44 && x16 && x54 && ~x29 && ~x33 && x49 && x27 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s870;
						end
					else if( ~x64 && ~x44 && x16 && x54 && ~x29 && ~x33 && x49 && ~x27 )
						nx_state = s802;
					else if( ~x64 && ~x44 && x16 && x54 && ~x29 && ~x33 && ~x49 && x27 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x64 && ~x44 && x16 && x54 && ~x29 && ~x33 && ~x49 && ~x27 )
						nx_state = s802;
					else if( ~x64 && ~x44 && x16 && ~x54 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x64 && ~x44 && ~x16 && x37 && x55 && x1 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x64 && ~x44 && ~x16 && x37 && x55 && ~x1 )
						nx_state = s802;
					else if( ~x64 && ~x44 && ~x16 && x37 && ~x55 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x64 && ~x44 && ~x16 && ~x37 && x25 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x64 && ~x44 && ~x16 && ~x37 && ~x25 && x5 && x4 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( ~x64 && ~x44 && ~x16 && ~x37 && ~x25 && x5 && ~x4 )
						nx_state = s802;
					else if( ~x64 && ~x44 && ~x16 && ~x37 && ~x25 && ~x5 && x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x64 && ~x44 && ~x16 && ~x37 && ~x25 && ~x5 && ~x4 )
						nx_state = s802;
					else nx_state = s802;
				s803 : if( x62 && x61 && x19 && x13 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x62 && x61 && x19 && ~x13 && x32 && x18 && x12 )
						nx_state = s803;
					else if( x62 && x61 && x19 && ~x13 && x32 && x18 && ~x12 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s875;
						end
					else if( x62 && x61 && x19 && ~x13 && x32 && ~x18 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( x62 && x61 && x19 && ~x13 && ~x32 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s840;
						end
					else if( x62 && x61 && ~x19 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( x62 && ~x61 && x17 && x19 && x10 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( x62 && ~x61 && x17 && x19 && ~x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s875;
						end
					else if( x62 && ~x61 && x17 && ~x19 )
						nx_state = s803;
					else if( x62 && ~x61 && ~x17 && x20 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s1097;
						end
					else if( x62 && ~x61 && ~x17 && ~x20 && x2 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( x62 && ~x61 && ~x17 && ~x20 && ~x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x62 && x63 && x55 && x19 && x44 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s443;
						end
					else if( ~x62 && x63 && x55 && x19 && ~x44 && x32 && x18 && x12 )
						nx_state = s803;
					else if( ~x62 && x63 && x55 && x19 && ~x44 && x32 && x18 && ~x12 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s914;
						end
					else if( ~x62 && x63 && x55 && x19 && ~x44 && x32 && ~x18 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( ~x62 && x63 && x55 && x19 && ~x44 && ~x32 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x62 && x63 && x55 && ~x19 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( ~x62 && x63 && ~x55 && x17 && x50 && x10 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s734;
						end
					else if( ~x62 && x63 && ~x55 && x17 && x50 && ~x10 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s914;
						end
					else if( ~x62 && x63 && ~x55 && x17 && ~x50 )
						nx_state = s803;
					else if( ~x62 && x63 && ~x55 && ~x17 && x51 )
						begin
							y11 = 1'b1;	
							nx_state = s250;
						end
					else if( ~x62 && x63 && ~x55 && ~x17 && ~x51 && x33 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x62 && x63 && ~x55 && ~x17 && ~x51 && ~x33 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x62 && ~x63 && x40 && x19 && x13 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s443;
						end
					else if( ~x62 && ~x63 && x40 && x19 && ~x13 && x32 && x18 && x12 )
						nx_state = s803;
					else if( ~x62 && ~x63 && x40 && x19 && ~x13 && x32 && x18 && ~x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s915;
						end
					else if( ~x62 && ~x63 && x40 && x19 && ~x13 && x32 && ~x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( ~x62 && ~x63 && x40 && x19 && ~x13 && ~x32 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x62 && ~x63 && x40 && ~x19 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x62 && ~x63 && ~x40 && x17 && x19 && x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s736;
						end
					else if( ~x62 && ~x63 && ~x40 && x17 && x19 && ~x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s915;
						end
					else if( ~x62 && ~x63 && ~x40 && x17 && ~x19 )
						nx_state = s803;
					else if( ~x62 && ~x63 && ~x40 && ~x17 && x20 )
						begin
							y11 = 1'b1;	
							nx_state = s250;
						end
					else if( ~x62 && ~x63 && ~x40 && ~x17 && ~x20 && x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x62 && ~x63 && ~x40 && ~x17 && ~x20 && ~x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else nx_state = s803;
				s804 : if( x15 && x64 && x1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1000;
						end
					else if( x15 && x64 && ~x1 )
						begin
							y11 = 1'b1;	
							nx_state = s248;
						end
					else if( x15 && ~x64 && x37 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1000;
						end
					else if( x15 && ~x64 && ~x37 )
						begin
							y11 = 1'b1;	
							nx_state = s248;
						end
					else if( ~x15 )
						begin
							y11 = 1'b1;	
							nx_state = s248;
						end
					else nx_state = s804;
				s805 : if( x21 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x21 && x22 && x23 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && x6 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && x22 && ~x23 && x6 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && x22 && ~x23 && x6 && ~x18 && x19 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && x22 && ~x23 && x6 && ~x18 && x19 && ~x15 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x21 && x22 && ~x23 && x6 && ~x18 && ~x19 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s465;
						end
					else if( ~x21 && x22 && ~x23 && ~x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s107;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x20 && x16 && x18 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x20 && x16 && ~x18 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x20 && ~x16 && x17 && x18 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s296;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x20 && ~x16 && x17 && ~x18 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y20 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s795;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x20 && ~x16 && ~x17 && x18 && x11 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s666;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x20 && ~x16 && ~x17 && x18 && ~x11 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x20 && ~x16 && ~x17 && x18 && ~x11 && x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && x19 && x20 && ~x16 && ~x17 && x18 && ~x11 && ~x9 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && x19 && x20 && ~x16 && ~x17 && ~x18 && x10 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s666;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x20 && ~x16 && ~x17 && ~x18 && ~x10 && x9 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x20 && ~x16 && ~x17 && ~x18 && ~x10 && x9 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && x19 && x20 && ~x16 && ~x17 && ~x18 && ~x10 && ~x9 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && x19 && ~x20 && x17 && x16 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x20 && x17 && ~x16 && x18 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x20 && x17 && ~x16 && ~x18 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s796;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x20 && ~x17 && x18 && x16 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x20 && ~x17 && x18 && ~x16 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s797;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x20 && ~x17 && ~x18 && x3 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x20 && ~x17 && ~x18 && ~x3 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x20 && ~x17 && ~x18 && ~x3 && ~x5 && x16 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s795;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x20 && ~x17 && ~x18 && ~x3 && ~x5 && ~x16 )
						begin
							y16 = 1'b1;	y20 = 1'b1;	
							nx_state = s795;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && x16 && x3 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && x16 && ~x3 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && x16 && ~x3 && ~x5 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && x17 && x18 && x3 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && x17 && x18 && ~x3 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && x17 && x18 && ~x3 && ~x5 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s795;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && x17 && ~x18 && x15 && x3 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && x17 && ~x18 && x15 && ~x3 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && x17 && ~x18 && x15 && ~x3 && ~x5 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s795;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && x17 && ~x18 && ~x15 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x17 && x18 && x13 && x3 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x17 && x18 && x13 && ~x3 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x17 && x18 && x13 && ~x3 && ~x5 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s795;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x17 && x18 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x17 && ~x18 && x12 && x3 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x17 && ~x18 && x12 && ~x3 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x17 && ~x18 && ~x12 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x17 && ~x18 && ~x12 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x17 && ~x18 && ~x12 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x17 && ~x18 && ~x12 && ~x9 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x19 && ~x20 && x3 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && ~x20 && ~x3 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s799;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && ~x20 && ~x3 && ~x5 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( ~x21 && ~x22 && ~x23 )
						nx_state = s1;
					else nx_state = s805;
				s806 : if( 1'b1 )
						begin
							y7 = 1'b1;	
							nx_state = s747;
						end
					else nx_state = s806;
				s807 : if( x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s643;
						end
					else if( x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x8 )
						nx_state = s1;
					else nx_state = s807;
				s808 : if( 1'b1 )
						begin
							y3 = 1'b1;	y12 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s1304;
						end
					else nx_state = s808;
				s809 : if( x22 && x21 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( x22 && ~x21 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1305;
						end
					else if( ~x22 && x19 && x21 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( ~x22 && x19 && ~x21 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1305;
						end
					else if( ~x22 && ~x19 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else nx_state = s809;
				s810 : if( x21 && x18 && x16 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( x21 && x18 && ~x16 && x13 && x15 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( x21 && x18 && ~x16 && x13 && ~x15 && x17 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1305;
						end
					else if( x21 && x18 && ~x16 && x13 && ~x15 && ~x17 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( x21 && x18 && ~x16 && ~x13 && x17 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1305;
						end
					else if( x21 && x18 && ~x16 && ~x13 && ~x17 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( x21 && ~x18 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1305;
						end
					else if( ~x21 && x19 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( ~x21 && ~x19 && x22 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( ~x21 && ~x19 && ~x22 && x20 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1305;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x20 && x16 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && x15 && x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && x15 && ~x13 && x17 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1305;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && x15 && ~x13 && ~x17 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && ~x15 && x17 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1305;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && ~x15 && ~x17 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else nx_state = s810;
				s811 : if( x60 && x61 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s554;
						end
					else if( x60 && ~x61 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x60 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else nx_state = s811;
				s812 : if( x60 && x61 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s555;
						end
					else if( x60 && ~x61 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x60 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else nx_state = s812;
				s813 : if( x20 && x17 && x15 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s556;
						end
					else if( x20 && x17 && ~x15 && x16 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s131;
						end
					else if( x20 && x17 && ~x15 && ~x16 )
						begin
							y7 = 1'b1;	y12 = 1'b1;	
							nx_state = s610;
						end
					else if( x20 && ~x17 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	y22 = 1'b1;	
							nx_state = s1070;
						end
					else if( ~x20 && x21 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	y22 = 1'b1;	
							nx_state = s1070;
						end
					else if( ~x20 && ~x21 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s369;
						end
					else nx_state = s813;
				s814 : if( 1'b1 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else nx_state = s814;
				s815 : if( 1'b1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s328;
						end
					else nx_state = s815;
				s816 : if( x70 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s216;
						end
					else if( ~x70 && x7 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s216;
						end
					else if( ~x70 && ~x7 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s96;
						end
					else nx_state = s816;
				s817 : if( x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s216;
						end
					else if( ~x15 && x13 && x11 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s767;
						end
					else if( ~x15 && x13 && ~x11 && x6 && x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s1284;
						end
					else if( ~x15 && x13 && ~x11 && x6 && ~x4 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s761;
						end
					else if( ~x15 && x13 && ~x11 && ~x6 && x5 )
						begin
							y2 = 1'b1;	
							nx_state = s768;
						end
					else if( ~x15 && x13 && ~x11 && ~x6 && ~x5 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s1280;
						end
					else if( ~x15 && ~x13 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s766;
						end
					else if( ~x15 && ~x13 && ~x14 && x9 )
						begin
							y10 = 1'b1;	
							nx_state = s766;
						end
					else if( ~x15 && ~x13 && ~x14 && ~x9 && x6 && x2 )
						begin
							y10 = 1'b1;	
							nx_state = s766;
						end
					else if( ~x15 && ~x13 && ~x14 && ~x9 && x6 && ~x2 )
						nx_state = s817;
					else if( ~x15 && ~x13 && ~x14 && ~x9 && ~x6 && x8 )
						begin
							y10 = 1'b1;	
							nx_state = s766;
						end
					else if( ~x15 && ~x13 && ~x14 && ~x9 && ~x6 && ~x8 )
						nx_state = s817;
					else nx_state = s817;
				s818 : if( x69 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s1182;
						end
					else if( ~x69 && x10 && x6 && x7 && x33 && x3 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( ~x69 && x10 && x6 && x7 && x33 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x69 && x10 && x6 && x7 && x33 && ~x3 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x69 && x10 && x6 && x7 && ~x33 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( ~x69 && x10 && x6 && ~x7 && x39 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s818;
						end
					else if( ~x69 && x10 && x6 && ~x7 && ~x39 && x33 && x3 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( ~x69 && x10 && x6 && ~x7 && ~x39 && x33 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x69 && x10 && x6 && ~x7 && ~x39 && x33 && ~x3 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x69 && x10 && x6 && ~x7 && ~x39 && ~x33 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( ~x69 && x10 && ~x6 && x2 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s818;
						end
					else if( ~x69 && x10 && ~x6 && ~x2 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x69 && ~x10 && x11 && x5 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s818;
						end
					else if( ~x69 && ~x10 && x11 && ~x5 && x37 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( ~x69 && ~x10 && x11 && ~x5 && ~x37 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && ~x10 && ~x11 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else nx_state = s818;
				s819 : if( 1'b1 )
						begin
							y8 = 1'b1;	y17 = 1'b1;	y23 = 1'b1;	
							nx_state = s303;
						end
					else nx_state = s819;
				s820 : if( x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x11 )
						nx_state = s1;
					else nx_state = s820;
				s821 : if( x19 && x18 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( x19 && ~x18 )
						begin
							y2 = 1'b1;	
							nx_state = s1306;
						end
					else if( ~x19 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else nx_state = s821;
				s822 : if( x70 && x62 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s822;
						end
					else if( x70 && x62 && x9 && ~x10 && x8 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	
							nx_state = s263;
						end
					else if( x70 && x62 && x9 && ~x10 && ~x8 )
						begin
							y4 = 1'b1;	y18 = 1'b1;	
							nx_state = s234;
						end
					else if( x70 && x62 && ~x9 )
						begin
							y13 = 1'b1;	
							nx_state = s800;
						end
					else if( x70 && ~x62 && x65 )
						begin
							y69 = 1'b1;	
							nx_state = s1123;
						end
					else if( x70 && ~x62 && ~x65 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s328;
						end
					else if( ~x70 && x65 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s167;
						end
					else if( ~x70 && ~x65 && x63 && x1 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s294;
						end
					else if( ~x70 && ~x65 && x63 && ~x1 && x18 && x15 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( ~x70 && ~x65 && x63 && ~x1 && x18 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x70 && ~x65 && x63 && ~x1 && x18 && ~x15 && x16 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x70 && ~x65 && x63 && ~x1 && x18 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s299;
						end
					else if( ~x70 && ~x65 && x63 && ~x1 && ~x18 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s295;
						end
					else if( ~x70 && ~x65 && ~x63 )
						begin
							y3 = 1'b1;	y22 = 1'b1;	y37 = 1'b1;	
							nx_state = s1035;
						end
					else nx_state = s822;
				s823 : if( x62 )
						begin
							y5 = 1'b1;	
							nx_state = s937;
						end
					else if( ~x62 )
						begin
							y7 = 1'b1;	y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s1307;
						end
					else nx_state = s823;
				s824 : if( 1'b1 )
						begin
							y13 = 1'b1;	y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s824;
				s825 : if( x21 && x20 && x18 && x15 && x10 && x11 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s600;
						end
					else if( x21 && x20 && x18 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s601;
						end
					else if( x21 && x20 && x18 && x15 && x10 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s776;
						end
					else if( x21 && x20 && x18 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( x21 && x20 && x18 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s602;
						end
					else if( x21 && x20 && x18 && ~x15 && x16 && x10 && x12 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( x21 && x20 && x18 && ~x15 && x16 && x10 && ~x12 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x21 && x20 && x18 && ~x15 && x16 && ~x10 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( x21 && x20 && x18 && ~x15 && ~x16 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s421;
						end
					else if( x21 && x20 && ~x18 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	
							nx_state = s826;
						end
					else if( x21 && ~x20 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s603;
						end
					else if( ~x21 && x18 && x15 && x10 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x21 && x18 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s605;
						end
					else if( ~x21 && x18 && x15 && x10 && ~x11 && ~x12 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s606;
						end
					else if( ~x21 && x18 && x15 && ~x10 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s359;
						end
					else if( ~x21 && x18 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s600;
						end
					else if( ~x21 && x18 && ~x15 && x16 && x10 && x12 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( ~x21 && x18 && ~x15 && x16 && x10 && ~x12 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( ~x21 && x18 && ~x15 && x16 && ~x10 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s563;
						end
					else if( ~x21 && x18 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s607;
						end
					else if( ~x21 && ~x18 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s129;
						end
					else nx_state = s825;
				s826 : if( x21 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s625;
						end
					else if( ~x21 )
						nx_state = s1;
					else nx_state = s826;
				s827 : if( 1'b1 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s149;
						end
					else nx_state = s827;
				s828 : if( x22 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x22 )
						begin
							y17 = 1'b1;	
							nx_state = s98;
						end
					else nx_state = s828;
				s829 : if( x21 && x16 && x15 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s181;
						end
					else if( x21 && x16 && x15 && ~x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s441;
						end
					else if( x21 && x16 && ~x15 && x10 )
						begin
							y18 = 1'b1;	
							nx_state = s63;
						end
					else if( x21 && x16 && ~x15 && ~x10 )
						begin
							y14 = 1'b1;	y16 = 1'b1;	
							nx_state = s492;
						end
					else if( x21 && ~x16 && x17 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s679;
						end
					else if( x21 && ~x16 && ~x17 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s680;
						end
					else if( x21 && ~x16 && ~x17 && ~x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s443;
						end
					else if( ~x21 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else nx_state = s829;
				s830 : if( 1'b1 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s559;
						end
					else nx_state = s830;
				s831 : if( 1'b1 )
						begin
							y47 = 1'b1;	y53 = 1'b1;	y61 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s1308;
						end
					else nx_state = s831;
				s832 : if( 1'b1 )
						begin
							y8 = 1'b1;	y22 = 1'b1;	
							nx_state = s570;
						end
					else nx_state = s832;
				s833 : if( x55 && x37 && x28 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s503;
						end
					else if( x55 && x37 && ~x28 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( x55 && ~x37 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x55 && x33 && x32 && x10 && x3 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( ~x55 && x33 && x32 && x10 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x55 && x33 && x32 && x10 && ~x3 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x55 && x33 && x32 && ~x10 )
						nx_state = s833;
					else if( ~x55 && x33 && ~x32 && x10 && x9 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s1125;
						end
					else if( ~x55 && x33 && ~x32 && x10 && ~x9 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x55 && x33 && ~x32 && ~x10 )
						nx_state = s833;
					else if( ~x55 && ~x33 && x32 && x10 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( ~x55 && ~x33 && x32 && ~x10 )
						nx_state = s833;
					else if( ~x55 && ~x33 && ~x32 && x10 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s498;
						end
					else if( ~x55 && ~x33 && ~x32 && ~x10 )
						nx_state = s833;
					else nx_state = s833;
				s834 : if( 1'b1 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else nx_state = s834;
				s835 : if( x70 && x64 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x70 && x64 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x70 && x64 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x70 && x64 && ~x14 )
						nx_state = s1;
					else if( x70 && ~x64 && x31 && x30 )
						begin
							y47 = 1'b1;	y52 = 1'b1;	y61 = 1'b1;	
							y66 = 1'b1;	
							nx_state = s54;
						end
					else if( x70 && ~x64 && x31 && ~x30 )
						begin
							y47 = 1'b1;	y52 = 1'b1;	y61 = 1'b1;	
							y68 = 1'b1;	
							nx_state = s1302;
						end
					else if( x70 && ~x64 && ~x31 && x30 )
						begin
							y47 = 1'b1;	y52 = 1'b1;	y61 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s353;
						end
					else if( x70 && ~x64 && ~x31 && ~x30 )
						begin
							y47 = 1'b1;	y56 = 1'b1;	y61 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s1110;
						end
					else if( ~x70 && x65 )
						nx_state = s47;
					else if( ~x70 && ~x65 && x66 && x23 && x18 && x15 && x7 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s151;
						end
					else if( ~x70 && ~x65 && x66 && x23 && x18 && x15 && ~x7 && x9 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && ~x65 && x66 && x23 && x18 && x15 && ~x7 && ~x9 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x70 && ~x65 && x66 && x23 && x18 && ~x15 && x7 && x9 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s274;
						end
					else if( ~x70 && ~x65 && x66 && x23 && x18 && ~x15 && x7 && ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x70 && ~x65 && x66 && x23 && x18 && ~x15 && ~x7 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s274;
						end
					else if( ~x70 && ~x65 && x66 && x23 && ~x18 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x70 && ~x65 && x66 && ~x23 && x9 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x65 && x66 && ~x23 && ~x9 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( ~x70 && ~x65 && x66 && ~x23 && ~x9 && ~x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x70 && ~x65 && ~x66 )
						begin
							y5 = 1'b1;	
							nx_state = s66;
						end
					else nx_state = s835;
				s836 : if( 1'b1 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y8 = 1'b1;	y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s1309;
						end
					else nx_state = s836;
				s837 : if( x61 && x16 && x17 && x11 && x13 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s251;
						end
					else if( x61 && x16 && x17 && x11 && ~x13 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s564;
						end
					else if( x61 && x16 && x17 && ~x11 && x12 && x13 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s565;
						end
					else if( x61 && x16 && x17 && ~x11 && x12 && ~x13 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s242;
						end
					else if( x61 && x16 && x17 && ~x11 && ~x12 && x13 && x15 )
						begin
							y15 = 1'b1;	
							nx_state = s243;
						end
					else if( x61 && x16 && x17 && ~x11 && ~x12 && x13 && ~x15 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x61 && x16 && x17 && ~x11 && ~x12 && x13 && ~x15 && x18 && ~x14 )
						nx_state = s1;
					else if( x61 && x16 && x17 && ~x11 && ~x12 && x13 && ~x15 && ~x18 )
						nx_state = s1;
					else if( x61 && x16 && x17 && ~x11 && ~x12 && ~x13 && x14 )
						begin
							y15 = 1'b1;	
							nx_state = s243;
						end
					else if( x61 && x16 && x17 && ~x11 && ~x12 && ~x13 && ~x14 && x18 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x61 && x16 && x17 && ~x11 && ~x12 && ~x13 && ~x14 && x18 && ~x15 )
						nx_state = s1;
					else if( x61 && x16 && x17 && ~x11 && ~x12 && ~x13 && ~x14 && ~x18 )
						nx_state = s1;
					else if( x61 && x16 && ~x17 && x12 && x11 && x13 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x61 && x16 && ~x17 && x12 && x11 && x13 && ~x3 && x2 )
						nx_state = s47;
					else if( x61 && x16 && ~x17 && x12 && x11 && x13 && ~x3 && ~x2 )
						begin
							y22 = 1'b1;	
							nx_state = s683;
						end
					else if( x61 && x16 && ~x17 && x12 && x11 && ~x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else if( x61 && x16 && ~x17 && x12 && ~x11 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else if( x61 && x16 && ~x17 && x12 && ~x11 && ~x13 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s566;
						end
					else if( x61 && x16 && ~x17 && ~x12 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x61 && x16 && ~x17 && ~x12 && ~x3 && x2 )
						nx_state = s47;
					else if( x61 && x16 && ~x17 && ~x12 && ~x3 && ~x2 && x13 && x11 )
						begin
							y22 = 1'b1;	
							nx_state = s130;
						end
					else if( x61 && x16 && ~x17 && ~x12 && ~x3 && ~x2 && x13 && ~x11 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x61 && x16 && ~x17 && ~x12 && ~x3 && ~x2 && ~x13 && x11 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y24 = 1'b1;	
							nx_state = s136;
						end
					else if( x61 && x16 && ~x17 && ~x12 && ~x3 && ~x2 && ~x13 && ~x11 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x61 && ~x16 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( x61 && ~x16 && ~x3 && x17 && x13 && x11 && x9 && x2 )
						nx_state = s47;
					else if( x61 && ~x16 && ~x3 && x17 && x13 && x11 && x9 && ~x2 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s707;
						end
					else if( x61 && ~x16 && ~x3 && x17 && x13 && x11 && ~x9 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x61 && ~x16 && ~x3 && x17 && x13 && x11 && ~x9 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x61 && ~x16 && ~x3 && x17 && x13 && x11 && ~x9 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x61 && ~x16 && ~x3 && x17 && x13 && x11 && ~x9 && ~x18 )
						nx_state = s1;
					else if( x61 && ~x16 && ~x3 && x17 && x13 && ~x11 && x12 && x2 )
						nx_state = s47;
					else if( x61 && ~x16 && ~x3 && x17 && x13 && ~x11 && x12 && ~x2 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s707;
						end
					else if( x61 && ~x16 && ~x3 && x17 && x13 && ~x11 && ~x12 && x8 && x2 )
						nx_state = s47;
					else if( x61 && ~x16 && ~x3 && x17 && x13 && ~x11 && ~x12 && x8 && ~x2 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s707;
						end
					else if( x61 && ~x16 && ~x3 && x17 && x13 && ~x11 && ~x12 && ~x8 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x61 && ~x16 && ~x3 && x17 && x13 && ~x11 && ~x12 && ~x8 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x61 && ~x16 && ~x3 && x17 && x13 && ~x11 && ~x12 && ~x8 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x61 && ~x16 && ~x3 && x17 && x13 && ~x11 && ~x12 && ~x8 && ~x18 )
						nx_state = s1;
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && x11 )
						nx_state = s47;
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && x12 && x10 && x2 )
						nx_state = s47;
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && x12 && x10 && ~x2 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s707;
						end
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && x12 && ~x10 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && x12 && ~x10 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && x12 && ~x10 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && x12 && ~x10 && ~x18 )
						nx_state = s1;
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && x7 && x2 )
						nx_state = s47;
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && x7 && ~x2 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s707;
						end
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && ~x7 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && ~x7 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && ~x7 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && ~x7 && ~x18 )
						nx_state = s1;
					else if( x61 && ~x16 && ~x3 && ~x17 && x2 )
						nx_state = s47;
					else if( x61 && ~x16 && ~x3 && ~x17 && ~x2 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x61 && x62 && x2 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s564;
						end
					else if( ~x61 && x62 && ~x2 && x19 && x15 && x12 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s491;
						end
					else if( ~x61 && x62 && ~x2 && x19 && x15 && x12 && ~x7 )
						begin
							y12 = 1'b1;	
							nx_state = s490;
						end
					else if( ~x61 && x62 && ~x2 && x19 && x15 && ~x12 && x7 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x61 && x62 && ~x2 && x19 && x15 && ~x12 && ~x7 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s566;
						end
					else if( ~x61 && x62 && ~x2 && x19 && ~x15 && x16 && x7 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s490;
						end
					else if( ~x61 && x62 && ~x2 && x19 && ~x15 && x16 && x7 && ~x12 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s565;
						end
					else if( ~x61 && x62 && ~x2 && x19 && ~x15 && x16 && ~x7 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s487;
						end
					else if( ~x61 && x62 && ~x2 && x19 && ~x15 && ~x16 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x61 && x62 && ~x2 && x19 && ~x15 && ~x16 && ~x7 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x61 && x62 && ~x2 && ~x19 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y23 = 1'b1;	
							nx_state = s993;
						end
					else if( ~x61 && ~x62 )
						nx_state = s1;
					else nx_state = s837;
				s838 : if( x70 && x63 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y22 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s1310;
						end
					else if( x70 && ~x63 )
						begin
							y37 = 1'b1;	
							nx_state = s888;
						end
					else if( ~x70 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s1311;
						end
					else nx_state = s838;
				s839 : if( 1'b1 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else nx_state = s839;
				s840 : if( x61 && x24 && x26 && x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( x61 && x24 && x26 && ~x7 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s280;
						end
					else if( x61 && x24 && ~x26 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s875;
						end
					else if( x61 && ~x24 && x28 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s215;
						end
					else if( x61 && ~x24 && ~x28 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( ~x61 && x31 && x19 && x10 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x61 && x31 && x19 && ~x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s875;
						end
					else if( ~x61 && x31 && ~x19 )
						nx_state = s840;
					else if( ~x61 && ~x31 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s875;
						end
					else nx_state = s840;
				s841 : if( x69 && x63 && x22 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	y38 = 1'b1;	
							nx_state = s1312;
						end
					else if( x69 && x63 && ~x22 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	y26 = 1'b1;	
							nx_state = s1313;
						end
					else if( x69 && ~x63 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s328;
						end
					else if( ~x69 && x61 && x22 && x2 && x33 )
						begin
							y10 = 1'b1;	
							nx_state = s841;
						end
					else if( ~x69 && x61 && x22 && x2 && ~x33 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( ~x69 && x61 && x22 && x2 && ~x33 && ~x13 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s840;
						end
					else if( ~x69 && x61 && x22 && ~x2 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( ~x69 && x61 && ~x22 && x31 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( ~x69 && x61 && ~x22 && ~x31 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( ~x69 && ~x61 && x46 && x3 && x23 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s874;
						end
					else if( ~x69 && ~x61 && x46 && x3 && ~x23 )
						nx_state = s841;
					else if( ~x69 && ~x61 && x46 && ~x3 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( ~x69 && ~x61 && ~x46 && x2 && x23 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s874;
						end
					else if( ~x69 && ~x61 && ~x46 && x2 && ~x23 )
						nx_state = s841;
					else if( ~x69 && ~x61 && ~x46 && ~x2 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else nx_state = s841;
				s842 : if( x9 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s733;
						end
					else if( ~x9 && x37 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s733;
						end
					else if( ~x9 && ~x37 )
						begin
							y10 = 1'b1;	
							nx_state = s841;
						end
					else nx_state = s842;
				s843 : if( x61 && x30 && x16 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( x61 && x30 && x16 && ~x6 && x8 && x19 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s320;
						end
					else if( x61 && x30 && x16 && ~x6 && x8 && ~x19 && x26 && x5 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( x61 && x30 && x16 && ~x6 && x8 && ~x19 && x26 && ~x5 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s733;
						end
					else if( x61 && x30 && x16 && ~x6 && x8 && ~x19 && ~x26 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s738;
						end
					else if( x61 && x30 && x16 && ~x6 && ~x8 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( x61 && x30 && ~x16 && x10 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s840;
						end
					else if( x61 && x30 && ~x16 && ~x10 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( x61 && ~x30 && x5 && x9 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( x61 && ~x30 && x5 && ~x9 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( x61 && ~x30 && ~x5 && x11 && x3 )
						nx_state = s843;
					else if( x61 && ~x30 && ~x5 && x11 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( x61 && ~x30 && ~x5 && ~x11 && x3 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( x61 && ~x30 && ~x5 && ~x11 && ~x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x61 && x51 && x24 && x5 && x36 )
						nx_state = s843;
					else if( ~x61 && x51 && x24 && x5 && ~x36 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x61 && x51 && x24 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( ~x61 && x51 && ~x24 && x31 && x29 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x61 && x51 && ~x24 && x31 && ~x29 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( ~x61 && x51 && ~x24 && ~x31 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x61 && ~x51 && x11 && x35 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x61 && ~x51 && x11 && x35 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( ~x61 && ~x51 && x11 && ~x35 && x60 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( ~x61 && ~x51 && x11 && ~x35 && ~x60 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( ~x61 && ~x51 && ~x11 && x52 && x35 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x61 && ~x51 && ~x11 && x52 && ~x35 && x60 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( ~x61 && ~x51 && ~x11 && x52 && ~x35 && ~x60 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( ~x61 && ~x51 && ~x11 && ~x52 && x3 && x6 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s215;
						end
					else if( ~x61 && ~x51 && ~x11 && ~x52 && x3 && ~x6 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( ~x61 && ~x51 && ~x11 && ~x52 && ~x3 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else nx_state = s843;
				s844 : if( x21 && x10 )
						begin
							y62 = 1'b1;	y65 = 1'b1;	y78 = 1'b1;	
							y90 = 1'b1;	
							nx_state = s1132;
						end
					else if( x21 && ~x10 && x14 && x11 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1130;
						end
					else if( x21 && ~x10 && x14 && ~x11 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1133;
						end
					else if( x21 && ~x10 && ~x14 && x11 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1134;
						end
					else if( x21 && ~x10 && ~x14 && ~x11 )
						begin
							y3 = 1'b1;	y74 = 1'b1;	
							nx_state = s1135;
						end
					else if( ~x21 && x22 && x10 && x11 && x14 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1134;
						end
					else if( ~x21 && x22 && x10 && x11 && ~x14 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1131;
						end
					else if( ~x21 && x22 && x10 && ~x11 && x14 && x19 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x21 && x22 && x10 && ~x11 && x14 && ~x19 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && x10 && ~x11 && x14 && ~x19 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && x10 && ~x11 && x14 && ~x19 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && x10 && ~x11 && x14 && ~x19 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && x10 && ~x11 && ~x14 && x18 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x21 && x22 && x10 && ~x11 && ~x14 && ~x18 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && x10 && ~x11 && ~x14 && ~x18 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && x10 && ~x11 && ~x14 && ~x18 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && x10 && ~x11 && ~x14 && ~x18 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x10 && x14 && x11 && x17 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x21 && x22 && ~x10 && x14 && x11 && ~x17 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && ~x10 && x14 && x11 && ~x17 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && ~x10 && x14 && x11 && ~x17 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x10 && x14 && x11 && ~x17 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x10 && x14 && ~x11 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x21 && x22 && ~x10 && ~x14 && x11 && x16 && x18 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x21 && x22 && ~x10 && ~x14 && x11 && x16 && ~x18 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && ~x10 && ~x14 && x11 && x16 && ~x18 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && ~x10 && ~x14 && x11 && x16 && ~x18 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x10 && ~x14 && x11 && x16 && ~x18 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x10 && ~x14 && x11 && ~x16 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && ~x10 && ~x14 && x11 && ~x16 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && ~x10 && ~x14 && x11 && ~x16 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x10 && ~x14 && x11 && ~x16 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x10 && ~x14 && ~x11 )
						begin
							y102 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x21 && ~x22 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1134;
						end
					else nx_state = s844;
				s845 : if( x62 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x62 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x62 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( x62 && ~x27 )
						nx_state = s1;
					else if( ~x62 && x63 && x67 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x62 && x63 && x67 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x62 && x63 && x67 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( ~x62 && x63 && x67 && ~x22 )
						nx_state = s1;
					else if( ~x62 && x63 && ~x67 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x62 && x63 && ~x67 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x62 && x63 && ~x67 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x62 && x63 && ~x67 && ~x11 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && ~x63 && x64 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && ~x63 && x64 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x64 && ~x6 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 && x65 && x31 )
						begin
							y25 = 1'b1;	
							nx_state = s238;
						end
					else if( ~x62 && ~x63 && ~x64 && x65 && ~x31 )
						begin
							y40 = 1'b1;	
							nx_state = s947;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x66 && x19 && x6 && x5 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x66 && x19 && x6 && ~x5 )
						begin
							y69 = 1'b1;	
							nx_state = s1123;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x66 && x19 && ~x6 && x8 && x9 && x5 )
						begin
							y51 = 1'b1;	
							nx_state = s391;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x66 && x19 && ~x6 && x8 && x9 && ~x5 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y62 = 1'b1;	
							y63 = 1'b1;	y65 = 1'b1;	y66 = 1'b1;	
							nx_state = s1314;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x66 && x19 && ~x6 && x8 && x9 && ~x5 && ~x7 )
						begin
							y5 = 1'b1;	y27 = 1'b1;	y57 = 1'b1;	
							y58 = 1'b1;	
							nx_state = s1314;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x66 && x19 && ~x6 && x8 && ~x9 && x5 )
						begin
							y3 = 1'b1;	y19 = 1'b1;	y53 = 1'b1;	
							nx_state = s1314;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x66 && x19 && ~x6 && x8 && ~x9 && ~x5 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y59 = 1'b1;	
							y60 = 1'b1;	y67 = 1'b1;	y68 = 1'b1;	
							nx_state = s1314;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x66 && x19 && ~x6 && x8 && ~x9 && ~x5 && ~x7 )
						begin
							y5 = 1'b1;	y27 = 1'b1;	y55 = 1'b1;	
							y56 = 1'b1;	
							nx_state = s1314;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x66 && x19 && ~x6 && ~x8 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1314;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x66 && x19 && ~x6 && ~x8 && ~x5 && x7 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y62 = 1'b1;	
							y63 = 1'b1;	y64 = 1'b1;	
							nx_state = s1314;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x66 && x19 && ~x6 && ~x8 && ~x5 && x7 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y59 = 1'b1;	
							y60 = 1'b1;	y61 = 1'b1;	
							nx_state = s1314;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x66 && x19 && ~x6 && ~x8 && ~x5 && ~x7 )
						begin
							y5 = 1'b1;	y27 = 1'b1;	y41 = 1'b1;	
							y54 = 1'b1;	
							nx_state = s1314;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && x66 && ~x19 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y49 = 1'b1;	
							y50 = 1'b1;	
							nx_state = s1315;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && ~x66 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && ~x66 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x62 && ~x63 && ~x64 && ~x65 && ~x66 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x64 && ~x65 && ~x66 && ~x17 )
						nx_state = s1;
					else nx_state = s845;
				s846 : if( x15 )
						begin
							y46 = 1'b1;	y47 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x15 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x15 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x15 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x15 && ~x6 )
						nx_state = s1;
					else nx_state = s846;
				s847 : if( x63 && x28 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x63 && ~x28 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x63 && x15 )
						begin
							y44 = 1'b1;	y45 = 1'b1;	
							nx_state = s392;
						end
					else if( ~x63 && ~x15 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && ~x15 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && ~x15 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x63 && ~x15 && ~x6 )
						nx_state = s1;
					else nx_state = s847;
				s848 : if( 1'b1 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1129;
						end
					else nx_state = s848;
				s849 : if( 1'b1 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1130;
						end
					else nx_state = s849;
				s850 : if( x65 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x65 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else nx_state = s850;
				s851 : if( x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x18 )
						nx_state = s1;
					else if( ~x21 && x23 && x22 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x21 && x23 && ~x22 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s362;
						end
					else if( ~x21 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else nx_state = s851;
				s852 : if( 1'b1 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s365;
						end
					else nx_state = s852;
				s853 : if( x23 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s275;
						end
					else if( ~x23 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else nx_state = s853;
				s854 : if( x64 )
						begin
							y6 = 1'b1;	
							nx_state = s431;
						end
					else if( ~x64 )
						begin
							y47 = 1'b1;	y51 = 1'b1;	y61 = 1'b1;	
							y68 = 1'b1;	
							nx_state = s1316;
						end
					else nx_state = s854;
				s855 : if( 1'b1 )
						begin
							y38 = 1'b1;	
							nx_state = s532;
						end
					else nx_state = s855;
				s856 : if( 1'b1 )
						begin
							y27 = 1'b1;	
							nx_state = s893;
						end
					else nx_state = s856;
				s857 : if( x30 )
						begin
							y24 = 1'b1;	
							nx_state = s1317;
						end
					else if( ~x30 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else nx_state = s857;
				s858 : if( x68 && x15 && x10 && x11 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s600;
						end
					else if( x68 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s601;
						end
					else if( x68 && x15 && x10 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y13 = 1'b1;	
							nx_state = s600;
						end
					else if( x68 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s260;
						end
					else if( x68 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s602;
						end
					else if( x68 && ~x15 && x16 && x10 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x68 && ~x15 && x16 && x10 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x68 && ~x15 && x16 && x10 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x68 && ~x15 && x16 && x10 && ~x19 )
						nx_state = s1;
					else if( x68 && ~x15 && x16 && ~x10 && x12 && x11 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s603;
						end
					else if( x68 && ~x15 && x16 && ~x10 && x12 && ~x11 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x68 && ~x15 && x16 && ~x10 && x12 && ~x11 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x68 && ~x15 && x16 && ~x10 && x12 && ~x11 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x68 && ~x15 && x16 && ~x10 && x12 && ~x11 && ~x19 )
						nx_state = s1;
					else if( x68 && ~x15 && x16 && ~x10 && ~x12 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x68 && ~x15 && x16 && ~x10 && ~x12 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x68 && ~x15 && x16 && ~x10 && ~x12 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x68 && ~x15 && x16 && ~x10 && ~x12 && ~x19 )
						nx_state = s1;
					else if( x68 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s604;
						end
					else if( ~x68 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s70;
						end
					else nx_state = s858;
				s859 : if( x19 && x20 && x11 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x19 && x20 && ~x11 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x19 && x20 && ~x11 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x19 && x20 && ~x11 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x19 && x20 && ~x11 && ~x5 )
						nx_state = s1;
					else if( x19 && ~x20 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x19 && ~x20 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x19 && ~x20 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x19 && ~x20 && ~x5 )
						nx_state = s1;
					else if( ~x19 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x19 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x19 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x19 && ~x5 )
						nx_state = s1;
					else nx_state = s859;
				s860 : if( x19 && x17 && x20 && x14 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x19 && x17 && x20 && ~x14 )
						begin
							y4 = 1'b1;	y29 = 1'b1;	y32 = 1'b1;	
							nx_state = s863;
						end
					else if( x19 && x17 && ~x20 && x14 )
						begin
							y4 = 1'b1;	y18 = 1'b1;	y29 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s863;
						end
					else if( x19 && x17 && ~x20 && ~x14 && x15 )
						begin
							y16 = 1'b1;	y28 = 1'b1;	
							nx_state = s865;
						end
					else if( x19 && x17 && ~x20 && ~x14 && ~x15 && x16 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	y32 = 1'b1;	
							nx_state = s863;
						end
					else if( x19 && x17 && ~x20 && ~x14 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s863;
						end
					else if( x19 && ~x17 && x18 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	y19 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s861;
						end
					else if( x19 && ~x17 && ~x18 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x19 && x20 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x19 && ~x20 && x17 && x16 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x19 && ~x20 && x17 && ~x16 && x15 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x19 && ~x20 && x17 && ~x16 && ~x15 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x19 && ~x20 && ~x17 && x18 && x4 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s868;
						end
					else if( ~x19 && ~x20 && ~x17 && x18 && ~x4 )
						begin
							y7 = 1'b1;	
							nx_state = s747;
						end
					else if( ~x19 && ~x20 && ~x17 && ~x18 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else nx_state = s860;
				s861 : if( x19 && x11 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x19 && ~x11 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x19 && ~x11 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x19 && ~x11 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x19 && ~x11 && ~x5 )
						nx_state = s1;
					else if( ~x19 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x19 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x19 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x19 && ~x5 )
						nx_state = s1;
					else nx_state = s861;
				s862 : if( x19 && x14 && x20 )
						begin
							y7 = 1'b1;	
							nx_state = s747;
						end
					else if( x19 && x14 && ~x20 )
						begin
							y2 = 1'b1;	y21 = 1'b1;	
							nx_state = s1318;
						end
					else if( x19 && ~x14 )
						begin
							y7 = 1'b1;	
							nx_state = s747;
						end
					else if( ~x19 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x19 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x19 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x19 && ~x5 )
						nx_state = s1;
					else nx_state = s862;
				s863 : if( x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x5 )
						nx_state = s1;
					else nx_state = s863;
				s864 : if( x70 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x70 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x70 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x70 && ~x5 )
						nx_state = s1;
					else nx_state = s864;
				s865 : if( x19 && x20 && x9 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s868;
						end
					else if( x19 && x20 && ~x9 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x19 && ~x20 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x19 && ~x20 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( x19 && ~x20 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x19 && ~x20 && ~x5 )
						nx_state = s1;
					else if( ~x19 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x19 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x19 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x19 && ~x5 )
						nx_state = s1;
					else nx_state = s865;
				s866 : if( 1'b1 )
						begin
							y14 = 1'b1;	
							nx_state = s1319;
						end
					else nx_state = s866;
				s867 : if( x44 && x19 && x28 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( x44 && x19 && x28 && ~x1 && x35 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x44 && x19 && x28 && ~x1 && ~x35 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s870;
						end
					else if( x44 && x19 && ~x28 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x44 && ~x19 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s870;
						end
					else if( ~x44 && x13 && x23 && x51 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x44 && x13 && x23 && ~x51 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x44 && x13 && ~x23 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x44 && ~x13 && x28 && x35 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x44 && ~x13 && x28 && x35 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( ~x44 && ~x13 && x28 && ~x35 && x45 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x44 && ~x13 && x28 && ~x35 && ~x45 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( ~x44 && ~x13 && ~x28 && x6 && x35 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s907;
						end
					else if( ~x44 && ~x13 && ~x28 && x6 && ~x35 && x45 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x44 && ~x13 && ~x28 && x6 && ~x35 && ~x45 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( ~x44 && ~x13 && ~x28 && ~x6 && x39 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( ~x44 && ~x13 && ~x28 && ~x6 && ~x39 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s737;
						end
					else nx_state = s867;
				s868 : if( x69 && x17 && x19 && x20 && x14 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x69 && x17 && x19 && x20 && ~x14 && x16 )
						begin
							y4 = 1'b1;	y29 = 1'b1;	y32 = 1'b1;	
							nx_state = s863;
						end
					else if( x69 && x17 && x19 && x20 && ~x14 && ~x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && x17 && x19 && ~x20 && x14 )
						begin
							y4 = 1'b1;	y18 = 1'b1;	y29 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s863;
						end
					else if( x69 && x17 && x19 && ~x20 && ~x14 && x16 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	y32 = 1'b1;	
							nx_state = s863;
						end
					else if( x69 && x17 && x19 && ~x20 && ~x14 && ~x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s863;
						end
					else if( x69 && x17 && ~x19 && x16 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s863;
						end
					else if( x69 && x17 && ~x19 && ~x16 && x20 )
						begin
							y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s863;
						end
					else if( x69 && x17 && ~x19 && ~x16 && ~x20 && x15 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x69 && x17 && ~x19 && ~x16 && ~x20 && ~x15 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x69 && ~x17 && x18 && x19 && x14 && x16 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	y19 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s861;
						end
					else if( x69 && ~x17 && x18 && x19 && x14 && ~x16 )
						begin
							y2 = 1'b1;	y21 = 1'b1;	
							nx_state = s1318;
						end
					else if( x69 && ~x17 && x18 && x19 && ~x14 )
						begin
							y7 = 1'b1;	
							nx_state = s747;
						end
					else if( x69 && ~x17 && x18 && ~x19 )
						begin
							y7 = 1'b1;	
							nx_state = s747;
						end
					else if( x69 && ~x17 && ~x18 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && x44 && x12 && x27 && x33 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( ~x69 && x44 && x12 && x27 && ~x33 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x69 && x44 && x12 && x27 && ~x33 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x69 && x44 && x12 && ~x27 && x37 && x29 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s871;
						end
					else if( ~x69 && x44 && x12 && ~x27 && x37 && ~x29 )
						nx_state = s868;
					else if( ~x69 && x44 && x12 && ~x27 && ~x37 )
						nx_state = s868;
					else if( ~x69 && x44 && ~x12 && x29 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( ~x69 && x44 && ~x12 && ~x29 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s910;
						end
					else if( ~x69 && ~x44 && x17 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s913;
						end
					else if( ~x69 && ~x44 && ~x17 && x49 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( ~x69 && ~x44 && ~x17 && ~x49 )
						nx_state = s868;
					else nx_state = s868;
				s869 : if( x62 && x2 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( x62 && ~x2 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s875;
						end
					else if( ~x62 && x64 && x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x62 && x64 && ~x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s915;
						end
					else if( ~x62 && ~x64 && x33 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x62 && ~x64 && ~x33 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s915;
						end
					else nx_state = s869;
				s870 : if( x44 && x19 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s907;
						end
					else if( x44 && x19 && ~x13 && x32 && x18 && x12 )
						nx_state = s870;
					else if( x44 && x19 && ~x13 && x32 && x18 && ~x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s915;
						end
					else if( x44 && x19 && ~x13 && x32 && ~x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x44 && x19 && ~x13 && ~x32 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x44 && ~x19 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x44 && x17 && x19 && x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s737;
						end
					else if( ~x44 && x17 && x19 && ~x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s915;
						end
					else if( ~x44 && x17 && ~x19 )
						nx_state = s870;
					else if( ~x44 && ~x17 && x20 )
						begin
							y11 = 1'b1;	
							nx_state = s250;
						end
					else if( ~x44 && ~x17 && ~x20 && x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x44 && ~x17 && ~x20 && ~x2 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s867;
						end
					else nx_state = s870;
				s871 : if( x44 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else if( x44 && ~x5 && x34 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s737;
						end
					else if( x44 && ~x5 && ~x34 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( ~x44 && x35 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x44 && ~x35 && x13 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s868;
						end
					else if( ~x44 && ~x35 && ~x13 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else nx_state = s871;
				s872 : if( 1'b1 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else nx_state = s872;
				s873 : if( x18 && x19 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y21 = 1'b1;	
							nx_state = s820;
						end
					else if( x18 && ~x19 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	y21 = 1'b1;	
							y42 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x18 && x19 )
						begin
							y23 = 1'b1;	y29 = 1'b1;	y48 = 1'b1;	
							nx_state = s1320;
						end
					else if( ~x18 && ~x19 && x2 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s1321;
						end
					else if( ~x18 && ~x19 && ~x2 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	y34 = 1'b1;	
							nx_state = s820;
						end
					else nx_state = s873;
				s874 : if( x61 && x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s965;
						end
					else if( x61 && ~x5 && x34 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( x61 && ~x5 && ~x34 )
						begin
							y10 = 1'b1;	
							nx_state = s841;
						end
					else if( ~x61 && x35 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( ~x61 && ~x35 && x13 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s215;
						end
					else if( ~x61 && ~x35 && ~x13 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s320;
						end
					else nx_state = s874;
				s875 : if( x61 && x25 && x22 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( x61 && x25 && ~x22 && x6 && x8 )
						begin
							y10 = 1'b1;	
							nx_state = s841;
						end
					else if( x61 && x25 && ~x22 && x6 && ~x8 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( x61 && x25 && ~x22 && ~x6 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s733;
						end
					else if( x61 && ~x25 && x29 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							nx_state = s869;
						end
					else if( x61 && ~x25 && ~x29 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s874;
						end
					else if( ~x61 && x38 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s733;
						end
					else if( ~x61 && ~x38 && x50 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x61 && ~x38 && ~x50 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else nx_state = s875;
				s876 : if( x15 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s761;
						end
					else if( x15 && ~x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s1322;
						end
					else if( ~x15 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s1322;
						end
					else nx_state = s876;
				s877 : if( x18 && x19 && x14 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( x18 && x19 && ~x14 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x18 && x19 && ~x14 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x18 && x19 && ~x14 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x18 && x19 && ~x14 && ~x11 )
						nx_state = s1;
					else if( x18 && ~x19 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x18 && ~x19 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x18 && ~x19 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x18 && ~x19 && ~x11 )
						nx_state = s1;
					else if( ~x18 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x18 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x18 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x18 && ~x11 )
						nx_state = s1;
					else nx_state = s877;
				s878 : if( 1'b1 )
						begin
							y30 = 1'b1;	
							nx_state = s291;
						end
					else nx_state = s878;
				s879 : if( x1 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s178;
						end
					else nx_state = s879;
				s880 : if( x19 && x18 && x14 )
						begin
							y7 = 1'b1;	
							nx_state = s747;
						end
					else if( x19 && x18 && ~x14 && x17 )
						begin
							y7 = 1'b1;	
							nx_state = s747;
						end
					else if( x19 && x18 && ~x14 && ~x17 && x20 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x19 && x18 && ~x14 && ~x17 && ~x20 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else if( x19 && ~x18 )
						begin
							y7 = 1'b1;	
							nx_state = s747;
						end
					else if( ~x19 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else nx_state = s880;
				s881 : if( 1'b1 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s818;
						end
					else nx_state = s881;
				s882 : if( x69 && x13 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s994;
						end
					else if( x69 && ~x13 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s995;
						end
					else if( ~x69 && x39 && x1 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y33 = 1'b1;	
							nx_state = s506;
						end
					else if( ~x69 && x39 && ~x1 && x4 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y31 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s1126;
						end
					else if( ~x69 && x39 && ~x1 && ~x4 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s501;
						end
					else if( ~x69 && ~x39 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else nx_state = s882;
				s883 : if( x69 && x14 )
						begin
							y3 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							nx_state = s881;
						end
					else if( x69 && ~x14 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s882;
						end
					else if( ~x69 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y33 = 1'b1;	
							nx_state = s1236;
						end
					else nx_state = s883;
				s884 : if( x69 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s498;
						end
					else if( ~x69 && x55 && x40 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && x55 && ~x40 && x37 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( ~x69 && x55 && ~x40 && ~x37 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s818;
						end
					else if( ~x69 && ~x55 && x10 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && ~x55 && ~x10 && x42 && x32 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s882;
						end
					else if( ~x69 && ~x55 && ~x10 && x42 && ~x32 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x69 && ~x55 && ~x10 && x42 && ~x32 && ~x3 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x69 && ~x55 && ~x10 && ~x42 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else nx_state = s884;
				s885 : if( x63 && x20 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							nx_state = s1323;
						end
					else if( x63 && ~x20 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s936;
						end
					else if( ~x63 )
						begin
							y33 = 1'b1;	
							nx_state = s589;
						end
					else nx_state = s885;
				s886 : if( x64 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( ~x64 && x4 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	y29 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x64 && ~x4 && x31 && x30 )
						begin
							y5 = 1'b1;	
							nx_state = s937;
						end
					else if( ~x64 && ~x4 && x31 && ~x30 )
						begin
							y5 = 1'b1;	
							nx_state = s562;
						end
					else if( ~x64 && ~x4 && ~x31 && x30 )
						begin
							y5 = 1'b1;	
							nx_state = s945;
						end
					else if( ~x64 && ~x4 && ~x31 && ~x30 )
						begin
							y5 = 1'b1;	
							nx_state = s950;
						end
					else nx_state = s886;
				s887 : if( 1'b1 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else nx_state = s887;
				s888 : if( x63 )
						begin
							y25 = 1'b1;	y27 = 1'b1;	y48 = 1'b1;	
							nx_state = s1324;
						end
					else if( ~x63 )
						begin
							y48 = 1'b1;	y53 = 1'b1;	y61 = 1'b1;	
							nx_state = s1325;
						end
					else nx_state = s888;
				s889 : if( 1'b1 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else nx_state = s889;
				s890 : if( x20 && x15 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s556;
						end
					else if( x20 && ~x15 && x16 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s131;
						end
					else if( x20 && ~x15 && ~x16 )
						begin
							y7 = 1'b1;	y12 = 1'b1;	
							nx_state = s610;
						end
					else if( ~x20 && x21 && x17 && x15 && x8 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x20 && x21 && x17 && x15 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s556;
						end
					else if( ~x20 && x21 && x17 && ~x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x20 && x21 && x17 && ~x15 && ~x16 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x20 && x21 && ~x17 )
						nx_state = s47;
					else if( ~x20 && ~x21 && x3 )
						nx_state = s47;
					else if( ~x20 && ~x21 && ~x3 && x18 && x15 && x8 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x20 && ~x21 && ~x3 && x18 && x15 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s556;
						end
					else if( ~x20 && ~x21 && ~x3 && x18 && ~x15 && x16 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x20 && ~x21 && ~x3 && x18 && ~x15 && ~x16 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x20 && ~x21 && ~x3 && ~x18 )
						nx_state = s118;
					else nx_state = s890;
				s891 : if( x62 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x62 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x62 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( x62 && ~x27 )
						nx_state = s1;
					else if( ~x62 && x63 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x62 && x63 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x62 && x63 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x62 && x63 && ~x14 )
						nx_state = s1;
					else if( ~x62 && ~x63 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x62 && ~x63 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x62 && ~x63 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x62 && ~x63 && ~x18 )
						nx_state = s1;
					else nx_state = s891;
				s892 : if( x63 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x63 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y55 = 1'b1;	
							nx_state = s1078;
						end
					else nx_state = s892;
				s893 : if( x63 && x10 && x2 )
						nx_state = s1;
					else if( x63 && x10 && ~x2 && x3 && x4 && x5 && x1 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x63 && x10 && ~x2 && x3 && x4 && x5 && ~x1 )
						begin
							y41 = 1'b1;	y45 = 1'b1;	y46 = 1'b1;	
							nx_state = s654;
						end
					else if( x63 && x10 && ~x2 && x3 && x4 && ~x5 && x1 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( x63 && x10 && ~x2 && x3 && x4 && ~x5 && ~x1 )
						begin
							y39 = 1'b1;	y43 = 1'b1;	y44 = 1'b1;	
							nx_state = s654;
						end
					else if( x63 && x10 && ~x2 && x3 && ~x4 && x5 && x1 )
						begin
							y51 = 1'b1;	
							nx_state = s655;
						end
					else if( x63 && x10 && ~x2 && x3 && ~x4 && x5 && ~x1 )
						begin
							y41 = 1'b1;	y42 = 1'b1;	
							nx_state = s654;
						end
					else if( x63 && x10 && ~x2 && x3 && ~x4 && ~x5 && x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y48 = 1'b1;	
							y50 = 1'b1;	
							nx_state = s654;
						end
					else if( x63 && x10 && ~x2 && x3 && ~x4 && ~x5 && ~x1 )
						begin
							y39 = 1'b1;	y40 = 1'b1;	
							nx_state = s654;
						end
					else if( x63 && x10 && ~x2 && ~x3 && x4 && x5 && x1 && x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s651;
						end
					else if( x63 && x10 && ~x2 && ~x3 && x4 && x5 && x1 && ~x6 && x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s651;
						end
					else if( x63 && x10 && ~x2 && ~x3 && x4 && x5 && x1 && ~x6 && ~x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s652;
						end
					else if( x63 && x10 && ~x2 && ~x3 && x4 && x5 && ~x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y47 = 1'b1;	y48 = 1'b1;	
							nx_state = s654;
						end
					else if( x63 && x10 && ~x2 && ~x3 && x4 && ~x5 && x1 && x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s653;
						end
					else if( x63 && x10 && ~x2 && ~x3 && x4 && ~x5 && x1 && ~x6 && x7 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s653;
						end
					else if( x63 && x10 && ~x2 && ~x3 && x4 && ~x5 && x1 && ~x6 && ~x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s654;
						end
					else if( x63 && x10 && ~x2 && ~x3 && x4 && ~x5 && ~x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y48 = 1'b1;	y49 = 1'b1;	
							nx_state = s654;
						end
					else if( x63 && x10 && ~x2 && ~x3 && ~x4 && x1 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s654;
						end
					else if( x63 && x10 && ~x2 && ~x3 && ~x4 && x1 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s654;
						end
					else if( x63 && x10 && ~x2 && ~x3 && ~x4 && ~x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y32 = 1'b1;	y48 = 1'b1;	
							nx_state = s654;
						end
					else if( x63 && ~x10 )
						begin
							y28 = 1'b1;	
							nx_state = s1326;
						end
					else if( ~x63 && x67 && x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x63 && x67 && x11 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x63 && x67 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x63 && x67 && ~x11 )
						nx_state = s1;
					else if( ~x63 && ~x67 )
						begin
							y38 = 1'b1;	
							nx_state = s532;
						end
					else nx_state = s893;
				s894 : if( x21 )
						nx_state = s1;
					else if( ~x21 && x22 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else if( ~x21 && ~x22 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s236;
						end
					else if( ~x21 && ~x22 && ~x5 && x7 && x18 && x15 )
						begin
							y8 = 1'b1;	y18 = 1'b1;	
							nx_state = s152;
						end
					else if( ~x21 && ~x22 && ~x5 && x7 && x18 && ~x15 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s6;
						end
					else if( ~x21 && ~x22 && ~x5 && x7 && ~x18 && x19 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s835;
						end
					else if( ~x21 && ~x22 && ~x5 && x7 && ~x18 && x19 && ~x15 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x21 && ~x22 && ~x5 && x7 && ~x18 && ~x19 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x21 && ~x22 && ~x5 && ~x7 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s376;
						end
					else nx_state = s894;
				s895 : if( x70 && x3 && x4 && x33 && x32 && x13 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s967;
						end
					else if( x70 && x3 && x4 && x33 && x32 && x13 && ~x15 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s968;
						end
					else if( x70 && x3 && x4 && x33 && x32 && ~x13 && x14 && x15 && x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s970;
						end
					else if( x70 && x3 && x4 && x33 && x32 && ~x13 && x14 && x15 && ~x12 && x10 && x11 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s470;
						end
					else if( x70 && x3 && x4 && x33 && x32 && ~x13 && x14 && x15 && ~x12 && x10 && ~x11 )
						nx_state = s1;
					else if( x70 && x3 && x4 && x33 && x32 && ~x13 && x14 && x15 && ~x12 && ~x10 )
						nx_state = s1;
					else if( x70 && x3 && x4 && x33 && x32 && ~x13 && x14 && ~x15 && x11 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s971;
						end
					else if( x70 && x3 && x4 && x33 && x32 && ~x13 && x14 && ~x15 && ~x11 && x10 && x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s470;
						end
					else if( x70 && x3 && x4 && x33 && x32 && ~x13 && x14 && ~x15 && ~x11 && x10 && ~x12 )
						nx_state = s1;
					else if( x70 && x3 && x4 && x33 && x32 && ~x13 && x14 && ~x15 && ~x11 && ~x10 )
						nx_state = s1;
					else if( x70 && x3 && x4 && x33 && x32 && ~x13 && ~x14 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x70 && x3 && x4 && x33 && x32 && ~x13 && ~x14 && ~x15 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s311;
						end
					else if( x70 && x3 && x4 && x33 && ~x32 )
						begin
							y15 = 1'b1;	
							nx_state = s22;
						end
					else if( x70 && x3 && x4 && ~x33 && x6 && x32 && x14 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1327;
						end
					else if( x70 && x3 && x4 && ~x33 && x6 && x32 && ~x14 )
						begin
							y6 = 1'b1;	y47 = 1'b1;	
							nx_state = s1328;
						end
					else if( x70 && x3 && x4 && ~x33 && x6 && ~x32 )
						begin
							y6 = 1'b1;	y35 = 1'b1;	y40 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s355;
						end
					else if( x70 && x3 && x4 && ~x33 && ~x6 )
						begin
							y15 = 1'b1;	
							nx_state = s22;
						end
					else if( x70 && x3 && ~x4 )
						begin
							y15 = 1'b1;	
							nx_state = s356;
						end
					else if( x70 && ~x3 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							nx_state = s1329;
						end
					else if( ~x70 && x21 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s358;
						end
					else if( ~x70 && ~x21 && x22 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x21 && x22 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x21 && x22 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x70 && ~x21 && x22 && ~x5 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 && x19 && x15 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s169;
						end
					else if( ~x70 && ~x21 && ~x22 && x19 && ~x15 && x12 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							nx_state = s315;
						end
					else if( ~x70 && ~x21 && ~x22 && x19 && ~x15 && ~x12 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s169;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x19 && x20 && x14 && x15 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s169;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x19 && x20 && x14 && ~x15 && x18 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s169;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x19 && x20 && x14 && ~x15 && ~x18 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x19 && x20 && x14 && ~x15 && ~x18 && x4 && ~x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x19 && x20 && x14 && ~x15 && ~x18 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 && ~x19 && x20 && x14 && ~x15 && ~x18 && ~x4 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 && ~x19 && x20 && ~x14 && x15 && x16 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s169;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x19 && x20 && ~x14 && x15 && ~x16 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x19 && x20 && ~x14 && x15 && ~x16 && x4 && ~x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x19 && x20 && ~x14 && x15 && ~x16 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 && ~x19 && x20 && ~x14 && x15 && ~x16 && ~x4 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 && ~x19 && x20 && ~x14 && ~x15 && x17 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s169;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x19 && x20 && ~x14 && ~x15 && ~x17 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x19 && x20 && ~x14 && ~x15 && ~x17 && x4 && ~x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x19 && x20 && ~x14 && ~x15 && ~x17 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 && ~x19 && x20 && ~x14 && ~x15 && ~x17 && ~x4 )
						nx_state = s1;
					else if( ~x70 && ~x21 && ~x22 && ~x19 && ~x20 && x12 )
						begin
							y6 = 1'b1;	y21 = 1'b1;	
							nx_state = s684;
						end
					else if( ~x70 && ~x21 && ~x22 && ~x19 && ~x20 && ~x12 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s169;
						end
					else nx_state = s895;
				s896 : if( 1'b1 )
						begin
							y21 = 1'b1;	
							nx_state = s90;
						end
					else nx_state = s896;
				s897 : if( x69 && x62 && x17 )
						begin
							y14 = 1'b1;	
							nx_state = s227;
						end
					else if( x69 && x62 && ~x17 )
						begin
							y1 = 1'b1;	y12 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1188;
						end
					else if( x69 && ~x62 && x63 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( x69 && ~x62 && ~x63 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s328;
						end
					else if( ~x69 && x63 && x4 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x69 && x63 && ~x4 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s577;
						end
					else if( ~x69 && ~x63 && x8 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( ~x69 && ~x63 && ~x8 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s1330;
						end
					else nx_state = s897;
				s898 : if( x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s1331;
						end
					else if( ~x3 && x8 && x21 && x16 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x3 && x8 && x21 && x16 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s261;
						end
					else if( ~x3 && x8 && x21 && ~x16 && x17 && x18 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s810;
						end
					else if( ~x3 && x8 && x21 && ~x16 && x17 && x18 && ~x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( ~x3 && x8 && x21 && ~x16 && x17 && ~x18 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( ~x3 && x8 && x21 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x3 && x8 && ~x21 && x22 && x16 && x19 && x18 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x3 && x8 && ~x21 && x22 && x16 && x19 && x18 && ~x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s264;
						end
					else if( ~x3 && x8 && ~x21 && x22 && x16 && x19 && ~x18 && x13 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x3 && x8 && ~x21 && x22 && x16 && x19 && ~x18 && ~x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x3 && x8 && ~x21 && x22 && x16 && ~x19 && x13 )
						begin
							y3 = 1'b1;	y16 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x3 && x8 && ~x21 && x22 && x16 && ~x19 && ~x13 && x18 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x3 && x8 && ~x21 && x22 && x16 && ~x19 && ~x13 && ~x18 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x3 && x8 && ~x21 && x22 && ~x16 && x17 && x19 && x18 && x10 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else if( ~x3 && x8 && ~x21 && x22 && ~x16 && x17 && x19 && x18 && ~x10 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x3 && x8 && ~x21 && x22 && ~x16 && x17 && x19 && ~x18 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else if( ~x3 && x8 && ~x21 && x22 && ~x16 && x17 && x19 && ~x18 && ~x13 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x3 && x8 && ~x21 && x22 && ~x16 && x17 && ~x19 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else if( ~x3 && x8 && ~x21 && x22 && ~x16 && x17 && ~x19 && ~x13 && x18 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x3 && x8 && ~x21 && x22 && ~x16 && x17 && ~x19 && ~x13 && ~x18 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x3 && x8 && ~x21 && x22 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && x19 && x17 && x13 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && x19 && x17 && ~x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && x19 && ~x17 && x18 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && x19 && ~x17 && x18 && ~x13 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && x19 && ~x17 && ~x18 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && ~x19 && x16 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && ~x19 && x16 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s261;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && ~x19 && ~x16 && x17 && x20 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && ~x19 && ~x16 && x17 && ~x20 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s810;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && ~x19 && ~x16 && x17 && ~x20 && ~x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && ~x19 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x3 && ~x8 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s1332;
						end
					else nx_state = s898;
				s899 : if( x68 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x68 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s497;
						end
					else nx_state = s899;
				s900 : if( x16 && x15 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s438;
						end
					else if( x16 && ~x15 && x4 && x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s438;
						end
					else if( x16 && ~x15 && x4 && ~x5 && x1 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s438;
						end
					else if( x16 && ~x15 && x4 && ~x5 && ~x1 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s194;
						end
					else if( x16 && ~x15 && ~x4 && x1 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s438;
						end
					else if( x16 && ~x15 && ~x4 && ~x1 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s448;
						end
					else if( ~x16 && x15 && x3 && x2 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s451;
						end
					else if( ~x16 && x15 && x3 && ~x2 )
						nx_state = s900;
					else if( ~x16 && x15 && ~x3 && x4 && x2 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s194;
						end
					else if( ~x16 && x15 && ~x3 && x4 && ~x2 )
						nx_state = s900;
					else if( ~x16 && x15 && ~x3 && ~x4 && x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x16 && x15 && ~x3 && ~x4 && ~x2 )
						nx_state = s900;
					else if( ~x16 && ~x15 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s438;
						end
					else nx_state = s900;
				s901 : if( x16 && x15 && x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( x16 && x15 && ~x5 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s627;
						end
					else if( x16 && ~x15 && x4 && x5 && x2 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s195;
						end
					else if( x16 && ~x15 && x4 && x5 && ~x2 && x1 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s448;
						end
					else if( x16 && ~x15 && x4 && x5 && ~x2 && ~x1 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else if( x16 && ~x15 && x4 && ~x5 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s195;
						end
					else if( x16 && ~x15 && ~x4 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s195;
						end
					else if( ~x16 && x15 && x13 && x11 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s436;
						end
					else if( ~x16 && x15 && x13 && ~x11 && x6 && x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s194;
						end
					else if( ~x16 && x15 && x13 && ~x11 && x6 && ~x4 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x16 && x15 && x13 && ~x11 && ~x6 && x5 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else if( ~x16 && x15 && x13 && ~x11 && ~x6 && ~x5 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s900;
						end
					else if( ~x16 && x15 && ~x13 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s193;
						end
					else if( ~x16 && x15 && ~x13 && ~x14 && x9 )
						begin
							y10 = 1'b1;	
							nx_state = s193;
						end
					else if( ~x16 && x15 && ~x13 && ~x14 && ~x9 && x6 && x2 )
						begin
							y10 = 1'b1;	
							nx_state = s193;
						end
					else if( ~x16 && x15 && ~x13 && ~x14 && ~x9 && x6 && ~x2 )
						nx_state = s901;
					else if( ~x16 && x15 && ~x13 && ~x14 && ~x9 && ~x6 && x8 )
						begin
							y10 = 1'b1;	
							nx_state = s193;
						end
					else if( ~x16 && x15 && ~x13 && ~x14 && ~x9 && ~x6 && ~x8 )
						nx_state = s901;
					else if( ~x16 && ~x15 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else nx_state = s901;
				s902 : if( x42 && x13 && x43 && x35 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( x42 && x13 && x43 && ~x35 )
						nx_state = s902;
					else if( x42 && x13 && ~x43 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( x42 && x13 && ~x43 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( x42 && x13 && ~x43 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( x42 && x13 && ~x43 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x42 && x13 && ~x43 && x15 && ~x47 && ~x1 )
						nx_state = s902;
					else if( x42 && x13 && ~x43 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x42 && x13 && ~x43 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x42 && x13 && ~x43 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x42 && ~x13 && x35 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( x42 && ~x13 && ~x35 )
						nx_state = s902;
					else if( ~x42 && x44 && x12 && x35 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x42 && x44 && x12 && ~x35 )
						nx_state = s902;
					else if( ~x42 && x44 && ~x12 && x14 && x35 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x42 && x44 && ~x12 && x14 && ~x35 )
						nx_state = s902;
					else if( ~x42 && x44 && ~x12 && ~x14 && x15 && x47 && x36 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x42 && x44 && ~x12 && ~x14 && x15 && x47 && ~x36 && x6 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x42 && x44 && ~x12 && ~x14 && x15 && x47 && ~x36 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x42 && x44 && ~x12 && ~x14 && x15 && ~x47 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && x44 && ~x12 && ~x14 && x15 && ~x47 && ~x1 )
						nx_state = s902;
					else if( ~x42 && x44 && ~x12 && ~x14 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && x44 && ~x12 && ~x14 && ~x15 && ~x16 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x42 && x44 && ~x12 && ~x14 && ~x15 && ~x16 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x42 && ~x44 && x35 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x42 && ~x44 && ~x35 )
						nx_state = s902;
					else nx_state = s902;
				s903 : if( x64 && x40 && x22 && x2 && x33 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( x64 && x40 && x22 && x2 && ~x33 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x64 && x40 && x22 && x2 && ~x33 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x64 && x40 && x22 && ~x2 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x64 && x40 && ~x22 && x31 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x64 && x40 && ~x22 && ~x31 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x64 && ~x40 && x46 && x3 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( x64 && ~x40 && x46 && x3 && ~x23 )
						nx_state = s903;
					else if( x64 && ~x40 && x46 && ~x3 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x64 && ~x40 && ~x46 && x2 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( x64 && ~x40 && ~x46 && x2 && ~x23 )
						nx_state = s903;
					else if( x64 && ~x40 && ~x46 && ~x2 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x64 && x44 && x22 && x2 && x33 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( ~x64 && x44 && x22 && x2 && ~x33 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x64 && x44 && x22 && x2 && ~x33 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x64 && x44 && x22 && ~x2 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x64 && x44 && ~x22 && x31 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x64 && x44 && ~x22 && ~x31 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x64 && ~x44 && x46 && x3 && x23 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s871;
						end
					else if( ~x64 && ~x44 && x46 && x3 && ~x23 )
						nx_state = s903;
					else if( ~x64 && ~x44 && x46 && ~x3 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x64 && ~x44 && ~x46 && x33 && x23 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s871;
						end
					else if( ~x64 && ~x44 && ~x46 && x33 && ~x23 )
						nx_state = s903;
					else if( ~x64 && ~x44 && ~x46 && ~x33 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else nx_state = s903;
				s904 : if( x16 && x37 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	y34 = 1'b1;	
							nx_state = s904;
						end
					else if( x16 && ~x37 && x39 && x19 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( x16 && ~x37 && x39 && ~x19 && x26 && x5 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s734;
						end
					else if( x16 && ~x37 && x39 && ~x19 && x26 && ~x5 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s735;
						end
					else if( x16 && ~x37 && x39 && ~x19 && ~x26 )
						begin
							y11 = 1'b1;	y36 = 1'b1;	
							nx_state = s739;
						end
					else if( x16 && ~x37 && ~x39 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( ~x16 && x41 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x16 && ~x41 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else nx_state = s904;
				s905 : if( x55 && x45 && x8 && x41 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x55 && x45 && x8 && ~x41 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( x55 && x45 && ~x8 && x30 && x32 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s909;
						end
					else if( x55 && x45 && ~x8 && x30 && ~x32 && x4 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s734;
						end
					else if( x55 && x45 && ~x8 && x30 && ~x32 && ~x4 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s914;
						end
					else if( x55 && x45 && ~x8 && ~x30 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x55 && ~x45 && x34 && x32 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s735;
						end
					else if( x55 && ~x45 && x34 && ~x32 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x55 && ~x45 && ~x34 )
						nx_state = s905;
					else if( ~x55 && x47 && x54 && x29 && x59 && x27 )
						begin
							y13 = 1'b1;	
							nx_state = s450;
						end
					else if( ~x55 && x47 && x54 && x29 && x59 && ~x27 )
						nx_state = s905;
					else if( ~x55 && x47 && x54 && x29 && ~x59 && x27 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x55 && x47 && x54 && x29 && ~x59 && ~x27 )
						nx_state = s905;
					else if( ~x55 && x47 && x54 && ~x29 && x33 && x27 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x55 && x47 && x54 && ~x29 && x33 && ~x27 )
						nx_state = s905;
					else if( ~x55 && x47 && x54 && ~x29 && ~x33 && x57 && x27 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( ~x55 && x47 && x54 && ~x29 && ~x33 && x57 && ~x27 )
						nx_state = s905;
					else if( ~x55 && x47 && x54 && ~x29 && ~x33 && ~x57 && x27 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x55 && x47 && x54 && ~x29 && ~x33 && ~x57 && ~x27 )
						nx_state = s905;
					else if( ~x55 && x47 && ~x54 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( ~x55 && ~x47 && x37 && x56 && x1 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x55 && ~x47 && x37 && x56 && ~x1 )
						nx_state = s905;
					else if( ~x55 && ~x47 && x37 && ~x56 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( ~x55 && ~x47 && ~x37 && x25 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( ~x55 && ~x47 && ~x37 && ~x25 && x36 && x35 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else if( ~x55 && ~x47 && ~x37 && ~x25 && x36 && ~x35 )
						nx_state = s905;
					else if( ~x55 && ~x47 && ~x37 && ~x25 && ~x36 && x35 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x55 && ~x47 && ~x37 && ~x25 && ~x36 && ~x35 )
						nx_state = s905;
					else nx_state = s905;
				s906 : if( x55 && x35 && x7 && x1 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s739;
						end
					else if( x55 && x35 && x7 && ~x1 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x55 && x35 && ~x7 )
						nx_state = s906;
					else if( x55 && ~x35 && x38 && x32 )
						nx_state = s906;
					else if( x55 && ~x35 && x38 && ~x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( x55 && ~x35 && ~x38 )
						nx_state = s906;
					else if( ~x55 && x34 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s908;
						end
					else if( ~x55 && ~x34 && x2 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s910;
						end
					else if( ~x55 && ~x34 && ~x2 && x28 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x55 && ~x34 && ~x2 && ~x28 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else nx_state = s906;
				s907 : if( x44 && x9 )
						begin
							y13 = 1'b1;	
							nx_state = s450;
						end
					else if( x44 && ~x9 && x3 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x44 && ~x9 && ~x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s737;
						end
					else if( ~x44 && x29 && x50 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s910;
						end
					else if( ~x44 && x29 && ~x50 )
						nx_state = s907;
					else if( ~x44 && ~x29 && x45 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x44 && ~x29 && ~x45 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s802;
						end
					else nx_state = s907;
				s908 : if( x55 && x22 && x2 && x33 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s908;
						end
					else if( x55 && x22 && x2 && ~x33 && x13 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( x55 && x22 && x2 && ~x33 && ~x13 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( x55 && x22 && ~x2 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( x55 && ~x22 && x31 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( x55 && ~x22 && ~x31 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x55 && x46 && x3 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s909;
						end
					else if( ~x55 && x46 && x3 && ~x23 )
						nx_state = s908;
					else if( ~x55 && x46 && ~x3 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( ~x55 && ~x46 && x33 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s909;
						end
					else if( ~x55 && ~x46 && x33 && ~x23 )
						nx_state = s908;
					else if( ~x55 && ~x46 && ~x33 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else nx_state = s908;
				s909 : if( x55 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s905;
						end
					else if( x55 && ~x5 && x34 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s734;
						end
					else if( x55 && ~x5 && ~x34 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s908;
						end
					else if( ~x55 && x35 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( ~x55 && ~x35 && x44 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s187;
						end
					else if( ~x55 && ~x35 && ~x44 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else nx_state = s909;
				s910 : if( x63 && x40 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s735;
						end
					else if( x63 && ~x40 && x37 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s735;
						end
					else if( x63 && ~x40 && ~x37 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s908;
						end
					else if( ~x63 && x64 && x37 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( ~x63 && x64 && ~x37 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( ~x63 && x64 && ~x37 && ~x9 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( ~x63 && ~x64 && x1 && x37 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( ~x63 && ~x64 && x1 && ~x37 && x9 )
						nx_state = s910;
					else if( ~x63 && ~x64 && x1 && ~x37 && ~x9 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x63 && ~x64 && ~x1 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( ~x63 && ~x64 && ~x1 && ~x9 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else nx_state = s910;
				s911 : if( 1'b1 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else nx_state = s911;
				s912 : if( x70 && x37 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s192;
						end
					else if( x70 && ~x37 && x9 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s192;
						end
					else if( x70 && ~x37 && ~x9 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s632;
						end
					else if( ~x70 && x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x70 && ~x4 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s732;
						end
					else nx_state = s912;
				s913 : if( x70 && x62 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s840;
						end
					else if( x70 && ~x62 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x70 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s189;
						end
					else nx_state = s913;
				s914 : if( x55 && x25 && x52 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( x55 && x25 && ~x52 && x6 && x39 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s908;
						end
					else if( x55 && x25 && ~x52 && x6 && ~x39 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s669;
						end
					else if( x55 && x25 && ~x52 && ~x6 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s735;
						end
					else if( x55 && ~x25 && x29 )
						begin
							y10 = 1'b1;	y26 = 1'b1;	y37 = 1'b1;	
							nx_state = s1184;
						end
					else if( x55 && ~x25 && ~x29 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s909;
						end
					else if( ~x55 && x38 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s735;
						end
					else if( ~x55 && ~x38 && x50 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x55 && ~x38 && ~x50 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s734;
						end
					else nx_state = s914;
				s915 : if( x64 && x40 && x25 && x22 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x64 && x40 && x25 && ~x22 && x6 && x8 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( x64 && x40 && x25 && ~x22 && x6 && ~x8 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( x64 && x40 && x25 && ~x22 && ~x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( x64 && x40 && ~x25 && x29 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							nx_state = s869;
						end
					else if( x64 && x40 && ~x25 && ~x29 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s185;
						end
					else if( x64 && ~x40 && x38 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( x64 && ~x40 && ~x38 && x50 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s108;
						end
					else if( x64 && ~x40 && ~x38 && ~x50 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s736;
						end
					else if( ~x64 && x44 && x25 && x22 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x64 && x44 && x25 && ~x22 && x6 && x8 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s903;
						end
					else if( ~x64 && x44 && x25 && ~x22 && x6 && ~x8 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s804;
						end
					else if( ~x64 && x44 && x25 && ~x22 && ~x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( ~x64 && x44 && ~x25 && x29 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							nx_state = s869;
						end
					else if( ~x64 && x44 && ~x25 && ~x29 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s871;
						end
					else if( ~x64 && ~x44 && x38 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s685;
						end
					else if( ~x64 && ~x44 && ~x38 && x50 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s867;
						end
					else if( ~x64 && ~x44 && ~x38 && ~x50 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s737;
						end
					else nx_state = s915;
				s916 : if( x16 && x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s519;
						end
					else if( x16 && ~x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s760;
						end
					else if( ~x16 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s868;
						end
					else nx_state = s916;
				s917 : if( x26 && x28 && x7 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s944;
						end
					else if( x26 && x28 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else if( x26 && ~x28 )
						nx_state = s1;
					else if( ~x26 && x27 && x25 && x9 )
						nx_state = s917;
					else if( ~x26 && x27 && x25 && ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else if( ~x26 && x27 && ~x25 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x26 && ~x27 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else nx_state = s917;
				s918 : if( x26 && x28 && x23 && x63 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s994;
						end
					else if( x26 && x28 && x23 && ~x63 && x64 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( x26 && x28 && x23 && ~x63 && ~x64 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s924;
						end
					else if( x26 && x28 && ~x23 && x25 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( x26 && x28 && ~x23 && ~x25 && x63 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( x26 && x28 && ~x23 && ~x25 && ~x63 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( x26 && ~x28 && x63 && x34 && x25 )
						nx_state = s918;
					else if( x26 && ~x28 && x63 && x34 && ~x25 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( x26 && ~x28 && x63 && ~x34 && x35 && x36 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else if( x26 && ~x28 && x63 && ~x34 && x35 && ~x36 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( x26 && ~x28 && x63 && ~x34 && ~x35 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( x26 && ~x28 && ~x63 && x3 && x25 )
						nx_state = s918;
					else if( x26 && ~x28 && ~x63 && x3 && ~x25 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( x26 && ~x28 && ~x63 && ~x3 && x4 && x5 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else if( x26 && ~x28 && ~x63 && ~x3 && x4 && ~x5 && x64 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( x26 && ~x28 && ~x63 && ~x3 && x4 && ~x5 && ~x64 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s917;
						end
					else if( x26 && ~x28 && ~x63 && ~x3 && ~x4 && x64 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( x26 && ~x28 && ~x63 && ~x3 && ~x4 && ~x64 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s944;
						end
					else if( ~x26 && x27 && x63 && x35 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else if( ~x26 && x27 && x63 && ~x35 )
						nx_state = s1;
					else if( ~x26 && x27 && ~x63 && x4 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else if( ~x26 && x27 && ~x63 && ~x4 )
						nx_state = s1;
					else if( ~x26 && ~x27 && x28 && x11 )
						nx_state = s1;
					else if( ~x26 && ~x27 && x28 && ~x11 && x63 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s679;
						end
					else if( ~x26 && ~x27 && x28 && ~x11 && ~x63 && x64 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s679;
						end
					else if( ~x26 && ~x27 && x28 && ~x11 && ~x63 && ~x64 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s1333;
						end
					else if( ~x26 && ~x27 && ~x28 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else nx_state = s918;
				s919 : if( x26 && x28 && x63 && x37 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( x26 && x28 && x63 && ~x37 && x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( x26 && x28 && x63 && ~x37 && ~x4 )
						nx_state = s1;
					else if( x26 && x28 && ~x63 && x6 && x64 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( x26 && x28 && ~x63 && x6 && ~x64 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s944;
						end
					else if( x26 && x28 && ~x63 && ~x6 && x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( x26 && x28 && ~x63 && ~x6 && ~x4 )
						nx_state = s1;
					else if( x26 && ~x28 )
						nx_state = s1;
					else if( ~x26 && x63 && x27 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s995;
						end
					else if( ~x26 && x63 && ~x27 && x28 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s1334;
						end
					else if( ~x26 && x63 && ~x27 && ~x28 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s995;
						end
					else if( ~x26 && ~x63 && x27 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else if( ~x26 && ~x63 && ~x27 && x28 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y29 = 1'b1;	
							nx_state = s1335;
						end
					else if( ~x26 && ~x63 && ~x27 && ~x28 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else nx_state = s919;
				s920 : if( x26 )
						begin
							y11 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x26 && x28 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s1336;
						end
					else if( ~x26 && x28 && ~x5 && x64 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s542;
						end
					else if( ~x26 && x28 && ~x5 && ~x64 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s801;
						end
					else if( ~x26 && ~x28 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else nx_state = s920;
				s921 : if( x26 && x21 )
						nx_state = s1;
					else if( x26 && ~x21 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else if( ~x26 && x27 )
						nx_state = s1;
					else if( ~x26 && ~x27 && x28 && x64 && x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( ~x26 && ~x27 && x28 && x64 && ~x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s922;
						end
					else if( ~x26 && ~x27 && x28 && ~x64 && x3 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s944;
						end
					else if( ~x26 && ~x27 && x28 && ~x64 && ~x3 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s923;
						end
					else if( ~x26 && ~x27 && ~x28 && x19 && x24 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s1185;
						end
					else if( ~x26 && ~x27 && ~x28 && x19 && ~x24 )
						nx_state = s1;
					else if( ~x26 && ~x27 && ~x28 && ~x19 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s920;
						end
					else nx_state = s921;
				s922 : if( x28 && x63 && x7 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s994;
						end
					else if( x28 && x63 && ~x7 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s1185;
						end
					else if( x28 && ~x63 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s635;
						end
					else if( x28 && ~x63 && ~x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s1185;
						end
					else if( ~x28 && x63 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x28 && ~x63 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else nx_state = s922;
				s923 : if( x28 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s924;
						end
					else if( x28 && ~x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s1185;
						end
					else if( ~x28 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else nx_state = s923;
				s924 : if( x26 && x8 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s944;
						end
					else if( x26 && x8 && ~x37 && x14 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s917;
						end
					else if( x26 && x8 && ~x37 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( x26 && ~x8 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s920;
						end
					else if( ~x26 && x28 )
						nx_state = s1;
					else if( ~x26 && ~x28 && x6 && x7 && x5 && x3 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s923;
						end
					else if( ~x26 && ~x28 && x6 && x7 && x5 && ~x3 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s924;
						end
					else if( ~x26 && ~x28 && x6 && x7 && x5 && ~x3 && ~x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else if( ~x26 && ~x28 && x6 && x7 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x26 && ~x28 && x6 && ~x7 && x8 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s1185;
						end
					else if( ~x26 && ~x28 && x6 && ~x7 && ~x8 && x5 && x3 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s923;
						end
					else if( ~x26 && ~x28 && x6 && ~x7 && ~x8 && x5 && ~x3 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s924;
						end
					else if( ~x26 && ~x28 && x6 && ~x7 && ~x8 && x5 && ~x3 && ~x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else if( ~x26 && ~x28 && x6 && ~x7 && ~x8 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x26 && ~x28 && ~x6 && x24 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s1185;
						end
					else if( ~x26 && ~x28 && ~x6 && ~x24 )
						nx_state = s1;
					else nx_state = s924;
				s925 : if( x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1337;
						end
					else if( ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1338;
						end
					else nx_state = s925;
				s926 : if( x22 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s1339;
						end
					else if( x22 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1091;
						end
					else if( ~x22 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s1092;
						end
					else if( ~x22 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1340;
						end
					else nx_state = s926;
				s927 : if( x16 && x15 && x5 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s194;
						end
					else if( x16 && x15 && ~x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s180;
						end
					else if( x16 && ~x15 && x4 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x16 && ~x15 && ~x4 && x2 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s451;
						end
					else if( x16 && ~x15 && ~x4 && ~x2 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s901;
						end
					else if( x16 && ~x15 && ~x4 && ~x2 && ~x1 )
						begin
							y10 = 1'b1;	
							nx_state = s193;
						end
					else if( ~x16 && x15 && x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s901;
						end
					else if( ~x16 && x15 && ~x12 )
						nx_state = s927;
					else if( ~x16 && ~x15 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s627;
						end
					else nx_state = s927;
				s928 : if( x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x15 && ~x16 && x13 && x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s194;
						end
					else if( x15 && ~x16 && x13 && ~x4 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x15 && ~x16 && ~x13 && x14 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s451;
						end
					else if( x15 && ~x16 && ~x13 && ~x14 && x9 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s451;
						end
					else if( x15 && ~x16 && ~x13 && ~x14 && ~x9 && x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s451;
						end
					else if( x15 && ~x16 && ~x13 && ~x14 && ~x9 && ~x7 && x8 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s451;
						end
					else if( x15 && ~x16 && ~x13 && ~x14 && ~x9 && ~x7 && ~x8 )
						nx_state = s928;
					else if( ~x15 && x16 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s450;
						end
					else if( ~x15 && x16 && ~x4 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x15 && ~x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else nx_state = s928;
				s929 : if( x15 && x63 && x16 && x5 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( x15 && x63 && x16 && ~x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x15 && x63 && ~x16 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( x15 && x63 && ~x16 && ~x12 )
						nx_state = s929;
					else if( x15 && ~x63 && x16 && x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( x15 && ~x63 && x16 && ~x5 && x64 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x15 && ~x63 && x16 && ~x5 && ~x64 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( x15 && ~x63 && ~x16 && x64 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( x15 && ~x63 && ~x16 && x64 && ~x12 )
						nx_state = s929;
					else if( x15 && ~x63 && ~x16 && ~x64 && x12 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s1143;
						end
					else if( x15 && ~x63 && ~x16 && ~x64 && ~x12 )
						nx_state = s929;
					else if( ~x15 && x63 && x47 && x35 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x15 && x63 && x47 && ~x35 && x33 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s322;
						end
					else if( ~x15 && x63 && x47 && ~x35 && ~x33 && x32 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( ~x15 && x63 && x47 && ~x35 && ~x33 && ~x32 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x15 && x63 && ~x47 )
						begin
							y21 = 1'b1;	y27 = 1'b1;	
							nx_state = s930;
						end
					else if( ~x15 && ~x63 && x16 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x15 && ~x63 && x16 && ~x4 && x64 && x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s326;
						end
					else if( ~x15 && ~x63 && x16 && ~x4 && x64 && ~x2 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( ~x15 && ~x63 && x16 && ~x4 && x64 && ~x2 && ~x1 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( ~x15 && ~x63 && x16 && ~x4 && ~x64 && x34 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s326;
						end
					else if( ~x15 && ~x63 && x16 && ~x4 && ~x64 && ~x34 && x37 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s1143;
						end
					else if( ~x15 && ~x63 && x16 && ~x4 && ~x64 && ~x34 && ~x37 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x15 && ~x63 && ~x16 )
						begin
							y21 = 1'b1;	y27 = 1'b1;	
							nx_state = s930;
						end
					else nx_state = s929;
				s930 : if( x16 && x63 && x46 )
						begin
							y15 = 1'b1;	y23 = 1'b1;	y31 = 1'b1;	
							nx_state = s1341;
						end
					else if( x16 && x63 && ~x46 && x2 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s440;
						end
					else if( x16 && x63 && ~x46 && ~x2 && x32 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( x16 && x63 && ~x46 && ~x2 && ~x32 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( x16 && ~x63 && x15 )
						begin
							y2 = 1'b1;	y15 = 1'b1;	y23 = 1'b1;	
							nx_state = s1342;
						end
					else if( x16 && ~x63 && ~x15 && x2 && x64 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s445;
						end
					else if( x16 && ~x63 && ~x15 && x2 && ~x64 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s931;
						end
					else if( x16 && ~x63 && ~x15 && ~x2 && x64 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( x16 && ~x63 && ~x15 && ~x2 && x64 && ~x1 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s196;
						end
					else if( x16 && ~x63 && ~x15 && ~x2 && ~x64 && x37 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s1143;
						end
					else if( x16 && ~x63 && ~x15 && ~x2 && ~x64 && ~x37 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x16 && x63 )
						begin
							y15 = 1'b1;	y23 = 1'b1;	y31 = 1'b1;	
							nx_state = s1341;
						end
					else if( ~x16 && ~x63 )
						begin
							y2 = 1'b1;	y15 = 1'b1;	y23 = 1'b1;	
							nx_state = s1342;
						end
					else nx_state = s930;
				s931 : if( x16 && x15 && x5 && x1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s326;
						end
					else if( x16 && x15 && x5 && ~x1 && x2 && x3 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s455;
						end
					else if( x16 && x15 && x5 && ~x1 && x2 && x3 && ~x4 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x16 && x15 && x5 && ~x1 && x2 && ~x3 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x16 && x15 && x5 && ~x1 && ~x2 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x16 && x15 && ~x5 && x6 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x16 && x15 && ~x5 && ~x6 && x37 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( x16 && x15 && ~x5 && ~x6 && ~x37 && x34 && x3 && x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s455;
						end
					else if( x16 && x15 && ~x5 && ~x6 && ~x37 && x34 && x3 && ~x4 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( x16 && x15 && ~x5 && ~x6 && ~x37 && x34 && ~x3 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x16 && x15 && ~x5 && ~x6 && ~x37 && ~x34 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x16 && ~x15 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s1143;
						end
					else if( ~x16 && x15 && x6 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s540;
						end
					else if( ~x16 && x15 && ~x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s446;
						end
					else if( ~x16 && ~x15 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else nx_state = s931;
				s932 : if( x15 && x16 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x15 && ~x16 && x63 && x13 && x4 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s323;
						end
					else if( x15 && ~x16 && x63 && x13 && ~x4 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x15 && ~x16 && x63 && x13 && ~x4 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x15 && ~x16 && x63 && ~x13 && x45 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s322;
						end
					else if( x15 && ~x16 && x63 && ~x13 && ~x45 && x9 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s322;
						end
					else if( x15 && ~x16 && x63 && ~x13 && ~x45 && ~x9 && x38 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s322;
						end
					else if( x15 && ~x16 && x63 && ~x13 && ~x45 && ~x9 && ~x38 && x39 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s322;
						end
					else if( x15 && ~x16 && x63 && ~x13 && ~x45 && ~x9 && ~x38 && ~x39 )
						nx_state = s932;
					else if( x15 && ~x16 && ~x63 && x13 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( x15 && ~x16 && ~x63 && x13 && ~x4 && x64 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( x15 && ~x16 && ~x63 && x13 && ~x4 && x64 && ~x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( x15 && ~x16 && ~x63 && x13 && ~x4 && ~x64 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( x15 && ~x16 && ~x63 && x13 && ~x4 && ~x64 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( x15 && ~x16 && ~x63 && ~x13 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s326;
						end
					else if( x15 && ~x16 && ~x63 && ~x13 && ~x14 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s326;
						end
					else if( x15 && ~x16 && ~x63 && ~x13 && ~x14 && ~x9 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s326;
						end
					else if( x15 && ~x16 && ~x63 && ~x13 && ~x14 && ~x9 && ~x7 && x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s326;
						end
					else if( x15 && ~x16 && ~x63 && ~x13 && ~x14 && ~x9 && ~x7 && ~x8 )
						nx_state = s932;
					else if( ~x15 && x63 && x47 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x15 && x63 && x47 && ~x4 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x15 && x63 && x47 && ~x4 && ~x32 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x15 && x63 && ~x47 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x15 && ~x63 && x16 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x15 && ~x63 && x16 && ~x4 && x64 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x15 && ~x63 && x16 && ~x4 && x64 && ~x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x15 && ~x63 && x16 && ~x4 && ~x64 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x15 && ~x63 && x16 && ~x4 && ~x64 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x15 && ~x63 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else nx_state = s932;
				s933 : if( x64 && x61 && x17 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s593;
						end
					else if( x64 && x61 && ~x17 && x57 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( x64 && x61 && ~x17 && ~x57 )
						nx_state = s933;
					else if( x64 && ~x61 && x6 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s593;
						end
					else if( x64 && ~x61 && ~x6 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s933;
						end
					else if( ~x64 && x14 && x17 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s593;
						end
					else if( ~x64 && x14 && ~x17 && x21 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( ~x64 && x14 && ~x17 && ~x21 )
						nx_state = s933;
					else if( ~x64 && ~x14 && x6 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s593;
						end
					else if( ~x64 && ~x14 && ~x6 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s933;
						end
					else nx_state = s933;
				s934 : if( x64 && x61 && x50 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s933;
						end
					else if( x64 && x61 && ~x50 )
						nx_state = s934;
					else if( x64 && ~x61 && x11 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else if( x64 && ~x61 && ~x11 && x9 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else if( x64 && ~x61 && ~x11 && ~x9 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( ~x64 && x14 && x42 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s933;
						end
					else if( ~x64 && x14 && ~x42 )
						nx_state = s934;
					else if( ~x64 && ~x14 && x11 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else if( ~x64 && ~x14 && ~x11 && x9 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else if( ~x64 && ~x14 && ~x11 && ~x9 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else nx_state = s934;
				s935 : if( x70 && x64 && x61 && x37 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( x70 && x64 && x61 && ~x37 && x9 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( x70 && x64 && x61 && ~x37 && ~x9 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && x64 && ~x61 && x10 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( x70 && x64 && ~x61 && ~x10 && x11 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s759;
						end
					else if( x70 && x64 && ~x61 && ~x10 && x11 && ~x1 && x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( x70 && x64 && ~x61 && ~x10 && x11 && ~x1 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x70 && x64 && ~x61 && ~x10 && ~x11 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x70 && ~x64 && x14 && x9 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( x70 && ~x64 && x14 && ~x9 && x37 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s202;
						end
					else if( x70 && ~x64 && x14 && ~x9 && ~x37 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x70 && ~x64 && ~x14 && x10 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( x70 && ~x64 && ~x14 && ~x10 && x11 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s759;
						end
					else if( x70 && ~x64 && ~x14 && ~x10 && x11 && ~x1 && x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s200;
						end
					else if( x70 && ~x64 && ~x14 && ~x10 && x11 && ~x1 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( x70 && ~x64 && ~x14 && ~x10 && ~x11 )
						begin
							y1 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x70 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s816;
						end
					else if( ~x70 && ~x9 && x5 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x70 && ~x9 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s203;
						end
					else nx_state = s935;
				s936 : if( 1'b1 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s426;
						end
					else nx_state = s936;
				s937 : if( x62 && x64 )
						begin
							y1 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s988;
						end
					else if( x62 && ~x64 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s1343;
						end
					else if( ~x62 && x64 && x21 && x20 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( ~x62 && x64 && x21 && ~x20 )
						begin
							y6 = 1'b1;	
							nx_state = s1049;
						end
					else if( ~x62 && x64 && ~x21 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( ~x62 && ~x64 && x30 && x31 )
						begin
							y47 = 1'b1;	y50 = 1'b1;	y61 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s1148;
						end
					else if( ~x62 && ~x64 && x30 && ~x31 )
						begin
							y47 = 1'b1;	y52 = 1'b1;	y61 = 1'b1;	
							y70 = 1'b1;	
							nx_state = s1298;
						end
					else if( ~x62 && ~x64 && ~x30 )
						begin
							y24 = 1'b1;	
							nx_state = s1317;
						end
					else nx_state = s937;
				s938 : if( x64 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y8 = 1'b1;	y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s1344;
						end
					else if( ~x64 && x19 && x20 && x5 && x6 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y23 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x64 && x19 && x20 && x5 && ~x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y25 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x64 && x19 && x20 && ~x5 )
						begin
							y3 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y30 = 1'b1;	y43 = 1'b1;	
							nx_state = s1345;
						end
					else if( ~x64 && x19 && ~x20 && x4 && x21 && x6 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s1270;
						end
					else if( ~x64 && x19 && ~x20 && x4 && x21 && x6 && ~x5 && x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x64 && x19 && ~x20 && x4 && x21 && x6 && ~x5 && ~x11 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x64 && x19 && ~x20 && x4 && x21 && x6 && ~x5 && ~x11 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x64 && x19 && ~x20 && x4 && x21 && x6 && ~x5 && ~x11 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x64 && x19 && ~x20 && x4 && x21 && x6 && ~x5 && ~x11 && ~x17 )
						nx_state = s1;
					else if( ~x64 && x19 && ~x20 && x4 && x21 && ~x6 && x5 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y15 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1347;
						end
					else if( ~x64 && x19 && ~x20 && x4 && x21 && ~x6 && ~x5 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x64 && x19 && ~x20 && x4 && x21 && ~x6 && ~x5 && ~x10 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x64 && x19 && ~x20 && x4 && x21 && ~x6 && ~x5 && ~x10 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x64 && x19 && ~x20 && x4 && x21 && ~x6 && ~x5 && ~x10 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x64 && x19 && ~x20 && x4 && x21 && ~x6 && ~x5 && ~x10 && ~x17 )
						nx_state = s1;
					else if( ~x64 && x19 && ~x20 && x4 && ~x21 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x64 && x19 && ~x20 && ~x4 && x21 && x6 && x5 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x64 && x19 && ~x20 && ~x4 && x21 && x6 && x5 && ~x13 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x64 && x19 && ~x20 && ~x4 && x21 && x6 && x5 && ~x13 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x64 && x19 && ~x20 && ~x4 && x21 && x6 && x5 && ~x13 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x64 && x19 && ~x20 && ~x4 && x21 && x6 && x5 && ~x13 && ~x17 )
						nx_state = s1;
					else if( ~x64 && x19 && ~x20 && ~x4 && x21 && x6 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x64 && x19 && ~x20 && ~x4 && x21 && ~x6 && x5 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x64 && x19 && ~x20 && ~x4 && x21 && ~x6 && x5 && ~x14 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x64 && x19 && ~x20 && ~x4 && x21 && ~x6 && x5 && ~x14 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x64 && x19 && ~x20 && ~x4 && x21 && ~x6 && x5 && ~x14 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x64 && x19 && ~x20 && ~x4 && x21 && ~x6 && x5 && ~x14 && ~x17 )
						nx_state = s1;
					else if( ~x64 && x19 && ~x20 && ~x4 && x21 && ~x6 && ~x5 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x64 && x19 && ~x20 && ~x4 && ~x21 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y23 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x64 && ~x19 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s1348;
						end
					else nx_state = s938;
				s939 : if( 1'b1 )
						begin
							y5 = 1'b1;	
							nx_state = s562;
						end
					else nx_state = s939;
				s940 : if( 1'b1 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else nx_state = s940;
				s941 : if( x26 && x28 && x23 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x26 && x28 && ~x23 && x25 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s941;
						end
					else if( x26 && x28 && ~x23 && ~x25 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( x26 && ~x28 && x3 && x25 )
						nx_state = s941;
					else if( x26 && ~x28 && x3 && ~x25 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( x26 && ~x28 && ~x3 && x4 && x5 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s942;
						end
					else if( x26 && ~x28 && ~x3 && x4 && ~x5 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( x26 && ~x28 && ~x3 && ~x4 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( ~x26 && x27 && x4 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s942;
						end
					else if( ~x26 && x27 && ~x4 )
						nx_state = s1;
					else if( ~x26 && ~x27 && x28 && x11 )
						nx_state = s1;
					else if( ~x26 && ~x27 && x28 && ~x11 )
						begin
							y13 = 1'b1;	
							nx_state = s897;
						end
					else if( ~x26 && ~x27 && ~x28 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s942;
						end
					else nx_state = s941;
				s942 : if( x26 && x28 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( x26 && x28 && ~x6 && x4 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s941;
						end
					else if( x26 && x28 && ~x6 && ~x4 )
						nx_state = s1;
					else if( x26 && ~x28 )
						nx_state = s1;
					else if( ~x26 && x28 && x27 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s614;
						end
					else if( ~x26 && x28 && ~x27 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s1349;
						end
					else if( ~x26 && ~x28 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s614;
						end
					else nx_state = s942;
				s943 : if( x26 && x28 && x9 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( x26 && x28 && ~x9 && x23 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s941;
						end
					else if( x26 && x28 && ~x9 && ~x23 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( x26 && ~x28 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( ~x26 && x27 && x1 && x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( ~x26 && x27 && x1 && ~x2 && x3 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s941;
						end
					else if( ~x26 && x27 && x1 && ~x2 && ~x3 )
						nx_state = s943;
					else if( ~x26 && x27 && ~x1 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( ~x26 && ~x27 && x1 && x5 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s613;
						end
					else if( ~x26 && ~x27 && x1 && x5 && ~x3 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x26 && ~x27 && x1 && x5 && ~x3 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s614;
						end
					else if( ~x26 && ~x27 && x1 && ~x5 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else if( ~x26 && ~x27 && ~x1 && x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( ~x26 && ~x27 && ~x1 && ~x2 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s941;
						end
					else nx_state = s943;
				s944 : if( x26 && x28 && x3 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s920;
						end
					else if( x26 && x28 && x3 && ~x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else if( x26 && x28 && ~x3 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else if( x26 && ~x28 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s917;
						end
					else if( ~x26 && x27 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x26 && ~x27 && x28 && x5 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( ~x26 && ~x27 && x28 && ~x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else if( ~x26 && ~x27 && ~x28 && x5 && x3 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s923;
						end
					else if( ~x26 && ~x27 && ~x28 && x5 && ~x3 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s924;
						end
					else if( ~x26 && ~x27 && ~x28 && x5 && ~x3 && ~x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s921;
						end
					else if( ~x26 && ~x27 && ~x28 && ~x5 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s917;
						end
					else nx_state = s944;
				s945 : if( x62 && x64 )
						begin
							y1 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s940;
						end
					else if( x62 && ~x64 && x66 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y37 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s1350;
						end
					else if( x62 && ~x64 && ~x66 && x6 && x3 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x62 && ~x64 && ~x66 && x6 && ~x3 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s18;
						end
					else if( x62 && ~x64 && ~x66 && x6 && ~x3 && ~x1 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s279;
						end
					else if( x62 && ~x64 && ~x66 && ~x6 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x62 && x30 )
						begin
							y47 = 1'b1;	y50 = 1'b1;	y61 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s1148;
						end
					else if( ~x62 && ~x30 && x31 )
						begin
							y47 = 1'b1;	y50 = 1'b1;	y61 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s1244;
						end
					else if( ~x62 && ~x30 && ~x31 )
						begin
							y33 = 1'b1;	
							nx_state = s589;
						end
					else nx_state = s945;
				s946 : if( 1'b1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							y8 = 1'b1;	
							nx_state = s1146;
						end
					else nx_state = s946;
				s947 : if( x63 && x11 )
						begin
							y14 = 1'b1;	y41 = 1'b1;	
							nx_state = s1351;
						end
					else if( x63 && ~x11 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s892;
						end
					else if( x63 && ~x11 && ~x15 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x63 && ~x11 && ~x15 && ~x18 )
						begin
							y44 = 1'b1;	y45 = 1'b1;	
							nx_state = s392;
						end
					else if( ~x63 )
						begin
							y25 = 1'b1;	
							nx_state = s1352;
						end
					else nx_state = s947;
				s948 : if( x63 )
						begin
							y9 = 1'b1;	y48 = 1'b1;	y49 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x63 )
						begin
							y6 = 1'b1;	
							nx_state = s659;
						end
					else nx_state = s948;
				s949 : if( x21 )
						begin
							y6 = 1'b1;	y17 = 1'b1;	y34 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s1211;
						end
					else if( ~x21 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x21 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x21 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x21 && ~x10 )
						nx_state = s1;
					else nx_state = s949;
				s950 : if( x64 && x62 )
						begin
							y1 = 1'b1;	y12 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1353;
						end
					else if( x64 && ~x62 && x21 )
						begin
							y4 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y93 = 1'b1;	
							nx_state = s516;
						end
					else if( x64 && ~x62 && ~x21 && x22 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y62 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s1189;
						end
					else if( x64 && ~x62 && ~x21 && ~x22 )
						begin
							y4 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y78 = 1'b1;	
							nx_state = s1354;
						end
					else if( ~x64 && x62 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s1355;
						end
					else if( ~x64 && ~x62 && x30 )
						begin
							y47 = 1'b1;	y56 = 1'b1;	y61 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s1110;
						end
					else if( ~x64 && ~x62 && ~x30 && x31 )
						begin
							y37 = 1'b1;	
							nx_state = s1356;
						end
					else if( ~x64 && ~x62 && ~x30 && ~x31 )
						begin
							y47 = 1'b1;	y50 = 1'b1;	y61 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s1148;
						end
					else nx_state = s950;
				s951 : if( x6 && x3 && x7 && x9 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x6 && x3 && x7 && ~x9 )
						begin
							y22 = 1'b1;	
							nx_state = s130;
						end
					else if( x6 && x3 && ~x7 && x8 && x9 && x11 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x6 && x3 && ~x7 && x8 && x9 && ~x11 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x6 && x3 && ~x7 && x8 && x9 && ~x11 && x14 && ~x10 )
						nx_state = s1;
					else if( x6 && x3 && ~x7 && x8 && x9 && ~x11 && ~x14 )
						nx_state = s1;
					else if( x6 && x3 && ~x7 && x8 && ~x9 && x10 )
						begin
							y7 = 1'b1;	
							nx_state = s109;
						end
					else if( x6 && x3 && ~x7 && x8 && ~x9 && ~x10 && x14 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x6 && x3 && ~x7 && x8 && ~x9 && ~x10 && x14 && ~x11 )
						nx_state = s1;
					else if( x6 && x3 && ~x7 && x8 && ~x9 && ~x10 && ~x14 )
						nx_state = s1;
					else if( x6 && x3 && ~x7 && ~x8 && x9 )
						begin
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s1357;
						end
					else if( x6 && x3 && ~x7 && ~x8 && ~x9 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s358;
						end
					else if( x6 && ~x3 && x8 && x9 && x15 && x16 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x6 && ~x3 && x8 && x9 && x15 && x16 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x6 && ~x3 && x8 && x9 && x15 && x16 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x6 && ~x3 && x8 && x9 && x15 && x16 && ~x14 )
						nx_state = s1;
					else if( x6 && ~x3 && x8 && x9 && x15 && ~x16 )
						begin
							y7 = 1'b1;	
							nx_state = s1358;
						end
					else if( x6 && ~x3 && x8 && x9 && ~x15 && x7 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x6 && ~x3 && x8 && x9 && ~x15 && ~x7 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	y31 = 1'b1;	
							nx_state = s1359;
						end
					else if( x6 && ~x3 && x8 && ~x9 && x15 && x17 )
						begin
							y7 = 1'b1;	
							nx_state = s1358;
						end
					else if( x6 && ~x3 && x8 && ~x9 && x15 && ~x17 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x6 && ~x3 && x8 && ~x9 && x15 && ~x17 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x6 && ~x3 && x8 && ~x9 && x15 && ~x17 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x6 && ~x3 && x8 && ~x9 && x15 && ~x17 && ~x14 )
						nx_state = s1;
					else if( x6 && ~x3 && x8 && ~x9 && ~x15 && x7 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x6 && ~x3 && x8 && ~x9 && ~x15 && ~x7 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s31;
						end
					else if( x6 && ~x3 && ~x8 && x9 && x15 && x18 )
						begin
							y7 = 1'b1;	
							nx_state = s1358;
						end
					else if( x6 && ~x3 && ~x8 && x9 && x15 && ~x18 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x6 && ~x3 && ~x8 && x9 && x15 && ~x18 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x6 && ~x3 && ~x8 && x9 && x15 && ~x18 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x6 && ~x3 && ~x8 && x9 && x15 && ~x18 && ~x14 )
						nx_state = s1;
					else if( x6 && ~x3 && ~x8 && x9 && ~x15 && x7 )
						begin
							y39 = 1'b1;	
							nx_state = s277;
						end
					else if( x6 && ~x3 && ~x8 && x9 && ~x15 && ~x7 )
						begin
							y25 = 1'b1;	
							nx_state = s1360;
						end
					else if( x6 && ~x3 && ~x8 && ~x9 && x15 && x18 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x6 && ~x3 && ~x8 && ~x9 && x15 && x18 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x6 && ~x3 && ~x8 && ~x9 && x15 && x18 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x6 && ~x3 && ~x8 && ~x9 && x15 && x18 && ~x14 )
						nx_state = s1;
					else if( x6 && ~x3 && ~x8 && ~x9 && x15 && ~x18 )
						begin
							y7 = 1'b1;	
							nx_state = s1358;
						end
					else if( x6 && ~x3 && ~x8 && ~x9 && ~x15 && x7 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x6 && ~x3 && ~x8 && ~x9 && ~x15 && ~x7 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x6 && x3 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s1361;
						end
					else if( ~x6 && ~x3 && x12 && x4 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s1362;
						end
					else if( ~x6 && ~x3 && x12 && ~x4 && x5 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s1363;
						end
					else if( ~x6 && ~x3 && x12 && ~x4 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y16 = 1'b1;	
							nx_state = s1359;
						end
					else if( ~x6 && ~x3 && ~x12 && x4 && x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y14 = 1'b1;	
							nx_state = s1359;
						end
					else if( ~x6 && ~x3 && ~x12 && x4 && ~x5 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s1364;
						end
					else if( ~x6 && ~x3 && ~x12 && ~x4 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s1365;
						end
					else nx_state = s951;
				s952 : if( x11 )
						begin
							y2 = 1'b1;	y22 = 1'b1;	
							nx_state = s952;
						end
					else if( ~x11 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else nx_state = s952;
				s953 : if( x62 && x20 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y8 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s1150;
						end
					else if( x62 && ~x20 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y15 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1192;
						end
					else if( ~x62 && x20 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							nx_state = s1213;
						end
					else if( ~x62 && ~x20 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							nx_state = s1366;
						end
					else nx_state = s953;
				s954 : if( 1'b1 )
						begin
							y26 = 1'b1;	
							nx_state = s262;
						end
					else nx_state = s954;
				s955 : if( x63 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x63 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x63 && x19 && ~x14 && ~x13 && x11 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( x63 && x19 && ~x14 && ~x13 && x11 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( x63 && x19 && ~x14 && ~x13 && ~x11 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( x63 && ~x19 )
						nx_state = s1;
					else if( ~x63 && x14 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x63 && x14 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x63 && x14 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x63 && x14 && ~x23 )
						nx_state = s1;
					else if( ~x63 && ~x14 )
						begin
							y39 = 1'b1;	
							nx_state = s1295;
						end
					else nx_state = s955;
				s956 : if( 1'b1 )
						begin
							y27 = 1'b1;	
							nx_state = s87;
						end
					else nx_state = s956;
				s957 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y70 = 1'b1;	
							y71 = 1'b1;	y72 = 1'b1;	
							nx_state = s1367;
						end
					else nx_state = s957;
				s958 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y70 = 1'b1;	
							y71 = 1'b1;	y72 = 1'b1;	
							nx_state = s1368;
						end
					else nx_state = s958;
				s959 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s1369;
						end
					else nx_state = s959;
				s960 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y61 = 1'b1;	
							y62 = 1'b1;	
							nx_state = s1370;
						end
					else nx_state = s960;
				s961 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y65 = 1'b1;	
							y66 = 1'b1;	
							nx_state = s1371;
						end
					else nx_state = s961;
				s962 : if( 1'b1 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else nx_state = s962;
				s963 : if( x62 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x62 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x62 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( x62 && ~x27 )
						nx_state = s1;
					else if( ~x62 && x64 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x62 && x64 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x62 && x64 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x62 && x64 && ~x11 )
						nx_state = s1;
					else if( ~x62 && ~x64 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( ~x62 && ~x64 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( ~x62 && ~x64 && x19 && ~x14 && ~x13 && x11 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( ~x62 && ~x64 && x19 && ~x14 && ~x13 && x11 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x62 && ~x64 && x19 && ~x14 && ~x13 && ~x11 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x62 && ~x64 && ~x19 )
						nx_state = s1;
					else nx_state = s963;
				s964 : if( 1'b1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s1372;
						end
					else nx_state = s964;
				s965 : if( x61 && x14 && x8 && x10 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s840;
						end
					else if( x61 && x14 && x8 && ~x10 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( x61 && x14 && ~x8 && x30 && x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s874;
						end
					else if( x61 && x14 && ~x8 && x30 && ~x1 && x4 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else if( x61 && x14 && ~x8 && x30 && ~x1 && ~x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s875;
						end
					else if( x61 && x14 && ~x8 && ~x30 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s840;
						end
					else if( x61 && ~x14 && x32 && x3 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s733;
						end
					else if( x61 && ~x14 && x32 && ~x3 )
						nx_state = s965;
					else if( x61 && ~x14 && ~x32 && x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s840;
						end
					else if( x61 && ~x14 && ~x32 && ~x3 )
						nx_state = s965;
					else if( ~x61 && x16 && x54 && x29 && x59 && x27 )
						begin
							y13 = 1'b1;	
							nx_state = s240;
						end
					else if( ~x61 && x16 && x54 && x29 && x59 && ~x27 )
						nx_state = s965;
					else if( ~x61 && x16 && x54 && x29 && ~x59 && x27 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( ~x61 && x16 && x54 && x29 && ~x59 && ~x27 )
						nx_state = s965;
					else if( ~x61 && x16 && x54 && ~x29 && x33 && x27 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( ~x61 && x16 && x54 && ~x29 && x33 && ~x27 )
						nx_state = s965;
					else if( ~x61 && x16 && x54 && ~x29 && ~x33 && x57 && x27 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( ~x61 && x16 && x54 && ~x29 && ~x33 && x57 && ~x27 )
						nx_state = s965;
					else if( ~x61 && x16 && x54 && ~x29 && ~x33 && ~x57 && x27 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( ~x61 && x16 && x54 && ~x29 && ~x33 && ~x57 && ~x27 )
						nx_state = s965;
					else if( ~x61 && x16 && ~x54 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( ~x61 && ~x16 && x37 && x56 && x1 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( ~x61 && ~x16 && x37 && x56 && ~x1 )
						nx_state = s965;
					else if( ~x61 && ~x16 && x37 && ~x56 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( ~x61 && ~x16 && ~x37 && x25 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	
							nx_state = s876;
						end
					else if( ~x61 && ~x16 && ~x37 && ~x25 && x5 && x4 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s320;
						end
					else if( ~x61 && ~x16 && ~x37 && ~x25 && x5 && ~x4 )
						nx_state = s965;
					else if( ~x61 && ~x16 && ~x37 && ~x25 && ~x5 && x4 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( ~x61 && ~x16 && ~x37 && ~x25 && ~x5 && ~x4 )
						nx_state = s965;
					else nx_state = s965;
				s966 : if( 1'b1 )
						begin
							y3 = 1'b1;	
							nx_state = s462;
						end
					else nx_state = s966;
				s967 : if( x62 && x33 && x32 && x10 && x11 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s470;
						end
					else if( x62 && x33 && x32 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s470;
						end
					else if( x62 && x33 && x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x62 && x33 && x32 && ~x10 )
						nx_state = s1;
					else if( x62 && x33 && ~x32 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s970;
						end
					else if( x62 && ~x33 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s970;
						end
					else if( ~x62 && x65 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x62 && x65 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x62 && x65 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x62 && x65 && ~x15 )
						nx_state = s1;
					else if( ~x62 && ~x65 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y56 = 1'b1;	
							nx_state = s1373;
						end
					else nx_state = s967;
				s968 : if( x33 && x32 && x10 && x11 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s470;
						end
					else if( x33 && x32 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s470;
						end
					else if( x33 && x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x33 && x32 && ~x10 )
						nx_state = s1;
					else if( x33 && ~x32 )
						begin
							y9 = 1'b1;	
							nx_state = s967;
						end
					else if( ~x33 )
						begin
							y9 = 1'b1;	
							nx_state = s967;
						end
					else nx_state = s968;
				s969 : if( x33 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s343;
						end
					else if( ~x33 && x32 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s343;
						end
					else if( ~x33 && ~x32 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x33 && ~x32 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x33 && ~x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x33 && ~x32 && ~x10 )
						nx_state = s1;
					else nx_state = s969;
				s970 : if( x33 && x32 && x10 && x11 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s470;
						end
					else if( x33 && x32 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s470;
						end
					else if( x33 && x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x33 && x32 && ~x10 )
						nx_state = s1;
					else if( x33 && ~x32 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s971;
						end
					else if( ~x33 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s971;
						end
					else nx_state = s970;
				s971 : if( x33 && x32 && x10 && x11 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s470;
						end
					else if( x33 && x32 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s470;
						end
					else if( x33 && x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x33 && x32 && ~x10 )
						nx_state = s1;
					else if( x33 && ~x32 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x33 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else nx_state = s971;
				s972 : if( x33 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s980;
						end
					else if( ~x33 && x32 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s980;
						end
					else if( ~x33 && ~x32 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x33 && ~x32 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x33 && ~x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x33 && ~x32 && ~x10 )
						nx_state = s1;
					else nx_state = s972;
				s973 : if( x32 )
						begin
							y31 = 1'b1;	y38 = 1'b1;	
							nx_state = s345;
						end
					else if( ~x32 && x33 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s977;
						end
					else if( ~x32 && ~x33 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x32 && ~x33 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x32 && ~x33 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x32 && ~x33 && ~x10 )
						nx_state = s1;
					else nx_state = s973;
				s974 : if( x32 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s345;
						end
					else if( ~x32 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s340;
						end
					else nx_state = s974;
				s975 : if( 1'b1 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s1374;
						end
					else nx_state = s975;
				s976 : if( x62 )
						begin
							y6 = 1'b1;	y47 = 1'b1;	
							nx_state = s1375;
						end
					else if( ~x62 && x63 )
						begin
							y26 = 1'b1;	
							nx_state = s262;
						end
					else if( ~x62 && ~x63 )
						begin
							y42 = 1'b1;	
							nx_state = s754;
						end
					else nx_state = s976;
				s977 : if( 1'b1 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s1376;
						end
					else nx_state = s977;
				s978 : if( 1'b1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1116;
						end
					else nx_state = s978;
				s979 : if( x32 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x32 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x32 && ~x10 )
						nx_state = s1;
					else if( ~x32 && x8 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s972;
						end
					else if( ~x32 && ~x8 && x33 )
						begin
							y53 = 1'b1;	
							nx_state = s1027;
						end
					else if( ~x32 && ~x8 && ~x33 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s972;
						end
					else nx_state = s979;
				s980 : if( 1'b1 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s352;
						end
					else nx_state = s980;
				s981 : if( 1'b1 )
						begin
							y4 = 1'b1;	y21 = 1'b1;	
							nx_state = s377;
						end
					else nx_state = s981;
				s982 : if( 1'b1 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else nx_state = s982;
				s983 : if( x14 )
						begin
							y26 = 1'b1;	
							nx_state = s1197;
						end
					else if( ~x14 && x7 )
						begin
							y25 = 1'b1;	
							nx_state = s238;
						end
					else if( ~x14 && ~x7 && x3 && x1 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x14 && ~x7 && x3 && x1 && ~x2 && x5 )
						nx_state = s983;
					else if( ~x14 && ~x7 && x3 && x1 && ~x2 && ~x5 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x14 && ~x7 && x3 && ~x1 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( ~x14 && ~x7 && ~x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else nx_state = s983;
				s984 : if( x11 )
						begin
							y18 = 1'b1;	y27 = 1'b1;	
							nx_state = s983;
						end
					else if( ~x11 )
						begin
							y10 = 1'b1;	y20 = 1'b1;	y26 = 1'b1;	
							nx_state = s984;
						end
					else nx_state = s984;
				s985 : if( x65 )
						begin
							y8 = 1'b1;	
							nx_state = s784;
						end
					else if( ~x65 )
						begin
							y7 = 1'b1;	
							nx_state = s891;
						end
					else nx_state = s985;
				s986 : if( x3 && x6 && x5 )
						nx_state = s1;
					else if( x3 && x6 && ~x5 && x8 && x7 && x10 && x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y17 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1379;
						end
					else if( x3 && x6 && ~x5 && x8 && x7 && x10 && ~x11 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1378;
						end
					else if( x3 && x6 && ~x5 && x8 && x7 && ~x10 )
						begin
							y72 = 1'b1;	
							nx_state = s1377;
						end
					else if( x3 && x6 && ~x5 && x8 && ~x7 && x9 && x18 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1378;
						end
					else if( x3 && x6 && ~x5 && x8 && ~x7 && x9 && ~x18 )
						nx_state = s1;
					else if( x3 && x6 && ~x5 && x8 && ~x7 && ~x9 && x17 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1378;
						end
					else if( x3 && x6 && ~x5 && x8 && ~x7 && ~x9 && ~x17 )
						nx_state = s1;
					else if( x3 && x6 && ~x5 && ~x8 && x9 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1378;
						end
					else if( x3 && x6 && ~x5 && ~x8 && ~x9 && x7 && x16 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1378;
						end
					else if( x3 && x6 && ~x5 && ~x8 && ~x9 && x7 && ~x16 )
						nx_state = s1;
					else if( x3 && x6 && ~x5 && ~x8 && ~x9 && ~x7 )
						begin
							y71 = 1'b1;	
							nx_state = s394;
						end
					else if( x3 && ~x6 && x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y17 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1379;
						end
					else if( x3 && ~x6 && ~x11 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1378;
						end
					else if( ~x3 && x4 )
						begin
							y14 = 1'b1;	
							nx_state = s124;
						end
					else if( ~x3 && ~x4 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s1380;
						end
					else nx_state = s986;
				s987 : if( 1'b1 )
						begin
							y22 = 1'b1;	
							nx_state = s1381;
						end
					else nx_state = s987;
				s988 : if( 1'b1 )
						begin
							y13 = 1'b1;	
							nx_state = s240;
						end
					else nx_state = s988;
				s989 : if( 1'b1 )
						begin
							y5 = 1'b1;	
							nx_state = s66;
						end
					else nx_state = s989;
				s990 : if( x17 )
						begin
							y3 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s1382;
						end
					else if( ~x17 )
						begin
							y5 = 1'b1;	y13 = 1'b1;	y17 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s990;
						end
					else nx_state = s990;
				s991 : if( x65 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	y21 = 1'b1;	
							nx_state = s1383;
						end
					else if( ~x65 && x20 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( ~x65 && ~x20 )
						begin
							y15 = 1'b1;	
							nx_state = s243;
						end
					else nx_state = s991;
				s992 : if( 1'b1 )
						begin
							y5 = 1'b1;	
							nx_state = s950;
						end
					else nx_state = s992;
				s993 : if( x61 )
						nx_state = s1;
					else if( ~x61 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	
							nx_state = s330;
						end
					else nx_state = s993;
				s994 : if( x69 )
						nx_state = s1;
					else if( ~x69 && x26 && x39 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( ~x69 && x26 && x39 && ~x32 && x14 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( ~x69 && x26 && x39 && ~x32 && ~x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x69 && x26 && ~x39 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s1124;
						end
					else if( ~x69 && ~x26 && x28 )
						nx_state = s1;
					else if( ~x69 && ~x26 && ~x28 && x6 && x38 && x5 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s922;
						end
					else if( ~x69 && ~x26 && ~x28 && x6 && x38 && x5 && ~x3 && x4 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s994;
						end
					else if( ~x69 && ~x26 && ~x28 && x6 && x38 && x5 && ~x3 && ~x4 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s995;
						end
					else if( ~x69 && ~x26 && ~x28 && x6 && x38 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x69 && ~x26 && ~x28 && x6 && ~x38 && x8 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s1185;
						end
					else if( ~x69 && ~x26 && ~x28 && x6 && ~x38 && ~x8 && x5 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s922;
						end
					else if( ~x69 && ~x26 && ~x28 && x6 && ~x38 && ~x8 && x5 && ~x3 && x4 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s994;
						end
					else if( ~x69 && ~x26 && ~x28 && x6 && ~x38 && ~x8 && x5 && ~x3 && ~x4 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s995;
						end
					else if( ~x69 && ~x26 && ~x28 && x6 && ~x38 && ~x8 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x69 && ~x26 && ~x28 && ~x6 && x24 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s1185;
						end
					else if( ~x69 && ~x26 && ~x28 && ~x6 && ~x24 )
						nx_state = s1;
					else nx_state = s994;
				s995 : if( x69 )
						nx_state = s1;
					else if( ~x69 && x26 && x21 )
						nx_state = s1;
					else if( ~x69 && x26 && ~x21 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else if( ~x69 && ~x26 && x27 )
						nx_state = s1;
					else if( ~x69 && ~x26 && ~x27 && x28 && x34 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( ~x69 && ~x26 && ~x27 && x28 && ~x34 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s922;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && x19 && x24 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s1185;
						end
					else if( ~x69 && ~x26 && ~x27 && ~x28 && x19 && ~x24 )
						nx_state = s1;
					else if( ~x69 && ~x26 && ~x27 && ~x28 && ~x19 )
						begin
							y27 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s1124;
						end
					else nx_state = s995;
				s996 : if( x46 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s697;
						end
					else if( ~x46 && x34 && x2 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s691;
						end
					else if( ~x46 && x34 && ~x2 )
						nx_state = s996;
					else if( ~x46 && ~x34 && x35 && x2 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s997;
						end
					else if( ~x46 && ~x34 && x35 && ~x2 )
						nx_state = s996;
					else if( ~x46 && ~x34 && ~x35 && x2 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s998;
						end
					else if( ~x46 && ~x34 && ~x35 && ~x2 )
						nx_state = s996;
					else nx_state = s996;
				s997 : if( x63 && x46 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( x63 && ~x46 && x37 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( x63 && ~x46 && ~x37 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s697;
						end
					else if( ~x63 && x15 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( ~x63 && ~x15 && x6 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x63 && ~x15 && ~x6 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s705;
						end
					else nx_state = s997;
				s998 : if( x15 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s996;
						end
					else if( ~x15 && x36 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( ~x15 && ~x36 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s996;
						end
					else nx_state = s998;
				s999 : if( x15 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( ~x15 && x6 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x15 && ~x6 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s705;
						end
					else nx_state = s999;
				s1000 : if( x15 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s477;
						end
					else if( ~x15 && x5 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( ~x15 && ~x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s477;
						end
					else nx_state = s1000;
				s1001 : if( x16 && x22 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x16 && ~x22 && x23 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( x16 && ~x22 && ~x23 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x16 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s604;
						end
					else nx_state = s1001;
				s1002 : if( 1'b1 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s251;
						end
					else nx_state = s1002;
				s1003 : if( x21 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s810;
						end
					else if( x21 && ~x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( ~x21 && x19 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else if( ~x21 && ~x19 && x22 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else if( ~x21 && ~x19 && ~x22 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s810;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else nx_state = s1003;
				s1004 : if( x21 && x18 && x16 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else if( x21 && x18 && ~x16 && x17 && x13 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else if( x21 && x18 && ~x16 && x17 && ~x13 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x21 && x18 && ~x16 && x17 && ~x13 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x21 && x18 && ~x16 && x17 && ~x13 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x21 && x18 && ~x16 && x17 && ~x13 && ~x4 )
						nx_state = s1;
					else if( x21 && x18 && ~x16 && ~x17 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else if( x21 && ~x18 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x21 && ~x18 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x21 && ~x18 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x21 && ~x18 && ~x4 )
						nx_state = s1;
					else if( ~x21 && x19 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x21 && ~x19 && x22 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x21 && ~x19 && ~x22 && x20 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && ~x19 && ~x22 && x20 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && ~x19 && ~x22 && x20 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x19 && ~x22 && x20 && ~x4 )
						nx_state = s1;
					else if( ~x21 && ~x19 && ~x22 && ~x20 && x16 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && x13 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && ~x13 && x17 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && ~x13 && x17 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && ~x13 && x17 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && ~x13 && x17 && ~x4 )
						nx_state = s1;
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && ~x13 && ~x17 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s1004;
				s1005 : if( 1'b1 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else nx_state = s1005;
				s1006 : if( 1'b1 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s1008;
						end
					else nx_state = s1006;
				s1007 : if( x65 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x65 )
						begin
							y51 = 1'b1;	
							nx_state = s655;
						end
					else nx_state = s1007;
				s1008 : if( 1'b1 )
						begin
							y2 = 1'b1;	y15 = 1'b1;	y31 = 1'b1;	
							nx_state = s1384;
						end
					else nx_state = s1008;
				s1009 : if( x63 && x17 )
						begin
							y13 = 1'b1;	
							nx_state = s763;
						end
					else if( x63 && ~x17 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x63 && ~x17 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x63 && ~x17 && x19 && ~x14 && ~x13 && x11 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( x63 && ~x17 && x19 && ~x14 && ~x13 && x11 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( x63 && ~x17 && x19 && ~x14 && ~x13 && ~x11 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( x63 && ~x17 && ~x19 )
						nx_state = s1;
					else if( ~x63 && x64 && x67 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x63 && x64 && x67 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x63 && x64 && x67 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( ~x63 && x64 && x67 && ~x14 )
						nx_state = s1;
					else if( ~x63 && x64 && ~x67 )
						begin
							y54 = 1'b1;	
							nx_state = s281;
						end
					else if( ~x63 && ~x64 )
						begin
							y38 = 1'b1;	
							nx_state = s845;
						end
					else nx_state = s1009;
				s1010 : if( x64 && x19 )
						begin
							y7 = 1'b1;	
							nx_state = s1385;
						end
					else if( x64 && ~x19 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x64 && ~x19 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x64 && ~x19 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x64 && ~x19 && ~x18 )
						nx_state = s1;
					else if( ~x64 && x14 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x64 && x14 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x64 && x14 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x64 && x14 && ~x23 )
						nx_state = s1;
					else if( ~x64 && ~x14 )
						begin
							y40 = 1'b1;	
							nx_state = s751;
						end
					else nx_state = s1010;
				s1011 : if( x17 )
						begin
							y24 = 1'b1;	
							nx_state = s1012;
						end
					else if( ~x17 )
						begin
							y5 = 1'b1;	y13 = 1'b1;	y17 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1011;
						end
					else nx_state = s1011;
				s1012 : if( x64 && x66 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y16 = 1'b1;	y27 = 1'b1;	
							nx_state = s1386;
						end
					else if( x64 && ~x66 )
						begin
							y2 = 1'b1;	y15 = 1'b1;	y31 = 1'b1;	
							nx_state = s1387;
						end
					else if( ~x64 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else nx_state = s1012;
				s1013 : if( x11 )
						begin
							y1 = 1'b1;	y22 = 1'b1;	
							nx_state = s1013;
						end
					else if( ~x11 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s8;
						end
					else nx_state = s1013;
				s1014 : if( 1'b1 )
						begin
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s1357;
						end
					else nx_state = s1014;
				s1015 : if( 1'b1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y20 = 1'b1;	
							y40 = 1'b1;	y42 = 1'b1;	
							nx_state = s1388;
						end
					else nx_state = s1015;
				s1016 : if( 1'b1 )
						begin
							y15 = 1'b1;	y20 = 1'b1;	
							nx_state = s665;
						end
					else nx_state = s1016;
				s1017 : if( x63 && x64 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s1389;
						end
					else if( x63 && ~x64 && x9 )
						begin
							y23 = 1'b1;	
							nx_state = s588;
						end
					else if( x63 && ~x64 && ~x9 )
						nx_state = s1017;
					else if( ~x63 )
						begin
							y27 = 1'b1;	
							nx_state = s648;
						end
					else nx_state = s1017;
				s1018 : if( 1'b1 )
						begin
							y13 = 1'b1;	
							nx_state = s769;
						end
					else nx_state = s1018;
				s1019 : if( x49 && x50 )
						begin
							y29 = 1'b1;	
							nx_state = s771;
						end
					else if( x49 && ~x50 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y37 = 1'b1;	
							y39 = 1'b1;	y44 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x49 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y35 = 1'b1;	
							y37 = 1'b1;	y39 = 1'b1;	
							nx_state = s584;
						end
					else nx_state = s1019;
				s1020 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s48;
						end
					else nx_state = s1020;
				s1021 : if( x17 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y18 = 1'b1;	
							nx_state = s1390;
						end
					else if( ~x17 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y13 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1021;
						end
					else nx_state = s1021;
				s1022 : if( x14 && x65 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x14 && x65 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x14 && x65 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x14 && ~x65 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x14 && ~x65 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x14 && ~x65 && ~x15 && ~x16 )
						nx_state = s1;
					else if( ~x14 )
						nx_state = s1;
					else nx_state = s1022;
				s1023 : if( x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x14 )
						nx_state = s1;
					else nx_state = s1023;
				s1024 : if( x63 )
						nx_state = s1;
					else if( ~x63 && x14 && x10 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x63 && x14 && ~x10 && x11 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x63 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x63 && ~x14 )
						nx_state = s1;
					else nx_state = s1024;
				s1025 : if( x63 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s1391;
						end
					else if( ~x63 )
						begin
							y5 = 1'b1;	
							nx_state = s937;
						end
					else nx_state = s1025;
				s1026 : if( x21 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s791;
						end
					else if( x21 && ~x3 )
						begin
							y4 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y93 = 1'b1;	
							nx_state = s1301;
						end
					else if( ~x21 && x22 && x3 )
						begin
							y62 = 1'b1;	y65 = 1'b1;	y78 = 1'b1;	
							y96 = 1'b1;	
							nx_state = s1392;
						end
					else if( ~x21 && x22 && ~x3 )
						begin
							y60 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y79 = 1'b1;	
							nx_state = s1392;
						end
					else if( ~x21 && ~x22 && x3 )
						begin
							y62 = 1'b1;	y65 = 1'b1;	y78 = 1'b1;	
							y96 = 1'b1;	
							nx_state = s1393;
						end
					else if( ~x21 && ~x22 && ~x3 )
						begin
							y60 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y79 = 1'b1;	
							nx_state = s1393;
						end
					else nx_state = s1026;
				s1027 : if( x62 && x33 )
						begin
							y6 = 1'b1;	y35 = 1'b1;	y40 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s355;
						end
					else if( x62 && ~x33 && x32 )
						begin
							y6 = 1'b1;	y35 = 1'b1;	y40 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s355;
						end
					else if( x62 && ~x33 && ~x32 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x62 && ~x33 && ~x32 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x62 && ~x33 && ~x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x62 && ~x33 && ~x32 && ~x10 )
						nx_state = s1;
					else if( ~x62 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x62 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x62 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x62 && ~x18 )
						nx_state = s1;
					else nx_state = s1027;
				s1028 : if( x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x10 )
						nx_state = s1;
					else nx_state = s1028;
				s1029 : if( 1'b1 )
						begin
							y6 = 1'b1;	y25 = 1'b1;	y31 = 1'b1;	
							y32 = 1'b1;	y45 = 1'b1;	
							nx_state = s1394;
						end
					else nx_state = s1029;
				s1030 : if( x62 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x62 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x62 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( x62 && ~x21 )
						nx_state = s1;
					else if( ~x62 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x62 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x62 && ~x9 )
						nx_state = s1;
					else nx_state = s1030;
				s1031 : if( 1'b1 )
						begin
							y35 = 1'b1;	
							nx_state = s718;
						end
					else nx_state = s1031;
				s1032 : if( 1'b1 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else nx_state = s1032;
				s1033 : if( x64 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( ~x64 && x66 && x4 )
						begin
							y29 = 1'b1;	y47 = 1'b1;	y49 = 1'b1;	
							y58 = 1'b1;	y61 = 1'b1;	y67 = 1'b1;	
							nx_state = s1395;
						end
					else if( ~x64 && x66 && ~x4 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x64 && ~x66 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y69 = 1'b1;	
							y70 = 1'b1;	y71 = 1'b1;	
							nx_state = s1396;
						end
					else nx_state = s1033;
				s1034 : if( x21 && x20 && x12 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x21 && x20 && x12 && ~x8 && x7 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x21 && x20 && x12 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x21 && x20 && ~x12 )
						nx_state = s1;
					else if( x21 && ~x20 && x6 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x21 && ~x20 && x6 && ~x7 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else if( x21 && ~x20 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x21 && ~x20 && ~x6 )
						nx_state = s1;
					else if( ~x21 )
						nx_state = s1;
					else nx_state = s1034;
				s1035 : if( x63 && x15 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s9;
						end
					else if( x63 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x63 && ~x15 && x16 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x63 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s299;
						end
					else if( ~x63 )
						nx_state = s1;
					else nx_state = s1035;
				s1036 : if( 1'b1 )
						begin
							y3 = 1'b1;	y17 = 1'b1;	y27 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s1397;
						end
					else nx_state = s1036;
				s1037 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1398;
						end
					else nx_state = s1037;
				s1038 : if( x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( x19 && ~x14 && ~x13 )
						nx_state = s1038;
					else if( ~x19 )
						nx_state = s1;
					else nx_state = s1038;
				s1039 : if( x66 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x66 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else nx_state = s1039;
				s1040 : if( 1'b1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s730;
						end
					else nx_state = s1040;
				s1041 : if( 1'b1 )
						begin
							y10 = 1'b1;	
							nx_state = s193;
						end
					else nx_state = s1041;
				s1042 : if( x63 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y44 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1399;
						end
					else if( ~x63 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y53 = 1'b1;	
							nx_state = s1400;
						end
					else nx_state = s1042;
				s1043 : if( x26 )
						begin
							y74 = 1'b1;	
							nx_state = s847;
						end
					else if( ~x26 && x27 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( ~x26 && ~x27 )
						begin
							y69 = 1'b1;	y73 = 1'b1;	
							nx_state = s1043;
						end
					else nx_state = s1043;
				s1044 : if( 1'b1 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	
							nx_state = s895;
						end
					else nx_state = s1044;
				s1045 : if( x16 && x15 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( x16 && ~x15 && x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s326;
						end
					else if( x16 && ~x15 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s929;
						end
					else if( ~x16 && x15 && x11 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x16 && x15 && ~x11 && x10 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s455;
						end
					else if( ~x16 && x15 && ~x11 && ~x10 )
						nx_state = s1045;
					else if( ~x16 && ~x15 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else nx_state = s1045;
				s1046 : if( 1'b1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s1249;
						end
					else nx_state = s1046;
				s1047 : if( 1'b1 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s140;
						end
					else nx_state = s1047;
				s1048 : if( x66 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s1401;
						end
					else if( ~x66 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s1249;
						end
					else nx_state = s1048;
				s1049 : if( x63 && x16 && x22 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x63 && x16 && ~x22 && x23 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( x63 && x16 && ~x22 && ~x23 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x63 && ~x16 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s604;
						end
					else if( ~x63 && x64 )
						begin
							y7 = 1'b1;	
							nx_state = s1385;
						end
					else if( ~x63 && ~x64 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s1402;
						end
					else nx_state = s1049;
				s1050 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s1046;
						end
					else nx_state = s1050;
				s1051 : if( x63 && x17 && x16 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x63 && x17 && x16 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x63 && x17 && x16 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x63 && x17 && ~x16 )
						nx_state = s1;
					else if( x63 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s1403;
						end
					else if( ~x63 && x65 && x3 && x6 && x5 && x9 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x63 && x65 && x3 && x6 && x5 && x9 && ~x7 && x8 && x17 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( ~x63 && x65 && x3 && x6 && x5 && x9 && ~x7 && x8 && ~x17 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x65 && x3 && x6 && x5 && x9 && ~x7 && x8 && ~x17 && x15 && ~x16 )
						nx_state = s1;
					else if( ~x63 && x65 && x3 && x6 && x5 && x9 && ~x7 && x8 && ~x17 && ~x15 )
						nx_state = s1;
					else if( ~x63 && x65 && x3 && x6 && x5 && x9 && ~x7 && ~x8 )
						begin
							y5 = 1'b1;	y31 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1400;
						end
					else if( ~x63 && x65 && x3 && x6 && x5 && ~x9 && x7 )
						begin
							y68 = 1'b1;	
							nx_state = s1404;
						end
					else if( ~x63 && x65 && x3 && x6 && x5 && ~x9 && ~x7 && x8 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( ~x63 && x65 && x3 && x6 && x5 && ~x9 && ~x7 && x8 && ~x18 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x65 && x3 && x6 && x5 && ~x9 && ~x7 && x8 && ~x18 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x65 && x3 && x6 && x5 && ~x9 && ~x7 && x8 && ~x18 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x63 && x65 && x3 && x6 && x5 && ~x9 && ~x7 && x8 && ~x18 && ~x15 )
						nx_state = s1;
					else if( ~x63 && x65 && x3 && x6 && x5 && ~x9 && ~x7 && ~x8 )
						begin
							y5 = 1'b1;	y34 = 1'b1;	y35 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1405;
						end
					else if( ~x63 && x65 && x3 && x6 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1406;
						end
					else if( ~x63 && x65 && x3 && ~x6 && x5 && x8 && x7 && x9 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x63 && x65 && x3 && ~x6 && x5 && x8 && x7 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( ~x63 && x65 && x3 && ~x6 && x5 && x8 && ~x7 && x11 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s1407;
						end
					else if( ~x63 && x65 && x3 && ~x6 && x5 && x8 && ~x7 && x11 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y28 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s1400;
						end
					else if( ~x63 && x65 && x3 && ~x6 && x5 && x8 && ~x7 && ~x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1408;
						end
					else if( ~x63 && x65 && x3 && ~x6 && x5 && ~x8 && x9 && x7 )
						begin
							y17 = 1'b1;	
							nx_state = s98;
						end
					else if( ~x63 && x65 && x3 && ~x6 && x5 && ~x8 && x9 && ~x7 && x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1400;
						end
					else if( ~x63 && x65 && x3 && ~x6 && x5 && ~x8 && x9 && ~x7 && ~x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1408;
						end
					else if( ~x63 && x65 && x3 && ~x6 && x5 && ~x8 && ~x9 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x63 && x65 && x3 && ~x6 && x5 && ~x8 && ~x9 && ~x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y22 = 1'b1;	
							nx_state = s1400;
						end
					else if( ~x63 && x65 && x3 && ~x6 && ~x5 && x11 && x8 && x9 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y47 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s1409;
						end
					else if( ~x63 && x65 && x3 && ~x6 && ~x5 && x11 && x8 && x9 && ~x7 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1400;
						end
					else if( ~x63 && x65 && x3 && ~x6 && ~x5 && x11 && x8 && ~x9 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y47 = 1'b1;	
							y58 = 1'b1;	
							nx_state = s1410;
						end
					else if( ~x63 && x65 && x3 && ~x6 && ~x5 && x11 && x8 && ~x9 && ~x7 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	y14 = 1'b1;	
							y20 = 1'b1;	y22 = 1'b1;	
							nx_state = s1400;
						end
					else if( ~x63 && x65 && x3 && ~x6 && ~x5 && x11 && ~x8 && x7 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y50 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s1411;
						end
					else if( ~x63 && x65 && x3 && ~x6 && ~x5 && x11 && ~x8 && x7 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y40 = 1'b1;	
							y59 = 1'b1;	
							nx_state = s1412;
						end
					else if( ~x63 && x65 && x3 && ~x6 && ~x5 && x11 && ~x8 && ~x7 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	y22 = 1'b1;	
							nx_state = s1400;
						end
					else if( ~x63 && x65 && x3 && ~x6 && ~x5 && ~x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1413;
						end
					else if( ~x63 && x65 && ~x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s1414;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && x20 && x4 && x6 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && x20 && x4 && ~x6 )
						begin
							y38 = 1'b1;	
							nx_state = s845;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && x20 && ~x4 && x5 && x6 && x9 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && x20 && ~x4 && x5 && x6 && ~x9 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && x20 && ~x4 && x5 && x6 && ~x9 && x17 && ~x8 )
						nx_state = s1;
					else if( ~x63 && ~x65 && x67 && x15 && x21 && x20 && ~x4 && x5 && x6 && ~x9 && ~x17 )
						nx_state = s1;
					else if( ~x63 && ~x65 && x67 && x15 && x21 && x20 && ~x4 && x5 && ~x6 && x8 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && x20 && ~x4 && x5 && ~x6 && ~x8 && x17 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && x20 && ~x4 && x5 && ~x6 && ~x8 && x17 && ~x9 )
						nx_state = s1;
					else if( ~x63 && ~x65 && x67 && x15 && x21 && x20 && ~x4 && x5 && ~x6 && ~x8 && ~x17 )
						nx_state = s1;
					else if( ~x63 && ~x65 && x67 && x15 && x21 && x20 && ~x4 && ~x5 && x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y39 = 1'b1;	y41 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && x20 && ~x4 && ~x5 && ~x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y13 = 1'b1;	
							y40 = 1'b1;	y42 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && x5 && x6 && x4 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s1270;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && x5 && x6 && ~x4 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && x5 && x6 && ~x4 && ~x13 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && x5 && x6 && ~x4 && ~x13 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && x5 && x6 && ~x4 && ~x13 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && x5 && x6 && ~x4 && ~x13 && ~x17 )
						nx_state = s1;
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && x5 && ~x6 && x4 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y15 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1347;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && x5 && ~x6 && ~x4 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && x5 && ~x6 && ~x4 && ~x14 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && x5 && ~x6 && ~x4 && ~x14 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && x5 && ~x6 && ~x4 && ~x14 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && x5 && ~x6 && ~x4 && ~x14 && ~x17 )
						nx_state = s1;
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && ~x5 && x6 && x4 && x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && ~x5 && x6 && x4 && ~x11 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && ~x5 && x6 && x4 && ~x11 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && ~x5 && x6 && x4 && ~x11 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && ~x5 && x6 && x4 && ~x11 && ~x17 )
						nx_state = s1;
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && ~x5 && x6 && ~x4 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && ~x5 && ~x6 && x4 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && ~x5 && ~x6 && x4 && ~x10 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && ~x5 && ~x6 && x4 && ~x10 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && ~x5 && ~x6 && x4 && ~x10 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && ~x5 && ~x6 && x4 && ~x10 && ~x17 )
						nx_state = s1;
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && x18 && ~x5 && ~x6 && ~x4 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x63 && ~x65 && x67 && x15 && x21 && ~x20 && ~x18 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s1415;
						end
					else if( ~x63 && ~x65 && x67 && x15 && ~x21 && x18 && x20 && x5 && x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x63 && ~x65 && x67 && x15 && ~x21 && x18 && x20 && x5 && ~x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1406;
						end
					else if( ~x63 && ~x65 && x67 && x15 && ~x21 && x18 && x20 && ~x5 )
						begin
							y3 = 1'b1;	y10 = 1'b1;	y30 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s1416;
						end
					else if( ~x63 && ~x65 && x67 && x15 && ~x21 && x18 && ~x20 && x4 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	y24 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x63 && ~x65 && x67 && x15 && ~x21 && x18 && ~x20 && ~x4 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	y23 = 1'b1;	
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x63 && ~x65 && x67 && x15 && ~x21 && ~x18 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s1415;
						end
					else if( ~x63 && ~x65 && x67 && ~x15 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s678;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && x5 && x21 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y13 = 1'b1;	
							y31 = 1'b1;	y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s1417;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && x5 && x21 && ~x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y13 = 1'b1;	
							y34 = 1'b1;	y36 = 1'b1;	
							nx_state = s1417;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && x5 && ~x21 && x22 && x10 && x24 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && x5 && ~x21 && x22 && x10 && ~x24 && x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && x5 && ~x21 && x22 && x10 && ~x24 && x26 && ~x25 )
						nx_state = s1;
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && x5 && ~x21 && x22 && x10 && ~x24 && ~x26 )
						nx_state = s1;
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && x5 && ~x21 && x22 && ~x10 && x25 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && x5 && ~x21 && x22 && ~x10 && ~x25 && x26 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && x5 && ~x21 && x22 && ~x10 && ~x25 && x26 && ~x24 )
						nx_state = s1;
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && x5 && ~x21 && x22 && ~x10 && ~x25 && ~x26 )
						nx_state = s1;
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && x5 && ~x21 && ~x22 && x23 && x10 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && x5 && ~x21 && ~x22 && x23 && ~x10 )
						begin
							y22 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && x5 && ~x21 && ~x22 && ~x23 && x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && x5 && ~x21 && ~x22 && ~x23 && x26 && ~x25 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && x5 && ~x21 && ~x22 && ~x23 && x26 && ~x25 && ~x24 )
						nx_state = s1;
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && x5 && ~x21 && ~x22 && ~x23 && ~x26 )
						nx_state = s1;
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && x9 && x8 && x14 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && x9 && x8 && ~x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s743;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && x9 && ~x8 && x10 && x11 && x14 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && x9 && ~x8 && x10 && x11 && ~x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s743;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && x9 && ~x8 && x10 && ~x11 && x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && x9 && ~x8 && x10 && ~x11 && x26 && ~x25 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && x9 && ~x8 && x10 && ~x11 && x26 && ~x25 && ~x24 )
						nx_state = s1;
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && x9 && ~x8 && x10 && ~x11 && ~x26 )
						nx_state = s1;
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && x9 && ~x8 && ~x10 && x12 && x14 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && x9 && ~x8 && ~x10 && x12 && ~x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s743;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && x9 && ~x8 && ~x10 && ~x12 && x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && x9 && ~x8 && ~x10 && ~x12 && x26 && ~x25 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && x9 && ~x8 && ~x10 && ~x12 && x26 && ~x25 && ~x24 )
						nx_state = s1;
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && x9 && ~x8 && ~x10 && ~x12 && ~x26 )
						nx_state = s1;
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && ~x9 && x10 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s1418;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && ~x9 && x10 && ~x8 && x14 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && ~x9 && x10 && ~x8 && ~x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s743;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && ~x9 && ~x10 && x8 && x13 && x14 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && ~x9 && ~x10 && x8 && x13 && ~x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s743;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && ~x9 && ~x10 && x8 && ~x13 && x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && ~x9 && ~x10 && x8 && ~x13 && x26 && ~x25 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && ~x9 && ~x10 && x8 && ~x13 && x26 && ~x25 && ~x24 )
						nx_state = s1;
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && ~x9 && ~x10 && x8 && ~x13 && ~x26 )
						nx_state = s1;
					else if( ~x63 && ~x65 && ~x67 && x3 && x6 && ~x5 && ~x9 && ~x10 && ~x8 )
						begin
							y30 = 1'b1;	
							nx_state = s291;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && ~x6 && x5 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y26 = 1'b1;	
							y37 = 1'b1;	y38 = 1'b1;	
							nx_state = s1417;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && ~x6 && x5 && ~x7 && x8 )
						begin
							y5 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s1417;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && ~x6 && x5 && ~x7 && ~x8 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s1417;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && ~x6 && x5 && ~x7 && ~x8 && ~x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s743;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && ~x6 && ~x5 && x8 )
						begin
							y5 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s1417;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && ~x6 && ~x5 && ~x8 && x14 )
						begin
							y25 = 1'b1;	y26 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s1417;
						end
					else if( ~x63 && ~x65 && ~x67 && x3 && ~x6 && ~x5 && ~x8 && ~x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s743;
						end
					else if( ~x63 && ~x65 && ~x67 && ~x3 )
						begin
							y5 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s1419;
						end
					else nx_state = s1051;
				s1052 : if( 1'b1 )
						begin
							y9 = 1'b1;	
							nx_state = s1420;
						end
					else nx_state = s1052;
				s1053 : if( x64 )
						begin
							y6 = 1'b1;	
							nx_state = s431;
						end
					else if( ~x64 && x30 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x64 && ~x30 )
						begin
							y5 = 1'b1;	
							nx_state = s937;
						end
					else nx_state = s1053;
				s1054 : if( 1'b1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y48 = 1'b1;	y50 = 1'b1;	
							nx_state = s1421;
						end
					else nx_state = s1054;
				s1055 : if( x33 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s350;
						end
					else if( ~x33 && x32 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s350;
						end
					else if( ~x33 && ~x32 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x33 && ~x32 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x33 && ~x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x33 && ~x32 && ~x10 )
						nx_state = s1;
					else nx_state = s1055;
				s1056 : if( 1'b1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s354;
						end
					else nx_state = s1056;
				s1057 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y33 = 1'b1;	
							y59 = 1'b1;	y60 = 1'b1;	y61 = 1'b1;	
							y62 = 1'b1;	
							nx_state = s1422;
						end
					else nx_state = s1057;
				s1058 : if( 1'b1 )
						begin
							y42 = 1'b1;	
							nx_state = s1423;
						end
					else nx_state = s1058;
				s1059 : if( x32 )
						begin
							y53 = 1'b1;	
							nx_state = s1424;
						end
					else if( ~x32 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y35 = 1'b1;	y40 = 1'b1;	
							nx_state = s351;
						end
					else nx_state = s1059;
				s1060 : if( 1'b1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	y40 = 1'b1;	
							nx_state = s1425;
						end
					else nx_state = s1060;
				s1061 : if( x32 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y27 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s339;
						end
					else if( ~x32 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x32 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x32 && ~x10 )
						nx_state = s1;
					else nx_state = s1061;
				s1062 : if( 1'b1 )
						begin
							y53 = 1'b1;	
							nx_state = s1027;
						end
					else nx_state = s1062;
				s1063 : if( x32 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x32 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x32 && ~x10 )
						nx_state = s1;
					else if( ~x32 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1327;
						end
					else nx_state = s1063;
				s1064 : if( 1'b1 )
						begin
							y8 = 1'b1;	y15 = 1'b1;	y19 = 1'b1;	
							nx_state = s1426;
						end
					else nx_state = s1064;
				s1065 : if( x16 )
						begin
							y6 = 1'b1;	y40 = 1'b1;	y41 = 1'b1;	
							y42 = 1'b1;	y50 = 1'b1;	
							nx_state = s1028;
						end
					else if( ~x16 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x16 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x16 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x16 && ~x10 )
						nx_state = s1;
					else nx_state = s1065;
				s1066 : if( 1'b1 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							nx_state = s1210;
						end
					else nx_state = s1066;
				s1067 : if( x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s609;
						end
					else if( ~x3 && x19 )
						begin
							y14 = 1'b1;	
							nx_state = s366;
						end
					else if( ~x3 && ~x19 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else nx_state = s1067;
				s1068 : if( 1'b1 )
						begin
							y28 = 1'b1;	
							nx_state = s1427;
						end
					else nx_state = s1068;
				s1069 : if( 1'b1 )
						begin
							y46 = 1'b1;	
							nx_state = s1428;
						end
					else nx_state = s1069;
				s1070 : if( x20 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s890;
						end
					else if( ~x20 )
						nx_state = s1;
					else nx_state = s1070;
				s1071 : if( x62 )
						begin
							y9 = 1'b1;	
							nx_state = s1429;
						end
					else if( ~x62 && x11 )
						begin
							y50 = 1'b1;	
							nx_state = s658;
						end
					else if( ~x62 && ~x11 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else nx_state = s1071;
				s1072 : if( x64 )
						begin
							y6 = 1'b1;	
							nx_state = s368;
						end
					else if( ~x64 )
						begin
							y42 = 1'b1;	
							nx_state = s754;
						end
					else nx_state = s1072;
				s1073 : if( 1'b1 )
						begin
							y6 = 1'b1;	
							nx_state = s368;
						end
					else nx_state = s1073;
				s1074 : if( 1'b1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1430;
						end
					else nx_state = s1074;
				s1075 : if( 1'b1 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else nx_state = s1075;
				s1076 : if( x27 )
						begin
							y21 = 1'b1;	
							nx_state = s317;
						end
					else if( ~x27 )
						begin
							y69 = 1'b1;	y73 = 1'b1;	
							nx_state = s1043;
						end
					else nx_state = s1076;
				s1077 : if( 1'b1 )
						begin
							y2 = 1'b1;	y37 = 1'b1;	y39 = 1'b1;	
							nx_state = s1144;
						end
					else nx_state = s1077;
				s1078 : if( x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x8 )
						nx_state = s1;
					else nx_state = s1078;
				s1079 : if( 1'b1 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s1182;
						end
					else nx_state = s1079;
				s1080 : if( 1'b1 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s131;
						end
					else nx_state = s1080;
				s1081 : if( x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							y18 = 1'b1;	y29 = 1'b1;	
							nx_state = s1001;
						end
					else if( ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1002;
						end
					else nx_state = s1081;
				s1082 : if( 1'b1 )
						begin
							y5 = 1'b1;	
							nx_state = s791;
						end
					else nx_state = s1082;
				s1083 : if( x63 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s1431;
						end
					else if( ~x63 && x64 && x21 && x10 )
						begin
							y5 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x63 && x64 && x21 && ~x10 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x63 && x64 && x21 && ~x10 && ~x12 && x17 && x16 && x19 && x11 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x63 && x64 && x21 && ~x10 && ~x12 && x17 && x16 && x19 && ~x11 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x64 && x21 && ~x10 && ~x12 && x17 && x16 && ~x19 && x18 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x63 && x64 && x21 && ~x10 && ~x12 && x17 && x16 && ~x19 && ~x18 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x64 && x21 && ~x10 && ~x12 && x17 && ~x16 && x11 )
						begin
							y3 = 1'b1;	
							nx_state = s788;
						end
					else if( ~x63 && x64 && x21 && ~x10 && ~x12 && x17 && ~x16 && ~x11 )
						begin
							y32 = 1'b1;	
							nx_state = s854;
						end
					else if( ~x63 && x64 && x21 && ~x10 && ~x12 && ~x17 && x16 && x19 && x14 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x63 && x64 && x21 && ~x10 && ~x12 && ~x17 && x16 && x19 && ~x14 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x64 && x21 && ~x10 && ~x12 && ~x17 && x16 && ~x19 && x13 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x63 && x64 && x21 && ~x10 && ~x12 && ~x17 && x16 && ~x19 && ~x13 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x64 && x21 && ~x10 && ~x12 && ~x17 && ~x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x64 && ~x21 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s937;
						end
					else if( ~x63 && x64 && ~x21 && ~x6 && x5 )
						begin
							y30 = 1'b1;	
							nx_state = s416;
						end
					else if( ~x63 && x64 && ~x21 && ~x6 && ~x5 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x63 && ~x64 )
						begin
							y42 = 1'b1;	
							nx_state = s1423;
						end
					else nx_state = s1083;
				s1084 : if( x17 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y16 = 1'b1;	y27 = 1'b1;	
							nx_state = s1432;
						end
					else if( ~x17 )
						begin
							y5 = 1'b1;	y13 = 1'b1;	y17 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1084;
						end
					else nx_state = s1084;
				s1085 : if( 1'b1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y12 = 1'b1;	
							y37 = 1'b1;	y38 = 1'b1;	
							nx_state = s1059;
						end
					else nx_state = s1085;
				s1086 : if( x16 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s442;
						end
					else if( ~x16 )
						begin
							y3 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s520;
						end
					else nx_state = s1086;
				s1087 : if( x16 && x22 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x16 && x22 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x16 && x22 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x16 && x22 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x16 && x22 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x16 && ~x22 )
						begin
							y3 = 1'b1;	y30 = 1'b1;	y31 = 1'b1;	
							nx_state = s741;
						end
					else if( ~x16 )
						begin
							y3 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s521;
						end
					else nx_state = s1087;
				s1088 : if( x22 )
						begin
							y17 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s418;
						end
					else if( ~x22 && x23 )
						begin
							y17 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s418;
						end
					else if( ~x22 && ~x23 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1433;
						end
					else nx_state = s1088;
				s1089 : if( x22 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1433;
						end
					else if( ~x22 && x23 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1433;
						end
					else if( ~x22 && ~x23 )
						begin
							y17 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s418;
						end
					else nx_state = s1089;
				s1090 : if( 1'b1 )
						begin
							y17 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s1434;
						end
					else nx_state = s1090;
				s1091 : if( x22 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1435;
						end
					else if( ~x22 )
						begin
							y17 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s1434;
						end
					else nx_state = s1091;
				s1092 : if( x22 && x16 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x22 && x16 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x22 && x16 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x22 && x16 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x22 && x16 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x22 && ~x16 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s657;
						end
					else if( ~x22 && x16 && x7 && x8 && x9 && x23 && x10 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y5 = 1'b1;	
							y22 = 1'b1;	y23 = 1'b1;	
							nx_state = s72;
						end
					else if( ~x22 && x16 && x7 && x8 && x9 && x23 && ~x10 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( ~x22 && x16 && x7 && x8 && x9 && ~x23 && x10 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y38 = 1'b1;	
							y46 = 1'b1;	
							nx_state = s741;
						end
					else if( ~x22 && x16 && x7 && x8 && x9 && ~x23 && ~x10 )
						begin
							y47 = 1'b1;	
							nx_state = s287;
						end
					else if( ~x22 && x16 && x7 && x8 && ~x9 && x23 && x10 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x22 && x16 && x7 && x8 && ~x9 && x23 && x10 && ~x13 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && x16 && x7 && x8 && ~x9 && x23 && x10 && ~x13 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && x16 && x7 && x8 && ~x9 && x23 && x10 && ~x13 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x22 && x16 && x7 && x8 && ~x9 && x23 && x10 && ~x13 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && x16 && x7 && x8 && ~x9 && x23 && x10 && ~x13 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x22 && x16 && x7 && x8 && ~x9 && x23 && ~x10 && x1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x22 && x16 && x7 && x8 && ~x9 && x23 && ~x10 && ~x1 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && x16 && x7 && x8 && ~x9 && x23 && ~x10 && ~x1 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && x16 && x7 && x8 && ~x9 && x23 && ~x10 && ~x1 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x22 && x16 && x7 && x8 && ~x9 && x23 && ~x10 && ~x1 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && x16 && x7 && x8 && ~x9 && x23 && ~x10 && ~x1 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x22 && x16 && x7 && x8 && ~x9 && ~x23 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y42 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s1042;
						end
					else if( ~x22 && x16 && x7 && ~x8 && x9 && x23 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x22 && x16 && x7 && ~x8 && x9 && ~x23 && x10 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y38 = 1'b1;	
							y40 = 1'b1;	y41 = 1'b1;	
							nx_state = s741;
						end
					else if( ~x22 && x16 && x7 && ~x8 && x9 && ~x23 && ~x10 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y38 = 1'b1;	
							y39 = 1'b1;	y41 = 1'b1;	
							nx_state = s741;
						end
					else if( ~x22 && x16 && x7 && ~x8 && ~x9 && x23 && x10 && x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x22 && x16 && x7 && ~x8 && ~x9 && x23 && x10 && ~x3 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && x16 && x7 && ~x8 && ~x9 && x23 && x10 && ~x3 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && x16 && x7 && ~x8 && ~x9 && x23 && x10 && ~x3 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x22 && x16 && x7 && ~x8 && ~x9 && x23 && x10 && ~x3 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && x16 && x7 && ~x8 && ~x9 && x23 && x10 && ~x3 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x22 && x16 && x7 && ~x8 && ~x9 && x23 && ~x10 && x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x22 && x16 && x7 && ~x8 && ~x9 && x23 && ~x10 && ~x15 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && x16 && x7 && ~x8 && ~x9 && x23 && ~x10 && ~x15 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && x16 && x7 && ~x8 && ~x9 && x23 && ~x10 && ~x15 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x22 && x16 && x7 && ~x8 && ~x9 && x23 && ~x10 && ~x15 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x22 && x16 && x7 && ~x8 && ~x9 && x23 && ~x10 && ~x15 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x22 && x16 && x7 && ~x8 && ~x9 && ~x23 )
						begin
							y5 = 1'b1;	y35 = 1'b1;	y36 = 1'b1;	
							y38 = 1'b1;	y41 = 1'b1;	
							nx_state = s741;
						end
					else if( ~x22 && x16 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s523;
						end
					else if( ~x22 && ~x16 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s524;
						end
					else nx_state = s1092;
				s1093 : if( 1'b1 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else nx_state = s1093;
				s1094 : if( 1'b1 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y21 = 1'b1;	
							nx_state = s1436;
						end
					else nx_state = s1094;
				s1095 : if( x3 && x9 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x3 && x9 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x3 && x9 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x3 && x9 && ~x14 )
						nx_state = s1;
					else if( x3 && ~x9 && x10 && x11 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y21 = 1'b1;	
							y26 = 1'b1;	y29 = 1'b1;	
							nx_state = s1430;
						end
					else if( x3 && ~x9 && x10 && ~x11 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y21 = 1'b1;	
							y26 = 1'b1;	y28 = 1'b1;	
							nx_state = s1430;
						end
					else if( x3 && ~x9 && ~x10 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y21 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s1430;
						end
					else if( ~x3 )
						begin
							y14 = 1'b1;	y37 = 1'b1;	y43 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s1437;
						end
					else nx_state = s1095;
				s1096 : if( x22 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							y18 = 1'b1;	y29 = 1'b1;	
							nx_state = s1001;
						end
					else if( x22 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1002;
						end
					else if( ~x22 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1002;
						end
					else if( ~x22 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							y18 = 1'b1;	y29 = 1'b1;	
							nx_state = s1001;
						end
					else nx_state = s1096;
				s1097 : if( x61 && x11 && x25 && x3 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( x61 && x11 && x25 && ~x3 && x5 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( x61 && x11 && x25 && ~x3 && ~x5 )
						nx_state = s1097;
					else if( x61 && x11 && ~x25 )
						begin
							y1 = 1'b1;	
							nx_state = s803;
						end
					else if( x61 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x61 && x53 && x47 )
						nx_state = s1097;
					else if( ~x61 && x53 && ~x47 && x59 && x51 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x61 && x53 && ~x47 && x59 && ~x51 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( ~x61 && x53 && ~x47 && ~x59 && x34 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s843;
						end
					else if( ~x61 && x53 && ~x47 && ~x59 && ~x34 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else if( ~x61 && ~x53 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s434;
						end
					else nx_state = s1097;
				s1098 : if( x63 && x65 && x20 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x63 && x65 && ~x20 )
						begin
							y62 = 1'b1;	
							nx_state = s1119;
						end
					else if( x63 && ~x65 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x65 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x65 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x63 && ~x65 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x65 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x63 && x64 && x65 && x10 )
						begin
							y62 = 1'b1;	
							nx_state = s1119;
						end
					else if( ~x63 && x64 && x65 && ~x10 && x4 && x5 && x3 && x12 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x63 && x64 && x65 && ~x10 && x4 && x5 && x3 && x12 && ~x8 && x7 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x63 && x64 && x65 && ~x10 && x4 && x5 && x3 && x12 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x63 && x64 && x65 && ~x10 && x4 && x5 && x3 && ~x12 )
						nx_state = s1;
					else if( ~x63 && x64 && x65 && ~x10 && x4 && x5 && ~x3 && x6 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x63 && x64 && x65 && ~x10 && x4 && x5 && ~x3 && x6 && ~x7 && x12 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x63 && x64 && x65 && ~x10 && x4 && x5 && ~x3 && x6 && ~x7 && x12 && ~x8 )
						nx_state = s1;
					else if( ~x63 && x64 && x65 && ~x10 && x4 && x5 && ~x3 && x6 && ~x7 && ~x12 )
						nx_state = s1;
					else if( ~x63 && x64 && x65 && ~x10 && x4 && x5 && ~x3 && ~x6 && x8 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x63 && x64 && x65 && ~x10 && x4 && x5 && ~x3 && ~x6 && ~x8 && x12 && x7 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x63 && x64 && x65 && ~x10 && x4 && x5 && ~x3 && ~x6 && ~x8 && x12 && ~x7 )
						nx_state = s1;
					else if( ~x63 && x64 && x65 && ~x10 && x4 && x5 && ~x3 && ~x6 && ~x8 && ~x12 )
						nx_state = s1;
					else if( ~x63 && x64 && x65 && ~x10 && x4 && ~x5 && x6 && x3 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x63 && x64 && x65 && ~x10 && x4 && ~x5 && x6 && ~x3 )
						begin
							y21 = 1'b1;	y38 = 1'b1;	
							nx_state = s412;
						end
					else if( ~x63 && x64 && x65 && ~x10 && x4 && ~x5 && ~x6 && x3 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x63 && x64 && x65 && ~x10 && x4 && ~x5 && ~x6 && ~x3 )
						begin
							y22 = 1'b1;	y29 = 1'b1;	
							nx_state = s412;
						end
					else if( ~x63 && x64 && x65 && ~x10 && ~x4 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x63 && x64 && ~x65 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s328;
						end
					else if( ~x63 && ~x64 && x65 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && ~x64 && x65 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && ~x64 && x65 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x63 && ~x64 && x65 && ~x15 )
						nx_state = s1;
					else if( ~x63 && ~x64 && ~x65 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x63 && ~x64 && ~x65 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x63 && ~x64 && ~x65 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x63 && ~x64 && ~x65 && ~x8 )
						nx_state = s1;
					else nx_state = s1098;
				s1099 : if( x3 )
						begin
							y5 = 1'b1;	
							nx_state = s560;
						end
					else if( ~x3 )
						begin
							y4 = 1'b1;	y62 = 1'b1;	y63 = 1'b1;	
							nx_state = s1145;
						end
					else nx_state = s1099;
				s1100 : if( x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y23 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1438;
						end
					else if( ~x8 && x10 && x9 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s1439;
						end
					else if( ~x8 && x10 && ~x9 )
						begin
							y58 = 1'b1;	
							nx_state = s1265;
						end
					else if( ~x8 && ~x10 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y26 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1440;
						end
					else if( ~x8 && ~x10 && ~x9 )
						begin
							y56 = 1'b1;	
							nx_state = s1219;
						end
					else nx_state = s1100;
				s1101 : if( 1'b1 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y21 = 1'b1;	
							y32 = 1'b1;	y35 = 1'b1;	
							nx_state = s1321;
						end
					else nx_state = s1101;
				s1102 : if( 1'b1 )
						begin
							y2 = 1'b1;	
							nx_state = s155;
						end
					else nx_state = s1102;
				s1103 : if( 1'b1 )
						begin
							y25 = 1'b1;	
							nx_state = s1441;
						end
					else nx_state = s1103;
				s1104 : if( x69 && x62 && x10 && x15 )
						nx_state = s1;
					else if( x69 && x62 && x10 && ~x15 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && x62 && ~x10 )
						nx_state = s1;
					else if( x69 && ~x62 && x17 && x18 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x5 && x6 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && ~x62 && x17 && x18 && ~x5 && ~x6 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( x69 && ~x62 && x17 && ~x18 && x3 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( x69 && ~x62 && x17 && ~x18 && ~x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( x69 && ~x62 && ~x17 && x18 && x1 )
						nx_state = s1;
					else if( x69 && ~x62 && ~x17 && x18 && ~x1 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( x69 && ~x62 && ~x17 && ~x18 )
						nx_state = s1;
					else if( ~x69 && x17 && x18 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1104;
						end
					else if( ~x69 && x17 && x18 && ~x5 && x6 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && x17 && x18 && ~x5 && ~x6 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x69 && x17 && ~x18 && x3 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s40;
						end
					else if( ~x69 && x17 && ~x18 && ~x3 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x69 && ~x17 && x16 && x18 && x1 && x15 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x69 && ~x17 && x16 && x18 && x1 && x15 && ~x5 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x69 && ~x17 && x16 && x18 && x1 && x15 && ~x5 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x69 && ~x17 && x16 && x18 && x1 && ~x15 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x17 && x16 && x18 && ~x1 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && ~x17 && x16 && ~x18 && x15 && x5 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x69 && ~x17 && x16 && ~x18 && x15 && ~x5 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x69 && ~x17 && x16 && ~x18 && x15 && ~x5 && ~x6 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x69 && ~x17 && x16 && ~x18 && ~x15 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x17 && ~x16 && x15 && x1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x17 && ~x16 && x15 && ~x1 && x18 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && ~x17 && ~x16 && x15 && ~x1 && ~x18 )
						nx_state = s1104;
					else if( ~x69 && ~x17 && ~x16 && ~x15 && x18 && x1 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x69 && ~x17 && ~x16 && ~x15 && x18 && x1 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x69 && ~x17 && ~x16 && ~x15 && x18 && ~x1 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x69 && ~x17 && ~x16 && ~x15 && ~x18 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x69 && ~x17 && ~x16 && ~x15 && ~x18 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else nx_state = s1104;
				s1105 : if( x62 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x62 && x64 && x40 && x50 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1106;
						end
					else if( ~x62 && x64 && x40 && ~x50 )
						nx_state = s1105;
					else if( ~x62 && x64 && ~x40 && x11 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s686;
						end
					else if( ~x62 && x64 && ~x40 && ~x11 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s686;
						end
					else if( ~x62 && x64 && ~x40 && ~x11 && ~x9 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x62 && ~x64 && x44 && x50 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s1107;
						end
					else if( ~x62 && ~x64 && x44 && ~x50 )
						nx_state = s1105;
					else if( ~x62 && ~x64 && ~x44 && x11 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s686;
						end
					else if( ~x62 && ~x64 && ~x44 && ~x11 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s686;
						end
					else if( ~x62 && ~x64 && ~x44 && ~x11 && ~x9 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else nx_state = s1105;
				s1106 : if( x40 && x17 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else if( x40 && ~x17 && x43 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( x40 && ~x17 && ~x43 )
						nx_state = s1106;
					else if( ~x40 && x6 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else if( ~x40 && ~x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1106;
						end
					else nx_state = s1106;
				s1107 : if( x44 && x17 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else if( x44 && ~x17 && x49 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( x44 && ~x17 && ~x49 )
						nx_state = s1107;
					else if( ~x44 && x6 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else if( ~x44 && ~x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s1107;
						end
					else nx_state = s1107;
				s1108 : if( x62 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s1442;
						end
					else if( ~x62 )
						begin
							y28 = 1'b1;	
							nx_state = s539;
						end
					else nx_state = s1108;
				s1109 : if( x65 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1443;
						end
					else if( ~x65 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else nx_state = s1109;
				s1110 : if( x31 && x30 )
						begin
							y30 = 1'b1;	
							nx_state = s976;
						end
					else if( x31 && ~x30 )
						begin
							y31 = 1'b1;	
							nx_state = s1072;
						end
					else if( ~x31 )
						begin
							y30 = 1'b1;	
							nx_state = s976;
						end
					else nx_state = s1110;
				s1111 : if( x63 && x19 && x18 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1286;
						end
					else if( x63 && x19 && ~x18 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s820;
						end
					else if( x63 && ~x19 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							y17 = 1'b1;	y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1238;
						end
					else if( ~x63 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							nx_state = s1444;
						end
					else nx_state = s1111;
				s1112 : if( 1'b1 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1286;
						end
					else nx_state = s1112;
				s1113 : if( 1'b1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y9 = 1'b1;	
							y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s433;
						end
					else nx_state = s1113;
				s1114 : if( 1'b1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s759;
						end
					else nx_state = s1114;
				s1115 : if( x63 && x20 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s936;
						end
					else if( x63 && ~x20 )
						begin
							y28 = 1'b1;	
							nx_state = s991;
						end
					else if( ~x63 )
						begin
							y6 = 1'b1;	
							nx_state = s239;
						end
					else nx_state = s1115;
				s1116 : if( 1'b1 )
						begin
							y28 = 1'b1;	
							nx_state = s1445;
						end
					else nx_state = s1116;
				s1117 : if( 1'b1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y48 = 1'b1;	y50 = 1'b1;	
							nx_state = s1446;
						end
					else nx_state = s1117;
				s1118 : if( x18 && x26 && x14 && x27 && x6 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s1448;
						end
					else if( x18 && x26 && x14 && x27 && x6 && ~x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s677;
						end
					else if( x18 && x26 && x14 && x27 && ~x6 && x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s1447;
						end
					else if( x18 && x26 && x14 && x27 && ~x6 && ~x5 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							nx_state = s1199;
						end
					else if( x18 && x26 && x14 && ~x27 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s1220;
						end
					else if( x18 && x26 && x14 && ~x27 && ~x5 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							nx_state = s1199;
						end
					else if( x18 && x26 && ~x14 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s1448;
						end
					else if( x18 && x26 && ~x14 && ~x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s677;
						end
					else if( x18 && ~x26 && x27 && x14 && x5 )
						begin
							y50 = 1'b1;	
							nx_state = s658;
						end
					else if( x18 && ~x26 && x27 && x14 && ~x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s1447;
						end
					else if( x18 && ~x26 && x27 && ~x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s1448;
						end
					else if( x18 && ~x26 && ~x27 && x7 && x6 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x18 && ~x26 && ~x27 && x7 && x6 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x18 && ~x26 && ~x27 && x7 && x6 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x18 && ~x26 && ~x27 && x7 && x6 && x22 && ~x23 )
						nx_state = s1;
					else if( x18 && ~x26 && ~x27 && x7 && x6 && ~x22 )
						nx_state = s1;
					else if( x18 && ~x26 && ~x27 && x7 && ~x6 && x8 && x15 )
						begin
							y10 = 1'b1;	
							nx_state = s405;
						end
					else if( x18 && ~x26 && ~x27 && x7 && ~x6 && x8 && ~x15 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x18 && ~x26 && ~x27 && x7 && ~x6 && x8 && ~x15 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x18 && ~x26 && ~x27 && x7 && ~x6 && x8 && ~x15 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x18 && ~x26 && ~x27 && x7 && ~x6 && x8 && ~x15 && x22 && ~x23 )
						nx_state = s1;
					else if( x18 && ~x26 && ~x27 && x7 && ~x6 && x8 && ~x15 && ~x22 )
						nx_state = s1;
					else if( x18 && ~x26 && ~x27 && x7 && ~x6 && ~x8 && x16 )
						begin
							y10 = 1'b1;	
							nx_state = s405;
						end
					else if( x18 && ~x26 && ~x27 && x7 && ~x6 && ~x8 && ~x16 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x18 && ~x26 && ~x27 && x7 && ~x6 && ~x8 && ~x16 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x18 && ~x26 && ~x27 && x7 && ~x6 && ~x8 && ~x16 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x18 && ~x26 && ~x27 && x7 && ~x6 && ~x8 && ~x16 && x22 && ~x23 )
						nx_state = s1;
					else if( x18 && ~x26 && ~x27 && x7 && ~x6 && ~x8 && ~x16 && ~x22 )
						nx_state = s1;
					else if( x18 && ~x26 && ~x27 && ~x7 && x8 && x6 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x18 && ~x26 && ~x27 && ~x7 && x8 && ~x6 )
						begin
							y5 = 1'b1;	y44 = 1'b1;	y55 = 1'b1;	
							y60 = 1'b1;	
							nx_state = s1220;
						end
					else if( x18 && ~x26 && ~x27 && ~x7 && ~x8 && x6 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x18 && ~x26 && ~x27 && ~x7 && ~x8 && ~x6 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y53 = 1'b1;	
							y54 = 1'b1;	
							nx_state = s1220;
						end
					else if( ~x18 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s1449;
						end
					else nx_state = s1118;
				s1119 : if( x63 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x63 && ~x18 )
						begin
							y44 = 1'b1;	
							nx_state = s755;
						end
					else if( ~x63 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else nx_state = s1119;
				s1120 : if( x63 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x63 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x63 )
						begin
							y63 = 1'b1;	
							nx_state = s483;
						end
					else nx_state = s1120;
				s1121 : if( x62 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							nx_state = s1450;
						end
					else if( ~x62 )
						begin
							y28 = 1'b1;	
							nx_state = s1326;
						end
					else nx_state = s1121;
				s1122 : if( 1'b1 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else nx_state = s1122;
				s1123 : if( x63 && x26 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( x63 && ~x26 )
						begin
							y66 = 1'b1;	
							nx_state = s726;
						end
					else if( ~x63 && x65 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x65 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x65 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x63 && x65 && ~x15 )
						nx_state = s1;
					else if( ~x63 && ~x65 && x20 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x63 && ~x65 && ~x20 )
						nx_state = s1;
					else nx_state = s1123;
				s1124 : if( x26 )
						begin
							y11 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x26 && x28 && x36 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s1170;
						end
					else if( ~x26 && x28 && ~x36 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s542;
						end
					else if( ~x26 && ~x28 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s995;
						end
					else nx_state = s1124;
				s1125 : if( x55 && x34 )
						begin
							y11 = 1'b1;	y29 = 1'b1;	
							nx_state = s818;
						end
					else if( x55 && ~x34 && x2 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x55 && ~x34 && ~x2 && x28 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s503;
						end
					else if( x55 && ~x34 && ~x2 && ~x28 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s502;
						end
					else if( ~x55 && x41 && x36 && x3 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( ~x55 && x41 && x36 && ~x3 && x4 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else if( ~x55 && x41 && x36 && ~x3 && ~x4 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s630;
						end
					else if( ~x55 && x41 && ~x36 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x55 && ~x41 && x11 && x32 )
						begin
							y10 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s882;
						end
					else if( ~x55 && ~x41 && x11 && ~x32 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s499;
						end
					else if( ~x55 && ~x41 && x11 && ~x32 && ~x3 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x55 && ~x41 && ~x11 )
						nx_state = s1125;
					else nx_state = s1125;
				s1126 : if( x55 && x50 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( x55 && ~x50 )
						nx_state = s1126;
					else if( ~x55 && x42 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s1125;
						end
					else if( ~x55 && ~x42 && x9 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s1125;
						end
					else if( ~x55 && ~x42 && ~x9 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s629;
						end
					else nx_state = s1126;
				s1127 : if( x44 && x1 && x37 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( x44 && x1 && ~x37 && x9 )
						nx_state = s1127;
					else if( x44 && x1 && ~x37 && ~x9 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s154;
						end
					else if( x44 && ~x1 && x9 )
						begin
							y2 = 1'b1;	y20 = 1'b1;	y25 = 1'b1;	
							nx_state = s500;
						end
					else if( x44 && ~x1 && ~x9 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x44 && x10 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else if( ~x44 && ~x10 && x11 && x37 )
						begin
							y3 = 1'b1;	y13 = 1'b1;	y22 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s640;
						end
					else if( ~x44 && ~x10 && x11 && ~x37 && x41 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s512;
						end
					else if( ~x44 && ~x10 && x11 && ~x37 && ~x41 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x44 && ~x10 && ~x11 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s138;
						end
					else nx_state = s1127;
				s1128 : if( 1'b1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s105;
						end
					else nx_state = s1128;
				s1129 : if( x3 )
						begin
							y5 = 1'b1;	
							nx_state = s645;
						end
					else if( ~x3 && x21 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y62 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s1189;
						end
					else if( ~x3 && ~x21 )
						begin
							y4 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y78 = 1'b1;	
							nx_state = s1190;
						end
					else nx_state = s1129;
				s1130 : if( x21 && x3 )
						begin
							y4 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y79 = 1'b1;	
							nx_state = s1451;
						end
					else if( x21 && ~x3 )
						begin
							y62 = 1'b1;	y65 = 1'b1;	y71 = 1'b1;	
							y90 = 1'b1;	
							nx_state = s1451;
						end
					else if( ~x21 && x22 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s950;
						end
					else if( ~x21 && x22 && ~x3 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y62 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s1189;
						end
					else if( ~x21 && ~x22 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x21 && ~x22 && ~x3 )
						begin
							y4 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y78 = 1'b1;	
							nx_state = s587;
						end
					else nx_state = s1130;
				s1131 : if( x21 && x3 )
						begin
							y62 = 1'b1;	y65 = 1'b1;	y78 = 1'b1;	
							y96 = 1'b1;	
							nx_state = s1392;
						end
					else if( x21 && ~x3 )
						begin
							y60 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y79 = 1'b1;	
							nx_state = s1392;
						end
					else if( ~x21 && x22 && x3 )
						begin
							y4 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y78 = 1'b1;	
							nx_state = s1393;
						end
					else if( ~x21 && x22 && ~x3 )
						begin
							y62 = 1'b1;	y81 = 1'b1;	
							nx_state = s1393;
						end
					else if( ~x21 && ~x22 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s791;
						end
					else if( ~x21 && ~x22 && ~x3 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y62 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s1189;
						end
					else nx_state = s1131;
				s1132 : if( 1'b1 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1026;
						end
					else nx_state = s1132;
				s1133 : if( x21 && x3 )
						begin
							y62 = 1'b1;	y64 = 1'b1;	y65 = 1'b1;	
							y78 = 1'b1;	
							nx_state = s1452;
						end
					else if( x21 && ~x3 )
						begin
							y62 = 1'b1;	y65 = 1'b1;	y79 = 1'b1;	
							y88 = 1'b1;	y102 = 1'b1;	
							nx_state = s1452;
						end
					else if( ~x21 && x3 )
						begin
							y62 = 1'b1;	y65 = 1'b1;	y78 = 1'b1;	
							y96 = 1'b1;	
							nx_state = s1392;
						end
					else if( ~x21 && ~x3 )
						begin
							y60 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y79 = 1'b1;	
							nx_state = s1392;
						end
					else nx_state = s1133;
				s1134 : if( x21 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s950;
						end
					else if( x21 && ~x3 )
						begin
							y4 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y93 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x21 && x22 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s791;
						end
					else if( ~x21 && x22 && ~x3 )
						begin
							y4 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y78 = 1'b1;	
							nx_state = s1190;
						end
					else if( ~x21 && ~x22 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s950;
						end
					else if( ~x21 && ~x22 && ~x3 )
						begin
							y4 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y78 = 1'b1;	
							nx_state = s1354;
						end
					else nx_state = s1134;
				s1135 : if( x3 )
						begin
							y5 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x3 )
						begin
							y4 = 1'b1;	y62 = 1'b1;	y73 = 1'b1;	
							nx_state = s1453;
						end
					else nx_state = s1135;
				s1136 : if( x21 && x10 )
						begin
							y62 = 1'b1;	y65 = 1'b1;	y78 = 1'b1;	
							y90 = 1'b1;	
							nx_state = s1132;
						end
					else if( x21 && ~x10 && x14 && x11 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1130;
						end
					else if( x21 && ~x10 && x14 && ~x11 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1133;
						end
					else if( x21 && ~x10 && ~x14 && x11 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1134;
						end
					else if( x21 && ~x10 && ~x14 && ~x11 )
						begin
							y3 = 1'b1;	y74 = 1'b1;	
							nx_state = s1135;
						end
					else if( ~x21 && x10 && x22 && x11 && x14 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1134;
						end
					else if( ~x21 && x10 && x22 && x11 && ~x14 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1131;
						end
					else if( ~x21 && x10 && x22 && ~x11 && x14 && x19 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x21 && x10 && x22 && ~x11 && x14 && ~x19 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x10 && x22 && ~x11 && x14 && ~x19 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x10 && x22 && ~x11 && x14 && ~x19 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x10 && x22 && ~x11 && x14 && ~x19 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x10 && x22 && ~x11 && ~x14 && x18 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x21 && x10 && x22 && ~x11 && ~x14 && ~x18 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x10 && x22 && ~x11 && ~x14 && ~x18 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x10 && x22 && ~x11 && ~x14 && ~x18 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x10 && x22 && ~x11 && ~x14 && ~x18 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x10 && ~x22 )
						begin
							y9 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y94 = 1'b1;	
							nx_state = s849;
						end
					else if( ~x21 && ~x10 && x22 && x14 && x11 && x17 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x21 && ~x10 && x22 && x14 && x11 && ~x17 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && ~x10 && x22 && x14 && x11 && ~x17 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && ~x10 && x22 && x14 && x11 && ~x17 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x10 && x22 && x14 && x11 && ~x17 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x10 && x22 && x14 && ~x11 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x21 && ~x10 && x22 && ~x14 && x11 && x16 && x18 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x21 && ~x10 && x22 && ~x14 && x11 && x16 && ~x18 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && ~x10 && x22 && ~x14 && x11 && x16 && ~x18 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && ~x10 && x22 && ~x14 && x11 && x16 && ~x18 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x10 && x22 && ~x14 && x11 && x16 && ~x18 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x10 && x22 && ~x14 && x11 && ~x16 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && ~x10 && x22 && ~x14 && x11 && ~x16 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && ~x10 && x22 && ~x14 && x11 && ~x16 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x10 && x22 && ~x14 && x11 && ~x16 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x10 && x22 && ~x14 && ~x11 )
						begin
							y102 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x21 && ~x10 && ~x22 )
						begin
							y9 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y94 = 1'b1;	
							nx_state = s844;
						end
					else nx_state = s1136;
				s1137 : if( x63 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x63 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x63 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x63 && ~x1 )
						nx_state = s1;
					else if( ~x63 && x64 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x63 && x64 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x63 && x64 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x63 && x64 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x63 && x64 && ~x22 )
						nx_state = s1;
					else if( ~x63 && ~x64 && x21 && x22 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x63 && ~x64 && x21 && ~x22 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x63 && ~x64 && x21 && ~x22 && ~x23 )
						nx_state = s1;
					else if( ~x63 && ~x64 && ~x21 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x63 && ~x64 && ~x21 && ~x23 )
						nx_state = s1;
					else nx_state = s1137;
				s1138 : if( x64 && x63 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x64 && x63 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x64 && x63 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x64 && x63 && ~x11 )
						nx_state = s1;
					else if( x64 && ~x63 && x65 )
						begin
							y4 = 1'b1;	y20 = 1'b1;	y31 = 1'b1;	
							nx_state = s1029;
						end
					else if( x64 && ~x63 && ~x65 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x64 && ~x63 && ~x65 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x64 && ~x63 && ~x65 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x64 && ~x63 && ~x65 && ~x14 )
						nx_state = s1;
					else if( ~x64 && x63 && x66 && x16 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x64 && x63 && x66 && x16 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x64 && x63 && x66 && x16 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x64 && x63 && x66 && ~x16 )
						nx_state = s1;
					else if( ~x64 && x63 && ~x66 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x64 && x63 && ~x66 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x64 && x63 && ~x66 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x64 && x63 && ~x66 && ~x1 )
						nx_state = s1;
					else if( ~x64 && ~x63 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else nx_state = s1138;
				s1139 : if( 1'b1 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1454;
						end
					else nx_state = s1139;
				s1140 : if( x3 && x5 && x7 && x9 && x11 )
						begin
							y26 = 1'b1;	
							nx_state = s262;
						end
					else if( x3 && x5 && x7 && x9 && ~x11 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( x3 && x5 && x7 && ~x9 && x10 && x11 && x12 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( x3 && x5 && x7 && ~x9 && x10 && x11 && ~x12 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x3 && x5 && x7 && ~x9 && x10 && x11 && ~x12 && x19 && ~x13 )
						nx_state = s1;
					else if( x3 && x5 && x7 && ~x9 && x10 && x11 && ~x12 && ~x19 )
						nx_state = s1;
					else if( x3 && x5 && x7 && ~x9 && x10 && ~x11 && x13 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( x3 && x5 && x7 && ~x9 && x10 && ~x11 && ~x13 && x19 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x3 && x5 && x7 && ~x9 && x10 && ~x11 && ~x13 && x19 && ~x12 )
						nx_state = s1;
					else if( x3 && x5 && x7 && ~x9 && x10 && ~x11 && ~x13 && ~x19 )
						nx_state = s1;
					else if( x3 && x5 && x7 && ~x9 && ~x10 && x11 )
						begin
							y5 = 1'b1;	y18 = 1'b1;	y27 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s1455;
						end
					else if( x3 && x5 && x7 && ~x9 && ~x10 && ~x11 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1455;
						end
					else if( x3 && x5 && ~x7 )
						begin
							y3 = 1'b1;	y6 = 1'b1;	y9 = 1'b1;	
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s1456;
						end
					else if( x3 && ~x5 && x8 && x7 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s1455;
						end
					else if( x3 && ~x5 && x8 && ~x7 && x9 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x3 && ~x5 && x8 && ~x7 && x9 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x3 && ~x5 && x8 && ~x7 && x9 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x3 && ~x5 && x8 && ~x7 && x9 && ~x19 )
						nx_state = s1;
					else if( x3 && ~x5 && x8 && ~x7 && ~x9 && x10 && x11 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s1455;
						end
					else if( x3 && ~x5 && x8 && ~x7 && ~x9 && x10 && ~x11 )
						begin
							y3 = 1'b1;	y18 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s1455;
						end
					else if( x3 && ~x5 && x8 && ~x7 && ~x9 && ~x10 )
						begin
							y3 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	y29 = 1'b1;	
							nx_state = s1455;
						end
					else if( x3 && ~x5 && ~x8 )
						begin
							y3 = 1'b1;	y6 = 1'b1;	y9 = 1'b1;	
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s1456;
						end
					else if( ~x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s1457;
						end
					else nx_state = s1140;
				s1141 : if( 1'b1 )
						begin
							y28 = 1'b1;	
							nx_state = s717;
						end
					else nx_state = s1141;
				s1142 : if( 1'b1 )
						begin
							y28 = 1'b1;	
							nx_state = s1458;
						end
					else nx_state = s1142;
				s1143 : if( x16 && x15 && x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( x16 && x15 && ~x5 )
						begin
							y21 = 1'b1;	y27 = 1'b1;	
							nx_state = s930;
						end
					else if( x16 && ~x15 && x4 && x5 && x34 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( x16 && ~x15 && x4 && x5 && ~x34 && x1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y15 = 1'b1;	
							nx_state = s455;
						end
					else if( x16 && ~x15 && x4 && x5 && ~x34 && ~x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s931;
						end
					else if( x16 && ~x15 && x4 && ~x5 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( x16 && ~x15 && ~x4 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x16 && x15 && x13 && x11 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s439;
						end
					else if( ~x16 && x15 && x13 && ~x11 && x6 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x16 && x15 && x13 && ~x11 && x6 && ~x4 && x37 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s550;
						end
					else if( ~x16 && x15 && x13 && ~x11 && x6 && ~x4 && ~x37 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s549;
						end
					else if( ~x16 && x15 && x13 && ~x11 && ~x6 && x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	y33 = 1'b1;	
							nx_state = s931;
						end
					else if( ~x16 && x15 && x13 && ~x11 && ~x6 && ~x5 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s325;
						end
					else if( ~x16 && x15 && ~x13 && x14 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x16 && x15 && ~x13 && ~x14 && x9 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x16 && x15 && ~x13 && ~x14 && ~x9 && x6 && x2 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x16 && x15 && ~x13 && ~x14 && ~x9 && x6 && ~x2 )
						nx_state = s1143;
					else if( ~x16 && x15 && ~x13 && ~x14 && ~x9 && ~x6 && x8 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s547;
						end
					else if( ~x16 && x15 && ~x13 && ~x14 && ~x9 && ~x6 && ~x8 )
						nx_state = s1143;
					else if( ~x16 && ~x15 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else nx_state = s1143;
				s1144 : if( 1'b1 )
						begin
							y13 = 1'b1;	
							nx_state = s800;
						end
					else nx_state = s1144;
				s1145 : if( x4 && x22 && x21 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x4 && x22 && ~x21 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( x4 && ~x22 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x4 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s146;
						end
					else nx_state = s1145;
				s1146 : if( 1'b1 )
						begin
							y5 = 1'b1;	
							nx_state = s266;
						end
					else nx_state = s1146;
				s1147 : if( 1'b1 )
						begin
							y5 = 1'b1;	
							nx_state = s64;
						end
					else nx_state = s1147;
				s1148 : if( 1'b1 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else nx_state = s1148;
				s1149 : if( 1'b1 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s367;
						end
					else nx_state = s1149;
				s1150 : if( 1'b1 )
						begin
							y6 = 1'b1;	
							nx_state = s431;
						end
					else nx_state = s1150;
				s1151 : if( x4 && x19 && x20 && x14 )
						begin
							y16 = 1'b1;	y28 = 1'b1;	
							nx_state = s1459;
						end
					else if( x4 && x19 && x20 && ~x14 && x16 )
						begin
							y16 = 1'b1;	y28 = 1'b1;	
							nx_state = s1459;
						end
					else if( x4 && x19 && x20 && ~x14 && ~x16 && x17 )
						begin
							y16 = 1'b1;	y28 = 1'b1;	
							nx_state = s865;
						end
					else if( x4 && x19 && x20 && ~x14 && ~x16 && ~x17 )
						begin
							y16 = 1'b1;	y28 = 1'b1;	
							nx_state = s1459;
						end
					else if( x4 && x19 && ~x20 )
						begin
							y16 = 1'b1;	y28 = 1'b1;	
							nx_state = s1459;
						end
					else if( x4 && ~x19 )
						begin
							y16 = 1'b1;	y28 = 1'b1;	
							nx_state = s1459;
						end
					else if( ~x4 && x9 && x17 && x19 && x20 && x14 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x4 && x9 && x17 && x19 && x20 && ~x14 && x16 )
						begin
							y4 = 1'b1;	y29 = 1'b1;	y32 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x4 && x9 && x17 && x19 && x20 && ~x14 && ~x16 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s868;
						end
					else if( ~x4 && x9 && x17 && x19 && ~x20 && x14 )
						begin
							y4 = 1'b1;	y18 = 1'b1;	y29 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x4 && x9 && x17 && x19 && ~x20 && ~x14 && x16 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	y32 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x4 && x9 && x17 && x19 && ~x20 && ~x14 && ~x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x4 && x9 && x17 && ~x19 && x16 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x4 && x9 && x17 && ~x19 && ~x16 && x20 )
						begin
							y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s863;
						end
					else if( ~x4 && x9 && x17 && ~x19 && ~x16 && ~x20 && x15 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x4 && x9 && x17 && ~x19 && ~x16 && ~x20 && ~x15 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x4 && x9 && ~x17 && x18 && x19 && x14 && x16 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	y19 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s861;
						end
					else if( ~x4 && x9 && ~x17 && x18 && x19 && x14 && ~x16 )
						begin
							y2 = 1'b1;	y21 = 1'b1;	
							nx_state = s1318;
						end
					else if( ~x4 && x9 && ~x17 && x18 && x19 && ~x14 )
						begin
							y7 = 1'b1;	
							nx_state = s747;
						end
					else if( ~x4 && x9 && ~x17 && x18 && ~x19 )
						begin
							y7 = 1'b1;	
							nx_state = s747;
						end
					else if( ~x4 && x9 && ~x17 && ~x18 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x4 && ~x9 && x19 && x20 && x17 && x16 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s868;
						end
					else if( ~x4 && ~x9 && x19 && x20 && x17 && ~x16 && x14 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s868;
						end
					else if( ~x4 && ~x9 && x19 && x20 && x17 && ~x16 && ~x14 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( ~x4 && ~x9 && x19 && x20 && ~x17 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s868;
						end
					else if( ~x4 && ~x9 && x19 && ~x20 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s868;
						end
					else if( ~x4 && ~x9 && ~x19 && x20 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s868;
						end
					else if( ~x4 && ~x9 && ~x19 && ~x20 && x17 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s868;
						end
					else if( ~x4 && ~x9 && ~x19 && ~x20 && ~x17 && x18 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x4 && ~x9 && ~x19 && ~x20 && ~x17 && ~x18 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s868;
						end
					else nx_state = s1151;
				s1152 : if( 1'b1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y37 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s1460;
						end
					else nx_state = s1152;
				s1153 : if( 1'b1 )
						begin
							y5 = 1'b1;	
							nx_state = s937;
						end
					else nx_state = s1153;
				s1154 : if( 1'b1 )
						begin
							y37 = 1'b1;	y40 = 1'b1;	y41 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s1461;
						end
					else nx_state = s1154;
				s1155 : if( 1'b1 )
						begin
							y5 = 1'b1;	
							nx_state = s560;
						end
					else nx_state = s1155;
				s1156 : if( x39 && x41 && x42 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y40 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s1154;
						end
					else if( x39 && x41 && ~x42 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y40 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s584;
						end
					else if( x39 && ~x41 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y37 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s939;
						end
					else if( ~x39 && x40 && x55 && x56 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x39 && x40 && x55 && ~x56 && x58 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( ~x39 && x40 && x55 && ~x56 && ~x58 && x59 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x39 && x40 && x55 && ~x56 && ~x58 && ~x59 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x39 && x40 && x55 && ~x56 && ~x58 && ~x59 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x39 && x40 && x55 && ~x56 && ~x58 && ~x59 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( ~x39 && x40 && x55 && ~x56 && ~x58 && ~x59 && ~x27 )
						nx_state = s1;
					else if( ~x39 && x40 && ~x55 && x54 && x57 && x28 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x39 && x40 && ~x55 && x54 && x57 && ~x28 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x39 && x40 && ~x55 && x54 && x57 && ~x28 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x39 && x40 && ~x55 && x54 && x57 && ~x28 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( ~x39 && x40 && ~x55 && x54 && x57 && ~x28 && ~x27 )
						nx_state = s1;
					else if( ~x39 && x40 && ~x55 && x54 && ~x57 && x29 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x39 && x40 && ~x55 && x54 && ~x57 && ~x29 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x39 && x40 && ~x55 && x54 && ~x57 && ~x29 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x39 && x40 && ~x55 && x54 && ~x57 && ~x29 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( ~x39 && x40 && ~x55 && x54 && ~x57 && ~x29 && ~x27 )
						nx_state = s1;
					else if( ~x39 && x40 && ~x55 && ~x54 && x53 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x39 && x40 && ~x55 && ~x54 && ~x53 )
						begin
							y30 = 1'b1;	
							nx_state = s291;
						end
					else if( ~x39 && ~x40 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y37 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s1155;
						end
					else nx_state = s1156;
				s1157 : if( x62 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else if( ~x62 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s1462;
						end
					else if( ~x62 && ~x14 )
						begin
							y47 = 1'b1;	y56 = 1'b1;	y61 = 1'b1;	
							y70 = 1'b1;	
							nx_state = s1463;
						end
					else nx_state = s1157;
				s1158 : if( 1'b1 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y44 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s1464;
						end
					else nx_state = s1158;
				s1159 : if( x51 && x41 && x42 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y40 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s1154;
						end
					else if( x51 && x41 && ~x42 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y40 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s584;
						end
					else if( x51 && ~x41 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y37 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s939;
						end
					else if( ~x51 && x52 && x55 && x56 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x51 && x52 && x55 && ~x56 && x58 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( ~x51 && x52 && x55 && ~x56 && ~x58 && x59 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x51 && x52 && x55 && ~x56 && ~x58 && ~x59 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x51 && x52 && x55 && ~x56 && ~x58 && ~x59 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x51 && x52 && x55 && ~x56 && ~x58 && ~x59 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( ~x51 && x52 && x55 && ~x56 && ~x58 && ~x59 && ~x27 )
						nx_state = s1;
					else if( ~x51 && x52 && ~x55 && x54 && x57 && x28 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x51 && x52 && ~x55 && x54 && x57 && ~x28 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x51 && x52 && ~x55 && x54 && x57 && ~x28 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x51 && x52 && ~x55 && x54 && x57 && ~x28 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( ~x51 && x52 && ~x55 && x54 && x57 && ~x28 && ~x27 )
						nx_state = s1;
					else if( ~x51 && x52 && ~x55 && x54 && ~x57 && x29 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x51 && x52 && ~x55 && x54 && ~x57 && ~x29 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x51 && x52 && ~x55 && x54 && ~x57 && ~x29 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x51 && x52 && ~x55 && x54 && ~x57 && ~x29 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( ~x51 && x52 && ~x55 && x54 && ~x57 && ~x29 && ~x27 )
						nx_state = s1;
					else if( ~x51 && x52 && ~x55 && ~x54 && x53 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s584;
						end
					else if( ~x51 && x52 && ~x55 && ~x54 && ~x53 )
						begin
							y30 = 1'b1;	
							nx_state = s291;
						end
					else if( ~x51 && ~x52 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y37 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s1147;
						end
					else nx_state = s1159;
				s1160 : if( 1'b1 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y39 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s1465;
						end
					else nx_state = s1160;
				s1161 : if( 1'b1 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y39 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s1466;
						end
					else nx_state = s1161;
				s1162 : if( 1'b1 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y39 = 1'b1;	
							nx_state = s584;
						end
					else nx_state = s1162;
				s1163 : if( 1'b1 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y39 = 1'b1;	
							nx_state = s584;
						end
					else nx_state = s1163;
				s1164 : if( x9 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x9 )
						nx_state = s1164;
					else nx_state = s1164;
				s1165 : if( x63 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x63 && ~x15 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x63 && x64 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && ~x64 )
						begin
							y4 = 1'b1;	
							nx_state = s403;
						end
					else nx_state = s1165;
				s1166 : if( x4 )
						begin
							y8 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x4 && x31 && x30 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x4 && x31 && ~x30 )
						begin
							y37 = 1'b1;	
							nx_state = s1467;
						end
					else if( ~x4 && ~x31 && x30 )
						begin
							y37 = 1'b1;	
							nx_state = s1467;
						end
					else if( ~x4 && ~x31 && ~x30 )
						begin
							y37 = 1'b1;	
							nx_state = s1356;
						end
					else nx_state = s1166;
				s1167 : if( x20 && x12 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x20 && ~x12 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x20 && ~x12 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x20 && ~x12 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x20 && ~x12 && x22 && ~x23 )
						nx_state = s1;
					else if( x20 && ~x12 && ~x22 )
						nx_state = s1;
					else if( ~x20 )
						begin
							y26 = 1'b1;	
							nx_state = s1468;
						end
					else nx_state = s1167;
				s1168 : if( 1'b1 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s894;
						end
					else nx_state = s1168;
				s1169 : if( x3 && x4 && x5 && x21 && x7 && x9 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x3 && x4 && x5 && x21 && x7 && ~x9 )
						begin
							y50 = 1'b1;	
							nx_state = s658;
						end
					else if( x3 && x4 && x5 && x21 && ~x7 && x8 && x9 && x12 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x3 && x4 && x5 && x21 && ~x7 && x8 && x9 && ~x12 && x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x3 && x4 && x5 && x21 && ~x7 && x8 && x9 && ~x12 && x10 && ~x11 )
						nx_state = s1;
					else if( x3 && x4 && x5 && x21 && ~x7 && x8 && x9 && ~x12 && ~x10 )
						nx_state = s1;
					else if( x3 && x4 && x5 && x21 && ~x7 && x8 && ~x9 && x11 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x3 && x4 && x5 && x21 && ~x7 && x8 && ~x9 && ~x11 && x10 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x3 && x4 && x5 && x21 && ~x7 && x8 && ~x9 && ~x11 && x10 && ~x12 )
						nx_state = s1;
					else if( x3 && x4 && x5 && x21 && ~x7 && x8 && ~x9 && ~x11 && ~x10 )
						nx_state = s1;
					else if( x3 && x4 && x5 && x21 && ~x7 && ~x8 && x9 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y39 = 1'b1;	y40 = 1'b1;	
							nx_state = s1263;
						end
					else if( x3 && x4 && x5 && x21 && ~x7 && ~x8 && ~x9 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y16 = 1'b1;	
							y42 = 1'b1;	y51 = 1'b1;	
							nx_state = s1263;
						end
					else if( x3 && x4 && x5 && ~x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s731;
						end
					else if( x3 && x4 && ~x5 && x13 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s1469;
						end
					else if( x3 && x4 && ~x5 && ~x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s731;
						end
					else if( x3 && ~x4 )
						begin
							y6 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s1470;
						end
					else if( ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s1471;
						end
					else nx_state = s1169;
				s1170 : if( 1'b1 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else nx_state = s1170;
				s1171 : if( x9 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s941;
						end
					else if( ~x9 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else nx_state = s1171;
				s1172 : if( x64 && x3 )
						begin
							y14 = 1'b1;	
							nx_state = s124;
						end
					else if( x64 && ~x3 )
						begin
							y31 = 1'b1;	
							nx_state = s1472;
						end
					else if( ~x64 )
						begin
							y47 = 1'b1;	y53 = 1'b1;	y61 = 1'b1;	
							y70 = 1'b1;	
							nx_state = s1473;
						end
					else nx_state = s1172;
				s1173 : if( x63 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	y25 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x63 && x30 )
						begin
							y47 = 1'b1;	y49 = 1'b1;	y58 = 1'b1;	
							y61 = 1'b1;	y68 = 1'b1;	
							nx_state = s1297;
						end
					else if( ~x63 && ~x30 && x31 )
						begin
							y35 = 1'b1;	
							nx_state = s414;
						end
					else if( ~x63 && ~x30 && ~x31 )
						begin
							y31 = 1'b1;	
							nx_state = s1053;
						end
					else nx_state = s1173;
				s1174 : if( 1'b1 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else nx_state = s1174;
				s1175 : if( x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x23 )
						nx_state = s1;
					else nx_state = s1175;
				s1176 : if( 1'b1 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else nx_state = s1176;
				s1177 : if( 1'b1 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							y17 = 1'b1;	y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1238;
						end
					else nx_state = s1177;
				s1178 : if( 1'b1 )
						begin
							y3 = 1'b1;	y17 = 1'b1;	y19 = 1'b1;	
							nx_state = s1474;
						end
					else nx_state = s1178;
				s1179 : if( x66 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x66 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s1179;
				s1180 : if( 1'b1 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else nx_state = s1180;
				s1181 : if( x20 && x21 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x20 && ~x21 && x4 && x6 && x14 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( x20 && ~x21 && x4 && x6 && ~x14 )
						begin
							y6 = 1'b1;	y40 = 1'b1;	y41 = 1'b1;	
							y42 = 1'b1;	
							nx_state = s1475;
						end
					else if( x20 && ~x21 && x4 && ~x6 )
						begin
							y20 = 1'b1;	
							nx_state = s1261;
						end
					else if( x20 && ~x21 && ~x4 )
						begin
							y20 = 1'b1;	
							nx_state = s1476;
						end
					else if( ~x20 && x4 && x6 && x13 && x21 && x14 && x15 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else if( ~x20 && x4 && x6 && x13 && x21 && x14 && ~x15 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( ~x20 && x4 && x6 && x13 && x21 && x14 && ~x15 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( ~x20 && x4 && x6 && x13 && x21 && ~x14 && x15 && x17 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( ~x20 && x4 && x6 && x13 && x21 && ~x14 && x15 && x17 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( ~x20 && x4 && x6 && x13 && x21 && ~x14 && x15 && ~x17 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && x4 && x6 && x13 && x21 && ~x14 && x15 && ~x17 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && x4 && x6 && x13 && x21 && ~x14 && x15 && ~x17 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x20 && x4 && x6 && x13 && x21 && ~x14 && x15 && ~x17 && ~x10 )
						nx_state = s1;
					else if( ~x20 && x4 && x6 && x13 && x21 && ~x14 && ~x15 && x9 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( ~x20 && x4 && x6 && x13 && x21 && ~x14 && ~x15 && x9 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( ~x20 && x4 && x6 && x13 && x21 && ~x14 && ~x15 && ~x9 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && x4 && x6 && x13 && x21 && ~x14 && ~x15 && ~x9 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && x4 && x6 && x13 && x21 && ~x14 && ~x15 && ~x9 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x20 && x4 && x6 && x13 && x21 && ~x14 && ~x15 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x20 && x4 && x6 && x13 && ~x21 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1259;
						end
					else if( ~x20 && x4 && x6 && ~x13 && x21 && x14 && x15 && x18 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( ~x20 && x4 && x6 && ~x13 && x21 && x14 && x15 && x18 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( ~x20 && x4 && x6 && ~x13 && x21 && x14 && x15 && ~x18 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && x4 && x6 && ~x13 && x21 && x14 && x15 && ~x18 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && x4 && x6 && ~x13 && x21 && x14 && x15 && ~x18 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x20 && x4 && x6 && ~x13 && x21 && x14 && x15 && ~x18 && ~x10 )
						nx_state = s1;
					else if( ~x20 && x4 && x6 && ~x13 && x21 && x14 && ~x15 && x19 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( ~x20 && x4 && x6 && ~x13 && x21 && x14 && ~x15 && x19 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( ~x20 && x4 && x6 && ~x13 && x21 && x14 && ~x15 && ~x19 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && x4 && x6 && ~x13 && x21 && x14 && ~x15 && ~x19 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && x4 && x6 && ~x13 && x21 && x14 && ~x15 && ~x19 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x20 && x4 && x6 && ~x13 && x21 && x14 && ~x15 && ~x19 && ~x10 )
						nx_state = s1;
					else if( ~x20 && x4 && x6 && ~x13 && x21 && ~x14 && x15 && x5 )
						begin
							y14 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x20 && x4 && x6 && ~x13 && x21 && ~x14 && x15 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1207;
						end
					else if( ~x20 && x4 && x6 && ~x13 && x21 && ~x14 && ~x15 && x7 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1208;
						end
					else if( ~x20 && x4 && x6 && ~x13 && x21 && ~x14 && ~x15 && ~x7 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1209;
						end
					else if( ~x20 && x4 && x6 && ~x13 && ~x21 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && x4 && x6 && ~x13 && ~x21 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && x4 && x6 && ~x13 && ~x21 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x20 && x4 && x6 && ~x13 && ~x21 && ~x10 )
						nx_state = s1;
					else if( ~x20 && x4 && ~x6 )
						begin
							y20 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x20 && ~x4 )
						begin
							y20 = 1'b1;	
							nx_state = s1261;
						end
					else nx_state = s1181;
				s1182 : if( x69 && x64 && x15 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( x69 && x64 && ~x15 && x14 && x13 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s691;
						end
					else if( x69 && x64 && ~x15 && x14 && ~x13 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s478;
						end
					else if( x69 && x64 && ~x15 && ~x14 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s638;
						end
					else if( x69 && ~x64 && x14 && x13 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s691;
						end
					else if( x69 && ~x64 && x14 && ~x13 && x66 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s498;
						end
					else if( x69 && ~x64 && x14 && ~x13 && ~x66 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x69 && ~x64 && ~x14 && x66 )
						begin
							y19 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s994;
						end
					else if( x69 && ~x64 && ~x14 && ~x66 )
						begin
							y12 = 1'b1;	
							nx_state = s246;
						end
					else if( ~x69 && x62 && x15 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s451;
						end
					else if( ~x69 && x62 && ~x15 && x14 && x13 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s1105;
						end
					else if( ~x69 && x62 && ~x15 && x14 && ~x13 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s901;
						end
					else if( ~x69 && x62 && ~x15 && ~x14 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x69 && ~x62 && x63 && x46 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y33 = 1'b1;	
							nx_state = s1236;
						end
					else if( ~x69 && ~x62 && x63 && ~x46 && x44 && x11 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( ~x69 && ~x62 && x63 && ~x46 && x44 && ~x11 && x6 && x35 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s997;
						end
					else if( ~x69 && ~x62 && x63 && ~x46 && x44 && ~x11 && x6 && ~x35 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y27 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s998;
						end
					else if( ~x69 && ~x62 && x63 && ~x46 && x44 && ~x11 && ~x6 && x36 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( ~x69 && ~x62 && x63 && ~x46 && x44 && ~x11 && ~x6 && ~x36 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y31 = 1'b1;	y35 = 1'b1;	
							nx_state = s996;
						end
					else if( ~x69 && ~x62 && x63 && ~x46 && ~x44 && x14 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s693;
						end
					else if( ~x69 && ~x62 && x63 && ~x46 && ~x44 && ~x14 && x9 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s693;
						end
					else if( ~x69 && ~x62 && x63 && ~x46 && ~x44 && ~x14 && ~x9 && x37 && x33 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s693;
						end
					else if( ~x69 && ~x62 && x63 && ~x46 && ~x44 && ~x14 && ~x9 && x37 && ~x33 )
						nx_state = s1182;
					else if( ~x69 && ~x62 && x63 && ~x46 && ~x44 && ~x14 && ~x9 && ~x37 && x8 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s693;
						end
					else if( ~x69 && ~x62 && x63 && ~x46 && ~x44 && ~x14 && ~x9 && ~x37 && ~x8 )
						nx_state = s1182;
					else if( ~x69 && ~x62 && ~x63 && x14 && x13 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s691;
						end
					else if( ~x69 && ~x62 && ~x63 && x14 && ~x13 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s1234;
						end
					else if( ~x69 && ~x62 && ~x63 && ~x14 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s704;
						end
					else nx_state = s1182;
				s1183 : if( x14 && x13 )
						begin
							y19 = 1'b1;	y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s1215;
						end
					else if( x14 && ~x13 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s1234;
						end
					else if( ~x14 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s704;
						end
					else nx_state = s1183;
				s1184 : if( x33 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x33 )
						begin
							y20 = 1'b1;	y23 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s914;
						end
					else nx_state = s1184;
				s1185 : if( x25 )
						nx_state = s1;
					else if( ~x25 && x28 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( ~x25 && ~x28 )
						nx_state = s1;
					else nx_state = s1185;
				s1186 : if( 1'b1 )
						begin
							y6 = 1'b1;	
							nx_state = s649;
						end
					else nx_state = s1186;
				s1187 : if( 1'b1 )
						begin
							y27 = 1'b1;	
							nx_state = s1083;
						end
					else nx_state = s1187;
				s1188 : if( 1'b1 )
						begin
							y13 = 1'b1;	
							nx_state = s897;
						end
					else nx_state = s1188;
				s1189 : if( x13 && x21 && x10 )
						begin
							y62 = 1'b1;	y65 = 1'b1;	y78 = 1'b1;	
							y90 = 1'b1;	
							nx_state = s1132;
						end
					else if( x13 && x21 && ~x10 && x14 && x11 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1130;
						end
					else if( x13 && x21 && ~x10 && x14 && ~x11 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1133;
						end
					else if( x13 && x21 && ~x10 && ~x14 && x11 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1134;
						end
					else if( x13 && x21 && ~x10 && ~x14 && ~x11 )
						begin
							y3 = 1'b1;	y74 = 1'b1;	
							nx_state = s1135;
						end
					else if( x13 && ~x21 && x10 && x22 && x11 && x14 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1134;
						end
					else if( x13 && ~x21 && x10 && x22 && x11 && ~x14 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1131;
						end
					else if( x13 && ~x21 && x10 && x22 && ~x11 && x14 && x19 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( x13 && ~x21 && x10 && x22 && ~x11 && x14 && ~x19 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x13 && ~x21 && x10 && x22 && ~x11 && x14 && ~x19 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x13 && ~x21 && x10 && x22 && ~x11 && x14 && ~x19 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x13 && ~x21 && x10 && x22 && ~x11 && x14 && ~x19 && ~x6 )
						nx_state = s1;
					else if( x13 && ~x21 && x10 && x22 && ~x11 && ~x14 && x18 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( x13 && ~x21 && x10 && x22 && ~x11 && ~x14 && ~x18 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x13 && ~x21 && x10 && x22 && ~x11 && ~x14 && ~x18 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x13 && ~x21 && x10 && x22 && ~x11 && ~x14 && ~x18 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x13 && ~x21 && x10 && x22 && ~x11 && ~x14 && ~x18 && ~x6 )
						nx_state = s1;
					else if( x13 && ~x21 && x10 && ~x22 )
						begin
							y9 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y94 = 1'b1;	
							nx_state = s849;
						end
					else if( x13 && ~x21 && ~x10 && x22 && x14 && x11 && x17 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( x13 && ~x21 && ~x10 && x22 && x14 && x11 && ~x17 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x13 && ~x21 && ~x10 && x22 && x14 && x11 && ~x17 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x13 && ~x21 && ~x10 && x22 && x14 && x11 && ~x17 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x13 && ~x21 && ~x10 && x22 && x14 && x11 && ~x17 && ~x6 )
						nx_state = s1;
					else if( x13 && ~x21 && ~x10 && x22 && x14 && ~x11 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( x13 && ~x21 && ~x10 && x22 && ~x14 && x11 && x16 && x18 )
						begin
							y12 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s516;
						end
					else if( x13 && ~x21 && ~x10 && x22 && ~x14 && x11 && x16 && ~x18 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x13 && ~x21 && ~x10 && x22 && ~x14 && x11 && x16 && ~x18 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x13 && ~x21 && ~x10 && x22 && ~x14 && x11 && x16 && ~x18 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x13 && ~x21 && ~x10 && x22 && ~x14 && x11 && x16 && ~x18 && ~x6 )
						nx_state = s1;
					else if( x13 && ~x21 && ~x10 && x22 && ~x14 && x11 && ~x16 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x13 && ~x21 && ~x10 && x22 && ~x14 && x11 && ~x16 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x13 && ~x21 && ~x10 && x22 && ~x14 && x11 && ~x16 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x13 && ~x21 && ~x10 && x22 && ~x14 && x11 && ~x16 && ~x6 )
						nx_state = s1;
					else if( x13 && ~x21 && ~x10 && x22 && ~x14 && ~x11 )
						begin
							y102 = 1'b1;	
							nx_state = s516;
						end
					else if( x13 && ~x21 && ~x10 && ~x22 )
						begin
							y9 = 1'b1;	y62 = 1'b1;	y65 = 1'b1;	
							y94 = 1'b1;	
							nx_state = s844;
						end
					else if( ~x13 )
						begin
							y9 = 1'b1;	y65 = 1'b1;	y84 = 1'b1;	
							y86 = 1'b1;	y91 = 1'b1;	
							nx_state = s1136;
						end
					else nx_state = s1189;
				s1190 : if( x22 )
						begin
							y54 = 1'b1;	
							nx_state = s281;
						end
					else if( ~x22 )
						begin
							y60 = 1'b1;	y65 = 1'b1;	y78 = 1'b1;	
							y92 = 1'b1;	
							nx_state = s1477;
						end
					else nx_state = s1190;
				s1191 : if( x10 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s1478;
						end
					else if( ~x10 )
						begin
							y28 = 1'b1;	
							nx_state = s991;
						end
					else nx_state = s1191;
				s1192 : if( 1'b1 )
						begin
							y14 = 1'b1;	
							nx_state = s366;
						end
					else nx_state = s1192;
				s1193 : if( x18 )
						begin
							y19 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x18 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x18 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x18 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x18 && ~x19 )
						nx_state = s1;
					else nx_state = s1193;
				s1194 : if( x65 )
						begin
							y8 = 1'b1;	
							nx_state = s642;
						end
					else if( ~x65 )
						begin
							y7 = 1'b1;	
							nx_state = s1358;
						end
					else nx_state = s1194;
				s1195 : if( 1'b1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1479;
						end
					else nx_state = s1195;
				s1196 : if( 1'b1 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else nx_state = s1196;
				s1197 : if( x64 )
						begin
							y27 = 1'b1;	
							nx_state = s893;
						end
					else if( ~x64 && x66 && x14 )
						begin
							y29 = 1'b1;	
							nx_state = s1017;
						end
					else if( ~x64 && x66 && ~x14 )
						begin
							y28 = 1'b1;	y30 = 1'b1;	
							nx_state = s1164;
						end
					else if( ~x64 && ~x66 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else nx_state = s1197;
				s1198 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	y26 = 1'b1;	
							nx_state = s1313;
						end
					else nx_state = s1198;
				s1199 : if( x26 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x26 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x26 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x26 && x22 && ~x23 )
						nx_state = s1;
					else if( x26 && ~x22 )
						nx_state = s1;
					else if( ~x26 && x12 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x26 && x12 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x26 && x12 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x26 && x12 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x26 && x12 && ~x22 )
						nx_state = s1;
					else if( ~x26 && ~x12 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else nx_state = s1199;
				s1200 : if( x65 )
						begin
							y8 = 1'b1;	
							nx_state = s786;
						end
					else if( ~x65 )
						begin
							y7 = 1'b1;	
							nx_state = s1194;
						end
					else nx_state = s1200;
				s1201 : if( 1'b1 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else nx_state = s1201;
				s1202 : if( 1'b1 )
						begin
							y4 = 1'b1;	y18 = 1'b1;	y20 = 1'b1;	
							nx_state = s1480;
						end
					else nx_state = s1202;
				s1203 : if( x7 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1481;
						end
					else if( ~x7 && x8 && x20 && x14 && x15 )
						begin
							y6 = 1'b1;	y11 = 1'b1;	y26 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1307;
						end
					else if( ~x7 && x8 && x20 && x14 && ~x15 )
						begin
							y6 = 1'b1;	y11 = 1'b1;	y42 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1068;
						end
					else if( ~x7 && x8 && x20 && ~x14 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y44 = 1'b1;	
							y45 = 1'b1;	y49 = 1'b1;	
							nx_state = s1482;
						end
					else if( ~x7 && x8 && ~x20 && x13 && x21 && x14 && x15 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else if( ~x7 && x8 && ~x20 && x13 && x21 && x14 && ~x15 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( ~x7 && x8 && ~x20 && x13 && x21 && x14 && ~x15 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( ~x7 && x8 && ~x20 && x13 && x21 && ~x14 && x15 && x17 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( ~x7 && x8 && ~x20 && x13 && x21 && ~x14 && x15 && x17 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( ~x7 && x8 && ~x20 && x13 && x21 && ~x14 && x15 && ~x17 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x7 && x8 && ~x20 && x13 && x21 && ~x14 && x15 && ~x17 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x7 && x8 && ~x20 && x13 && x21 && ~x14 && x15 && ~x17 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x7 && x8 && ~x20 && x13 && x21 && ~x14 && x15 && ~x17 && ~x10 )
						nx_state = s1;
					else if( ~x7 && x8 && ~x20 && x13 && x21 && ~x14 && ~x15 && x9 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( ~x7 && x8 && ~x20 && x13 && x21 && ~x14 && ~x15 && x9 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( ~x7 && x8 && ~x20 && x13 && x21 && ~x14 && ~x15 && ~x9 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x7 && x8 && ~x20 && x13 && x21 && ~x14 && ~x15 && ~x9 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x7 && x8 && ~x20 && x13 && x21 && ~x14 && ~x15 && ~x9 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x7 && x8 && ~x20 && x13 && x21 && ~x14 && ~x15 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x7 && x8 && ~x20 && x13 && ~x21 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							nx_state = s1213;
						end
					else if( ~x7 && x8 && ~x20 && ~x13 && x14 && x21 && x15 && x18 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( ~x7 && x8 && ~x20 && ~x13 && x14 && x21 && x15 && x18 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( ~x7 && x8 && ~x20 && ~x13 && x14 && x21 && x15 && ~x18 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x7 && x8 && ~x20 && ~x13 && x14 && x21 && x15 && ~x18 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x7 && x8 && ~x20 && ~x13 && x14 && x21 && x15 && ~x18 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x7 && x8 && ~x20 && ~x13 && x14 && x21 && x15 && ~x18 && ~x10 )
						nx_state = s1;
					else if( ~x7 && x8 && ~x20 && ~x13 && x14 && x21 && ~x15 && x19 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( ~x7 && x8 && ~x20 && ~x13 && x14 && x21 && ~x15 && x19 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( ~x7 && x8 && ~x20 && ~x13 && x14 && x21 && ~x15 && ~x19 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x7 && x8 && ~x20 && ~x13 && x14 && x21 && ~x15 && ~x19 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x7 && x8 && ~x20 && ~x13 && x14 && x21 && ~x15 && ~x19 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x7 && x8 && ~x20 && ~x13 && x14 && x21 && ~x15 && ~x19 && ~x10 )
						nx_state = s1;
					else if( ~x7 && x8 && ~x20 && ~x13 && x14 && ~x21 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y22 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s722;
						end
					else if( ~x7 && x8 && ~x20 && ~x13 && ~x14 && x21 && x15 && x5 )
						begin
							y14 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x7 && x8 && ~x20 && ~x13 && ~x14 && x21 && x15 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1207;
						end
					else if( ~x7 && x8 && ~x20 && ~x13 && ~x14 && x21 && ~x15 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1209;
						end
					else if( ~x7 && x8 && ~x20 && ~x13 && ~x14 && ~x21 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x7 && x8 && ~x20 && ~x13 && ~x14 && ~x21 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x7 && x8 && ~x20 && ~x13 && ~x14 && ~x21 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x7 && x8 && ~x20 && ~x13 && ~x14 && ~x21 && ~x10 )
						nx_state = s1;
					else if( ~x7 && ~x8 )
						begin
							y6 = 1'b1;	y9 = 1'b1;	y25 = 1'b1;	
							y56 = 1'b1;	
							nx_state = s1483;
						end
					else nx_state = s1203;
				s1204 : if( 1'b1 )
						begin
							y14 = 1'b1;	
							nx_state = s124;
						end
					else nx_state = s1204;
				s1205 : if( x20 && x21 )
						begin
							y6 = 1'b1;	y17 = 1'b1;	y34 = 1'b1;	
							nx_state = s226;
						end
					else if( x20 && ~x21 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s1484;
						end
					else if( ~x20 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s1485;
						end
					else nx_state = s1205;
				s1206 : if( 1'b1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1205;
						end
					else nx_state = s1206;
				s1207 : if( 1'b1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1486;
						end
					else nx_state = s1207;
				s1208 : if( x21 && x20 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1205;
						end
					else if( x21 && ~x20 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1487;
						end
					else if( ~x21 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1205;
						end
					else nx_state = s1208;
				s1209 : if( 1'b1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y22 = 1'b1;	
							y32 = 1'b1;	y33 = 1'b1;	
							nx_state = s949;
						end
					else nx_state = s1209;
				s1210 : if( x20 )
						begin
							y6 = 1'b1;	y41 = 1'b1;	y43 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s1488;
						end
					else if( ~x20 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s1381;
						end
					else if( ~x20 && ~x9 )
						begin
							y22 = 1'b1;	
							nx_state = s823;
						end
					else nx_state = s1210;
				s1211 : if( x21 && x20 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x21 && x20 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x21 && x20 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x21 && x20 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x20 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y22 = 1'b1;	
							y32 = 1'b1;	y33 = 1'b1;	
							nx_state = s1489;
						end
					else if( ~x21 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x21 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x21 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x21 && ~x10 )
						nx_state = s1;
					else nx_state = s1211;
				s1212 : if( 1'b1 )
						begin
							y55 = 1'b1;	
							nx_state = s773;
						end
					else nx_state = s1212;
				s1213 : if( x20 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y22 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s722;
						end
					else if( ~x20 && x21 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s953;
						end
					else if( ~x20 && x21 && ~x9 && x17 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y22 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s722;
						end
					else if( ~x20 && x21 && ~x9 && ~x17 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && x21 && ~x9 && ~x17 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && x21 && ~x9 && ~x17 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x20 && x21 && ~x9 && ~x17 && ~x10 )
						nx_state = s1;
					else if( ~x20 && ~x21 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && ~x21 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && ~x21 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x20 && ~x21 && ~x10 )
						nx_state = s1;
					else nx_state = s1213;
				s1214 : if( 1'b1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	y44 = 1'b1;	
							nx_state = s1490;
						end
					else nx_state = s1214;
				s1215 : if( 1'b1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s216;
						end
					else nx_state = s1215;
				s1216 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y33 = 1'b1;	
							y60 = 1'b1;	y61 = 1'b1;	y62 = 1'b1;	
							nx_state = s1491;
						end
					else nx_state = s1216;
				s1217 : if( 1'b1 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s1492;
						end
					else nx_state = s1217;
				s1218 : if( x6 && x8 && x7 )
						begin
							y63 = 1'b1;	
							nx_state = s483;
						end
					else if( x6 && x8 && ~x7 && x9 && x18 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y45 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s672;
						end
					else if( x6 && x8 && ~x7 && x9 && ~x18 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x6 && x8 && ~x7 && x9 && ~x18 && x20 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x6 && x8 && ~x7 && x9 && ~x18 && x20 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x6 && x8 && ~x7 && x9 && ~x18 && ~x20 )
						nx_state = s1;
					else if( x6 && x8 && ~x7 && ~x9 && x19 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y45 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s672;
						end
					else if( x6 && x8 && ~x7 && ~x9 && ~x19 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x6 && x8 && ~x7 && ~x9 && ~x19 && x20 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x6 && x8 && ~x7 && ~x9 && ~x19 && x20 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x6 && x8 && ~x7 && ~x9 && ~x19 && ~x20 )
						nx_state = s1;
					else if( x6 && ~x8 && x9 && x7 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y5 = 1'b1;	
							y74 = 1'b1;	
							nx_state = s1217;
						end
					else if( x6 && ~x8 && x9 && ~x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y45 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s672;
						end
					else if( x6 && ~x8 && ~x9 && x7 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y45 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s672;
						end
					else if( x6 && ~x8 && ~x9 && x7 && ~x17 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x6 && ~x8 && ~x9 && x7 && ~x17 && x20 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x6 && ~x8 && ~x9 && x7 && ~x17 && x20 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x6 && ~x8 && ~x9 && x7 && ~x17 && ~x20 )
						nx_state = s1;
					else if( x6 && ~x8 && ~x9 && ~x7 )
						begin
							y65 = 1'b1;	
							nx_state = s393;
						end
					else if( ~x6 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else nx_state = s1218;
				s1219 : if( x63 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y38 = 1'b1;	
							y57 = 1'b1;	
							nx_state = s741;
						end
					else if( ~x63 )
						begin
							y55 = 1'b1;	
							nx_state = s526;
						end
					else nx_state = s1219;
				s1220 : if( x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x22 && ~x23 )
						nx_state = s1;
					else if( ~x22 )
						nx_state = s1;
					else nx_state = s1220;
				s1221 : if( 1'b1 )
						begin
							y11 = 1'b1;	
							nx_state = s91;
						end
					else nx_state = s1221;
				s1222 : if( x8 )
						begin
							y5 = 1'b1;	y17 = 1'b1;	y32 = 1'b1;	
							y42 = 1'b1;	
							nx_state = s1220;
						end
					else if( ~x8 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x8 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x8 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x8 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x8 && ~x22 )
						nx_state = s1;
					else nx_state = s1222;
				s1223 : if( x63 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x63 && ~x18 )
						begin
							y44 = 1'b1;	
							nx_state = s755;
						end
					else if( ~x63 )
						begin
							y58 = 1'b1;	
							nx_state = s1265;
						end
					else nx_state = s1223;
				s1224 : if( x63 )
						begin
							y68 = 1'b1;	
							nx_state = s1404;
						end
					else if( ~x63 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s328;
						end
					else nx_state = s1224;
				s1225 : if( x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x17 )
						nx_state = s1;
					else nx_state = s1225;
				s1226 : if( x66 && x11 && x13 && x15 && x14 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	
							nx_state = s220;
						end
					else if( x66 && x11 && x13 && x15 && ~x14 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y58 = 1'b1;	
							nx_state = s1493;
						end
					else if( x66 && x11 && x13 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y59 = 1'b1;	
							nx_state = s1494;
						end
					else if( x66 && x11 && x13 && ~x15 && ~x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y29 = 1'b1;	
							nx_state = s1495;
						end
					else if( x66 && x11 && ~x13 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && x11 && ~x13 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && x11 && ~x13 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x66 && x11 && ~x13 && ~x8 )
						nx_state = s1;
					else if( x66 && ~x11 && x12 && x15 && x13 && x14 )
						begin
							y61 = 1'b1;	
							nx_state = s1098;
						end
					else if( x66 && ~x11 && x12 && x15 && x13 && ~x14 && x16 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( x66 && ~x11 && x12 && x15 && x13 && ~x14 && ~x16 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && ~x11 && x12 && x15 && x13 && ~x14 && ~x16 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && ~x11 && x12 && x15 && x13 && ~x14 && ~x16 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x66 && ~x11 && x12 && x15 && x13 && ~x14 && ~x16 && ~x8 )
						nx_state = s1;
					else if( x66 && ~x11 && x12 && x15 && ~x13 && x14 && x18 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1078;
						end
					else if( x66 && ~x11 && x12 && x15 && ~x13 && x14 && ~x18 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && ~x11 && x12 && x15 && ~x13 && x14 && ~x18 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && ~x11 && x12 && x15 && ~x13 && x14 && ~x18 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x66 && ~x11 && x12 && x15 && ~x13 && x14 && ~x18 && ~x8 )
						nx_state = s1;
					else if( x66 && ~x11 && x12 && x15 && ~x13 && ~x14 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x66 && ~x11 && x12 && ~x15 && x13 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( x66 && ~x11 && x12 && ~x15 && x13 && ~x14 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( x66 && ~x11 && x12 && ~x15 && x13 && ~x14 && ~x17 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && ~x11 && x12 && ~x15 && x13 && ~x14 && ~x17 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && ~x11 && x12 && ~x15 && x13 && ~x14 && ~x17 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x66 && ~x11 && x12 && ~x15 && x13 && ~x14 && ~x17 && ~x8 )
						nx_state = s1;
					else if( x66 && ~x11 && x12 && ~x15 && ~x13 && x14 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y62 = 1'b1;	
							nx_state = s1496;
						end
					else if( x66 && ~x11 && x12 && ~x15 && ~x13 && ~x14 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && ~x11 && x12 && ~x15 && ~x13 && ~x14 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && ~x11 && x12 && ~x15 && ~x13 && ~x14 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x66 && ~x11 && x12 && ~x15 && ~x13 && ~x14 && ~x8 )
						nx_state = s1;
					else if( x66 && ~x11 && ~x12 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y29 = 1'b1;	
							nx_state = s1497;
						end
					else if( ~x66 && x20 && x5 && x6 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y23 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x66 && x20 && x5 && ~x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y25 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x66 && x20 && ~x5 )
						begin
							y3 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y30 = 1'b1;	y43 = 1'b1;	
							nx_state = s1345;
						end
					else if( ~x66 && ~x20 && x4 && x21 && x6 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s1270;
						end
					else if( ~x66 && ~x20 && x4 && x21 && x6 && ~x5 && x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x66 && ~x20 && x4 && x21 && x6 && ~x5 && ~x11 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x66 && ~x20 && x4 && x21 && x6 && ~x5 && ~x11 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x66 && ~x20 && x4 && x21 && x6 && ~x5 && ~x11 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x66 && ~x20 && x4 && x21 && x6 && ~x5 && ~x11 && ~x17 )
						nx_state = s1;
					else if( ~x66 && ~x20 && x4 && x21 && ~x6 && x5 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y15 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1347;
						end
					else if( ~x66 && ~x20 && x4 && x21 && ~x6 && ~x5 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x66 && ~x20 && x4 && x21 && ~x6 && ~x5 && ~x10 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x66 && ~x20 && x4 && x21 && ~x6 && ~x5 && ~x10 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x66 && ~x20 && x4 && x21 && ~x6 && ~x5 && ~x10 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x66 && ~x20 && x4 && x21 && ~x6 && ~x5 && ~x10 && ~x17 )
						nx_state = s1;
					else if( ~x66 && ~x20 && x4 && ~x21 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x66 && ~x20 && ~x4 && x21 && x6 && x5 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x66 && ~x20 && ~x4 && x21 && x6 && x5 && ~x13 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x66 && ~x20 && ~x4 && x21 && x6 && x5 && ~x13 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x66 && ~x20 && ~x4 && x21 && x6 && x5 && ~x13 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x66 && ~x20 && ~x4 && x21 && x6 && x5 && ~x13 && ~x17 )
						nx_state = s1;
					else if( ~x66 && ~x20 && ~x4 && x21 && x6 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x66 && ~x20 && ~x4 && x21 && ~x6 && x5 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x66 && ~x20 && ~x4 && x21 && ~x6 && x5 && ~x14 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x66 && ~x20 && ~x4 && x21 && ~x6 && x5 && ~x14 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x66 && ~x20 && ~x4 && x21 && ~x6 && x5 && ~x14 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x66 && ~x20 && ~x4 && x21 && ~x6 && x5 && ~x14 && ~x17 )
						nx_state = s1;
					else if( ~x66 && ~x20 && ~x4 && x21 && ~x6 && ~x5 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x66 && ~x20 && ~x4 && ~x21 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y23 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s1225;
						end
					else nx_state = s1226;
				s1227 : if( x7 )
						begin
							y33 = 1'b1;	y34 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x7 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x7 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x7 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x7 && ~x17 )
						nx_state = s1;
					else nx_state = s1227;
				s1228 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1498;
						end
					else nx_state = s1228;
				s1229 : if( x7 )
						begin
							y31 = 1'b1;	y32 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x7 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x7 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x7 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x7 && ~x17 )
						nx_state = s1;
					else nx_state = s1229;
				s1230 : if( x63 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x63 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else nx_state = s1230;
				s1231 : if( x21 && x20 )
						begin
							y22 = 1'b1;	
							nx_state = s39;
						end
					else if( x21 && ~x20 )
						begin
							y22 = 1'b1;	
							nx_state = s1108;
						end
					else if( ~x21 )
						begin
							y22 = 1'b1;	
							nx_state = s39;
						end
					else nx_state = s1231;
				s1232 : if( x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s480;
						end
					else if( ~x3 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s628;
						end
					else nx_state = s1232;
				s1233 : if( x62 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s125;
						end
					else if( ~x62 && x15 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s627;
						end
					else if( ~x62 && ~x15 && x12 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s1234;
						end
					else if( ~x62 && ~x15 && ~x12 )
						nx_state = s1233;
					else nx_state = s1233;
				s1234 : if( x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s216;
						end
					else if( ~x15 && x13 && x11 && x64 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s694;
						end
					else if( ~x15 && x13 && x11 && ~x64 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y28 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s703;
						end
					else if( ~x15 && x13 && ~x11 && x6 && x4 && x64 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	
							nx_state = s997;
						end
					else if( ~x15 && x13 && ~x11 && x6 && x4 && ~x64 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s999;
						end
					else if( ~x15 && x13 && ~x11 && x6 && ~x4 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1000;
						end
					else if( ~x15 && x13 && ~x11 && ~x6 && x5 )
						begin
							y15 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s695;
						end
					else if( ~x15 && x13 && ~x11 && ~x6 && ~x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s477;
						end
					else if( ~x15 && ~x13 && x14 && x64 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s693;
						end
					else if( ~x15 && ~x13 && x14 && ~x64 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s702;
						end
					else if( ~x15 && ~x13 && ~x14 && x9 && x64 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s693;
						end
					else if( ~x15 && ~x13 && ~x14 && x9 && ~x64 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s702;
						end
					else if( ~x15 && ~x13 && ~x14 && ~x9 && x6 && x64 && x2 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s693;
						end
					else if( ~x15 && ~x13 && ~x14 && ~x9 && x6 && x64 && ~x2 )
						nx_state = s1234;
					else if( ~x15 && ~x13 && ~x14 && ~x9 && x6 && ~x64 && x33 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s702;
						end
					else if( ~x15 && ~x13 && ~x14 && ~x9 && x6 && ~x64 && ~x33 )
						nx_state = s1234;
					else if( ~x15 && ~x13 && ~x14 && ~x9 && ~x6 && x64 && x8 )
						begin
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s693;
						end
					else if( ~x15 && ~x13 && ~x14 && ~x9 && ~x6 && x64 && ~x8 )
						nx_state = s1234;
					else if( ~x15 && ~x13 && ~x14 && ~x9 && ~x6 && ~x64 && x8 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s702;
						end
					else if( ~x15 && ~x13 && ~x14 && ~x9 && ~x6 && ~x64 && ~x8 )
						nx_state = s1234;
					else nx_state = s1234;
				s1235 : if( 1'b1 )
						begin
							y22 = 1'b1;	
							nx_state = s683;
						end
					else nx_state = s1235;
				s1236 : if( x26 && x28 && x32 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( x26 && x28 && ~x32 && x2 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( x26 && x28 && ~x32 && ~x2 && x25 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( x26 && x28 && ~x32 && ~x2 && ~x25 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( x26 && ~x28 && x32 && x33 && x34 && x25 )
						nx_state = s1236;
					else if( x26 && ~x28 && x32 && x33 && x34 && ~x25 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( x26 && ~x28 && x32 && x33 && ~x34 && x35 && x36 )
						begin
							y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s919;
						end
					else if( x26 && ~x28 && x32 && x33 && ~x34 && x35 && ~x36 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( x26 && ~x28 && x32 && x33 && ~x34 && ~x35 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( x26 && ~x28 && x32 && ~x33 )
						begin
							y11 = 1'b1;	
							nx_state = s247;
						end
					else if( x26 && ~x28 && ~x32 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( ~x26 && x28 && x27 )
						begin
							y11 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x26 && x28 && ~x27 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s496;
						end
					else if( ~x26 && x28 && ~x27 && ~x1 && x4 )
						begin
							y16 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s918;
						end
					else if( ~x26 && x28 && ~x27 && ~x1 && ~x4 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x26 && ~x28 )
						begin
							y11 = 1'b1;	
							nx_state = s247;
						end
					else nx_state = s1236;
				s1237 : if( x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s216;
						end
					else if( ~x15 && x13 && x4 )
						begin
							y23 = 1'b1;	y30 = 1'b1;	
							nx_state = s999;
						end
					else if( ~x15 && x13 && ~x4 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1000;
						end
					else if( ~x15 && ~x13 && x14 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s700;
						end
					else if( ~x15 && ~x13 && ~x14 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s700;
						end
					else if( ~x15 && ~x13 && ~x14 && ~x9 && x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s700;
						end
					else if( ~x15 && ~x13 && ~x14 && ~x9 && ~x7 && x8 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s700;
						end
					else if( ~x15 && ~x13 && ~x14 && ~x9 && ~x7 && ~x8 )
						nx_state = s1237;
					else nx_state = s1237;
				s1238 : if( x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s21;
						end
					else if( ~x5 && x6 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s1499;
						end
					else if( ~x5 && ~x6 && x2 && x18 && x19 && x4 && x3 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y21 = 1'b1;	
							y32 = 1'b1;	y35 = 1'b1;	
							nx_state = s1500;
						end
					else if( ~x5 && ~x6 && x2 && x18 && x19 && x4 && ~x3 && x17 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x5 && ~x6 && x2 && x18 && x19 && x4 && ~x3 && ~x17 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x5 && ~x6 && x2 && x18 && x19 && x4 && ~x3 && ~x17 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x5 && ~x6 && x2 && x18 && x19 && x4 && ~x3 && ~x17 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x5 && ~x6 && x2 && x18 && x19 && x4 && ~x3 && ~x17 && ~x11 )
						nx_state = s1;
					else if( ~x5 && ~x6 && x2 && x18 && x19 && ~x4 && x3 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y19 = 1'b1;	
							nx_state = s872;
						end
					else if( ~x5 && ~x6 && x2 && x18 && x19 && ~x4 && ~x3 && x16 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x5 && ~x6 && x2 && x18 && x19 && ~x4 && ~x3 && ~x16 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x5 && ~x6 && x2 && x18 && x19 && ~x4 && ~x3 && ~x16 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x5 && ~x6 && x2 && x18 && x19 && ~x4 && ~x3 && ~x16 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x5 && ~x6 && x2 && x18 && x19 && ~x4 && ~x3 && ~x16 && ~x11 )
						nx_state = s1;
					else if( ~x5 && ~x6 && x2 && x18 && ~x19 && x3 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x5 && ~x6 && x2 && x18 && ~x19 && x3 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x5 && ~x6 && x2 && x18 && ~x19 && x3 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x5 && ~x6 && x2 && x18 && ~x19 && x3 && ~x11 )
						nx_state = s1;
					else if( ~x5 && ~x6 && x2 && x18 && ~x19 && ~x3 && x4 )
						begin
							y38 = 1'b1;	
							nx_state = s845;
						end
					else if( ~x5 && ~x6 && x2 && x18 && ~x19 && ~x3 && ~x4 )
						begin
							y39 = 1'b1;	
							nx_state = s277;
						end
					else if( ~x5 && ~x6 && x2 && ~x18 && x19 && x4 && x3 )
						begin
							y44 = 1'b1;	
							nx_state = s1138;
						end
					else if( ~x5 && ~x6 && x2 && ~x18 && x19 && x4 && ~x3 )
						begin
							y47 = 1'b1;	
							nx_state = s675;
						end
					else if( ~x5 && ~x6 && x2 && ~x18 && x19 && ~x4 && x3 )
						begin
							y45 = 1'b1;	
							nx_state = s286;
						end
					else if( ~x5 && ~x6 && x2 && ~x18 && x19 && ~x4 && ~x3 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s1501;
						end
					else if( ~x5 && ~x6 && x2 && ~x18 && ~x19 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y31 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x5 && ~x6 && ~x2 && x18 && x4 && x19 && x3 && x15 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x5 && ~x6 && ~x2 && x18 && x4 && x19 && x3 && ~x15 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x5 && ~x6 && ~x2 && x18 && x4 && x19 && x3 && ~x15 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x5 && ~x6 && ~x2 && x18 && x4 && x19 && x3 && ~x15 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x5 && ~x6 && ~x2 && x18 && x4 && x19 && x3 && ~x15 && ~x11 )
						nx_state = s1;
					else if( ~x5 && ~x6 && ~x2 && x18 && x4 && x19 && ~x3 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x5 && ~x6 && ~x2 && x18 && x4 && ~x19 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x5 && ~x6 && ~x2 && x18 && x4 && ~x19 && ~x3 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							y42 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x5 && ~x6 && ~x2 && x18 && ~x4 && x19 && x3 && x14 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x5 && ~x6 && ~x2 && x18 && ~x4 && x19 && x3 && ~x14 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x5 && ~x6 && ~x2 && x18 && ~x4 && x19 && x3 && ~x14 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x5 && ~x6 && ~x2 && x18 && ~x4 && x19 && x3 && ~x14 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x5 && ~x6 && ~x2 && x18 && ~x4 && x19 && x3 && ~x14 && ~x11 )
						nx_state = s1;
					else if( ~x5 && ~x6 && ~x2 && x18 && ~x4 && x19 && ~x3 )
						begin
							y47 = 1'b1;	
							nx_state = s287;
						end
					else if( ~x5 && ~x6 && ~x2 && x18 && ~x4 && ~x19 && x3 && x12 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x5 && ~x6 && ~x2 && x18 && ~x4 && ~x19 && x3 && ~x12 && x11 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x5 && ~x6 && ~x2 && x18 && ~x4 && ~x19 && x3 && ~x12 && x11 && ~x13 )
						nx_state = s1;
					else if( ~x5 && ~x6 && ~x2 && x18 && ~x4 && ~x19 && x3 && ~x12 && ~x11 )
						nx_state = s1;
					else if( ~x5 && ~x6 && ~x2 && x18 && ~x4 && ~x19 && ~x3 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x5 && ~x6 && ~x2 && ~x18 && x19 && x4 && x3 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x5 && ~x6 && ~x2 && ~x18 && x19 && x4 && ~x3 )
						begin
							y37 = 1'b1;	
							nx_state = s1173;
						end
					else if( ~x5 && ~x6 && ~x2 && ~x18 && x19 && ~x4 && x3 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x5 && ~x6 && ~x2 && ~x18 && x19 && ~x4 && ~x3 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s1502;
						end
					else if( ~x5 && ~x6 && ~x2 && ~x18 && ~x19 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							y31 = 1'b1;	y34 = 1'b1;	
							nx_state = s820;
						end
					else nx_state = s1238;
				s1239 : if( 1'b1 )
						begin
							y2 = 1'b1;	
							nx_state = s1111;
						end
					else nx_state = s1239;
				s1240 : if( x3 )
						begin
							y38 = 1'b1;	
							nx_state = s1503;
						end
					else if( ~x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y14 = 1'b1;	y43 = 1'b1;	
							nx_state = s1504;
						end
					else nx_state = s1240;
				s1241 : if( 1'b1 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s1495;
						end
					else nx_state = s1241;
				s1242 : if( 1'b1 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y58 = 1'b1;	
							nx_state = s1505;
						end
					else nx_state = s1242;
				s1243 : if( 1'b1 )
						begin
							y6 = 1'b1;	
							nx_state = s1506;
						end
					else nx_state = s1243;
				s1244 : if( 1'b1 )
						begin
							y32 = 1'b1;	
							nx_state = s1507;
						end
					else nx_state = s1244;
				s1245 : if( 1'b1 )
						begin
							y58 = 1'b1;	
							nx_state = s1508;
						end
					else nx_state = s1245;
				s1246 : if( 1'b1 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s1246;
				s1247 : if( x4 && x3 )
						begin
							y26 = 1'b1;	
							nx_state = s1468;
						end
					else if( x4 && ~x3 && x5 && x15 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s654;
						end
					else if( x4 && ~x3 && x5 && ~x15 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x4 && ~x3 && x5 && ~x15 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x4 && ~x3 && x5 && ~x15 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( x4 && ~x3 && x5 && ~x15 && ~x22 )
						nx_state = s1;
					else if( x4 && ~x3 && ~x5 && x17 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s654;
						end
					else if( x4 && ~x3 && ~x5 && ~x17 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x4 && ~x3 && ~x5 && ~x17 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x4 && ~x3 && ~x5 && ~x17 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( x4 && ~x3 && ~x5 && ~x17 && ~x22 )
						nx_state = s1;
					else if( ~x4 && x5 && x3 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1509;
						end
					else if( ~x4 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x4 && ~x5 && x3 && x16 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x4 && ~x5 && x3 && ~x16 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x4 && ~x5 && x3 && ~x16 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x4 && ~x5 && x3 && ~x16 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( ~x4 && ~x5 && x3 && ~x16 && ~x22 )
						nx_state = s1;
					else if( ~x4 && ~x5 && ~x3 )
						begin
							y38 = 1'b1;	
							nx_state = s845;
						end
					else nx_state = s1247;
				s1248 : if( x1 && x4 && x5 )
						begin
							y26 = 1'b1;	
							nx_state = s1197;
						end
					else if( x1 && x4 && ~x5 && x3 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( x1 && x4 && ~x5 && ~x3 && x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s653;
						end
					else if( x1 && x4 && ~x5 && ~x3 && ~x6 && x7 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s653;
						end
					else if( x1 && x4 && ~x5 && ~x3 && ~x6 && ~x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s654;
						end
					else if( x1 && ~x4 )
						begin
							y26 = 1'b1;	
							nx_state = s1197;
						end
					else if( ~x1 )
						begin
							y26 = 1'b1;	
							nx_state = s1197;
						end
					else nx_state = s1248;
				s1249 : if( x64 && x63 && x4 && x5 && x3 )
						begin
							y41 = 1'b1;	y45 = 1'b1;	y46 = 1'b1;	
							nx_state = s654;
						end
					else if( x64 && x63 && x4 && x5 && ~x3 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y47 = 1'b1;	y48 = 1'b1;	
							nx_state = s654;
						end
					else if( x64 && x63 && x4 && ~x5 && x3 )
						begin
							y39 = 1'b1;	y43 = 1'b1;	y44 = 1'b1;	
							nx_state = s654;
						end
					else if( x64 && x63 && x4 && ~x5 && ~x3 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y48 = 1'b1;	y49 = 1'b1;	
							nx_state = s654;
						end
					else if( x64 && x63 && ~x4 && x3 && x5 )
						begin
							y41 = 1'b1;	y42 = 1'b1;	
							nx_state = s654;
						end
					else if( x64 && x63 && ~x4 && x3 && ~x5 )
						begin
							y39 = 1'b1;	y40 = 1'b1;	
							nx_state = s654;
						end
					else if( x64 && x63 && ~x4 && ~x3 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y32 = 1'b1;	y48 = 1'b1;	
							nx_state = s654;
						end
					else if( x64 && ~x63 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x64 && x63 && x66 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s1051;
						end
					else if( ~x64 && x63 && ~x66 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s1510;
						end
					else if( ~x64 && ~x63 && x65 )
						begin
							y5 = 1'b1;	y42 = 1'b1;	y43 = 1'b1;	
							y68 = 1'b1;	
							nx_state = s889;
						end
					else if( ~x64 && ~x63 && ~x65 && x67 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x64 && ~x63 && ~x65 && ~x67 )
						begin
							y6 = 1'b1;	
							nx_state = s239;
						end
					else nx_state = s1249;
				s1250 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y12 = 1'b1;	
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s1511;
						end
					else nx_state = s1250;
				s1251 : if( 1'b1 )
						begin
							y6 = 1'b1;	y9 = 1'b1;	y25 = 1'b1;	
							y56 = 1'b1;	
							nx_state = s1512;
						end
					else nx_state = s1251;
				s1252 : if( x16 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x16 && ~x15 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x16 )
						begin
							y35 = 1'b1;	
							nx_state = s718;
						end
					else nx_state = s1252;
				s1253 : if( x15 )
						begin
							y34 = 1'b1;	
							nx_state = s1165;
						end
					else if( ~x15 )
						begin
							y35 = 1'b1;	
							nx_state = s718;
						end
					else nx_state = s1253;
				s1254 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s948;
						end
					else nx_state = s1254;
				s1255 : if( 1'b1 )
						begin
							y47 = 1'b1;	y55 = 1'b1;	y61 = 1'b1;	
							y71 = 1'b1;	
							nx_state = s1513;
						end
					else nx_state = s1255;
				s1256 : if( 1'b1 )
						begin
							y47 = 1'b1;	y56 = 1'b1;	y61 = 1'b1;	
							y70 = 1'b1;	
							nx_state = s1514;
						end
					else nx_state = s1256;
				s1257 : if( 1'b1 )
						begin
							y47 = 1'b1;	y55 = 1'b1;	y61 = 1'b1;	
							y68 = 1'b1;	
							nx_state = s1515;
						end
					else nx_state = s1257;
				s1258 : if( 1'b1 )
						begin
							y2 = 1'b1;	y37 = 1'b1;	y39 = 1'b1;	
							nx_state = s720;
						end
					else nx_state = s1258;
				s1259 : if( x20 && x21 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x20 && x21 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x20 && x21 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x20 && x21 && ~x10 )
						nx_state = s1;
					else if( x20 && ~x21 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y22 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1516;
						end
					else if( ~x20 && x21 )
						begin
							y22 = 1'b1;	
							nx_state = s1121;
						end
					else if( ~x20 && ~x21 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && ~x21 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && ~x21 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x20 && ~x21 && ~x10 )
						nx_state = s1;
					else nx_state = s1259;
				s1260 : if( 1'b1 )
						begin
							y22 = 1'b1;	y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s1024;
						end
					else nx_state = s1260;
				s1261 : if( x64 && x20 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1016;
						end
					else if( x64 && ~x20 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s1014;
						end
					else if( ~x64 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s822;
						end
					else if( ~x64 && ~x11 )
						begin
							y68 = 1'b1;	
							nx_state = s1404;
						end
					else nx_state = s1261;
				s1262 : if( x64 && x66 )
						begin
							y18 = 1'b1;	y27 = 1'b1;	y29 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s1517;
						end
					else if( x64 && ~x66 )
						begin
							y25 = 1'b1;	
							nx_state = s1010;
						end
					else if( ~x64 && x14 && x31 && x30 )
						begin
							y3 = 1'b1;	
							nx_state = s788;
						end
					else if( ~x64 && x14 && x31 && ~x30 )
						begin
							y3 = 1'b1;	
							nx_state = s1293;
						end
					else if( ~x64 && x14 && ~x31 && x30 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( ~x64 && x14 && ~x31 && ~x30 )
						begin
							y3 = 1'b1;	
							nx_state = s789;
						end
					else if( ~x64 && ~x14 )
						begin
							y25 = 1'b1;	
							nx_state = s838;
						end
					else nx_state = s1262;
				s1263 : if( x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x10 && ~x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x10 )
						nx_state = s1;
					else nx_state = s1263;
				s1264 : if( x21 && x9 )
						begin
							y44 = 1'b1;	
							nx_state = s755;
						end
					else if( x21 && ~x9 )
						begin
							y44 = 1'b1;	
							nx_state = s1138;
						end
					else if( ~x21 && x5 && x8 && x7 )
						begin
							y44 = 1'b1;	
							nx_state = s755;
						end
					else if( ~x21 && x5 && x8 && ~x7 && x9 && x18 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1263;
						end
					else if( ~x21 && x5 && x8 && ~x7 && x9 && ~x18 && x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x21 && x5 && x8 && ~x7 && x9 && ~x18 && x10 && ~x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x21 && x5 && x8 && ~x7 && x9 && ~x18 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x21 && x5 && x8 && ~x7 && x9 && ~x18 && ~x10 )
						nx_state = s1;
					else if( ~x21 && x5 && x8 && ~x7 && ~x9 && x19 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1263;
						end
					else if( ~x21 && x5 && x8 && ~x7 && ~x9 && ~x19 && x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x21 && x5 && x8 && ~x7 && ~x9 && ~x19 && x10 && ~x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x21 && x5 && x8 && ~x7 && ~x9 && ~x19 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x21 && x5 && x8 && ~x7 && ~x9 && ~x19 && ~x10 )
						nx_state = s1;
					else if( ~x21 && x5 && ~x8 && x7 && x9 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else if( ~x21 && x5 && ~x8 && x7 && ~x9 && x20 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1263;
						end
					else if( ~x21 && x5 && ~x8 && x7 && ~x9 && ~x20 && x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x21 && x5 && ~x8 && x7 && ~x9 && ~x20 && x10 && ~x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x21 && x5 && ~x8 && x7 && ~x9 && ~x20 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x21 && x5 && ~x8 && x7 && ~x9 && ~x20 && ~x10 )
						nx_state = s1;
					else if( ~x21 && x5 && ~x8 && ~x7 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1263;
						end
					else if( ~x21 && ~x5 )
						begin
							y44 = 1'b1;	
							nx_state = s755;
						end
					else nx_state = s1264;
				s1265 : if( x63 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y36 = 1'b1;	
							y59 = 1'b1;	
							nx_state = s741;
						end
					else if( ~x63 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s1518;
						end
					else nx_state = s1265;
				s1266 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y36 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s1519;
						end
					else nx_state = s1266;
				s1267 : if( x9 && x8 && x10 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y5 = 1'b1;	
							y22 = 1'b1;	y23 = 1'b1;	
							nx_state = s72;
						end
					else if( x9 && x8 && ~x10 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else if( x9 && ~x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x9 && x10 && x8 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x9 && x10 && x8 && ~x13 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x9 && x10 && x8 && ~x13 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x9 && x10 && x8 && ~x13 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x9 && x10 && x8 && ~x13 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x9 && x10 && x8 && ~x13 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x9 && x10 && ~x8 && x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x9 && x10 && ~x8 && ~x3 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x9 && x10 && ~x8 && ~x3 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x9 && x10 && ~x8 && ~x3 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x9 && x10 && ~x8 && ~x3 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x9 && x10 && ~x8 && ~x3 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x9 && ~x10 && x8 && x1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x9 && ~x10 && x8 && ~x1 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x9 && ~x10 && x8 && ~x1 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x9 && ~x10 && x8 && ~x1 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x9 && ~x10 && x8 && ~x1 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x9 && ~x10 && x8 && ~x1 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x9 && ~x10 && ~x8 && x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s522;
						end
					else if( ~x9 && ~x10 && ~x8 && ~x15 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x9 && ~x10 && ~x8 && ~x15 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x9 && ~x10 && ~x8 && ~x15 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x9 && ~x10 && ~x8 && ~x15 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x9 && ~x10 && ~x8 && ~x15 && ~x6 && ~x5 )
						nx_state = s1;
					else nx_state = s1267;
				s1268 : if( x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s1269;
						end
					else if( ~x16 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s1270;
						end
					else nx_state = s1268;
				s1269 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s1270;
						end
					else nx_state = s1269;
				s1270 : if( x67 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s1520;
						end
					else if( ~x67 )
						begin
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s1357;
						end
					else nx_state = s1270;
				s1271 : if( 1'b1 )
						begin
							y26 = 1'b1;	
							nx_state = s1468;
						end
					else nx_state = s1271;
				s1272 : if( x65 )
						begin
							y8 = 1'b1;	
							nx_state = s785;
						end
					else if( ~x65 )
						begin
							y7 = 1'b1;	
							nx_state = s985;
						end
					else nx_state = s1272;
				s1273 : if( 1'b1 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s1521;
						end
					else nx_state = s1273;
				s1274 : if( 1'b1 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s1522;
						end
					else nx_state = s1274;
				s1275 : if( 1'b1 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s1523;
						end
					else nx_state = s1275;
				s1276 : if( 1'b1 )
						begin
							y24 = 1'b1;	
							nx_state = s259;
						end
					else nx_state = s1276;
				s1277 : if( 1'b1 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y27 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s749;
						end
					else nx_state = s1277;
				s1278 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s1524;
						end
					else nx_state = s1278;
				s1279 : if( x15 && x5 )
						begin
							y44 = 1'b1;	y48 = 1'b1;	y49 = 1'b1;	
							nx_state = s1525;
						end
					else if( x15 && ~x5 && x21 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y27 = 1'b1;	
							y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s1263;
						end
					else if( x15 && ~x5 && ~x21 && x8 && x9 )
						begin
							y6 = 1'b1;	y30 = 1'b1;	y31 = 1'b1;	
							y32 = 1'b1;	y38 = 1'b1;	
							nx_state = s1263;
						end
					else if( x15 && ~x5 && ~x21 && x8 && ~x9 )
						begin
							y6 = 1'b1;	y30 = 1'b1;	y31 = 1'b1;	
							y32 = 1'b1;	y38 = 1'b1;	
							nx_state = s1263;
						end
					else if( x15 && ~x5 && ~x21 && ~x8 )
						begin
							y6 = 1'b1;	y30 = 1'b1;	y31 = 1'b1;	
							y32 = 1'b1;	y38 = 1'b1;	
							nx_state = s1263;
						end
					else if( ~x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	y46 = 1'b1;	
							nx_state = s1526;
						end
					else nx_state = s1279;
				s1280 : if( x15 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s770;
						end
					else if( ~x15 && x3 && x2 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s764;
						end
					else if( ~x15 && x3 && ~x2 )
						nx_state = s1280;
					else if( ~x15 && ~x3 && x4 && x2 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s1284;
						end
					else if( ~x15 && ~x3 && x4 && ~x2 )
						nx_state = s1280;
					else if( ~x15 && ~x3 && ~x4 && x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s761;
						end
					else if( ~x15 && ~x3 && ~x4 && ~x2 )
						nx_state = s1280;
					else nx_state = s1280;
				s1281 : if( x62 && x17 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							nx_state = s1527;
						end
					else if( x62 && ~x17 )
						begin
							y1 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1300;
						end
					else if( ~x62 )
						begin
							y13 = 1'b1;	
							nx_state = s1528;
						end
					else nx_state = s1281;
				s1282 : if( x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s216;
						end
					else if( ~x15 && x13 && x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s1284;
						end
					else if( ~x15 && x13 && ~x4 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s761;
						end
					else if( ~x15 && ~x13 && x14 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s764;
						end
					else if( ~x15 && ~x13 && ~x14 && x9 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s764;
						end
					else if( ~x15 && ~x13 && ~x14 && ~x9 && x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s764;
						end
					else if( ~x15 && ~x13 && ~x14 && ~x9 && ~x7 && x8 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s764;
						end
					else if( ~x15 && ~x13 && ~x14 && ~x9 && ~x7 && ~x8 )
						nx_state = s1282;
					else nx_state = s1282;
				s1283 : if( x15 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	
							nx_state = s1233;
						end
					else if( ~x15 && x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s817;
						end
					else if( ~x15 && ~x12 )
						nx_state = s1283;
					else nx_state = s1283;
				s1284 : if( x15 )
						begin
							y2 = 1'b1;	
							nx_state = s768;
						end
					else if( ~x15 && x6 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x15 && ~x6 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s770;
						end
					else nx_state = s1284;
				s1285 : if( 1'b1 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else nx_state = s1285;
				s1286 : if( x7 && x19 && x18 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x7 && x19 && x18 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x7 && x19 && x18 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x7 && x19 && x18 && ~x11 )
						nx_state = s1;
					else if( x7 && x19 && ~x18 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y20 = 1'b1;	
							nx_state = s820;
						end
					else if( x7 && ~x19 && x2 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x7 && ~x19 && x2 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x7 && ~x19 && x2 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x7 && ~x19 && x2 && ~x11 )
						nx_state = s1;
					else if( x7 && ~x19 && ~x2 && x18 && x3 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x7 && ~x19 && ~x2 && x18 && x3 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x7 && ~x19 && ~x2 && x18 && x3 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x7 && ~x19 && ~x2 && x18 && x3 && ~x11 )
						nx_state = s1;
					else if( x7 && ~x19 && ~x2 && x18 && ~x3 && x4 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	y20 = 1'b1;	
							y42 = 1'b1;	
							nx_state = s820;
						end
					else if( x7 && ~x19 && ~x2 && x18 && ~x3 && ~x4 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x7 && ~x19 && ~x2 && x18 && ~x3 && ~x4 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x7 && ~x19 && ~x2 && x18 && ~x3 && ~x4 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x7 && ~x19 && ~x2 && x18 && ~x3 && ~x4 && ~x11 )
						nx_state = s1;
					else if( x7 && ~x19 && ~x2 && ~x18 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y20 = 1'b1;	
							y31 = 1'b1;	y34 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x7 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y20 = 1'b1;	
							nx_state = s1529;
						end
					else nx_state = s1286;
				s1287 : if( x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1430;
						end
					else if( ~x3 )
						begin
							y14 = 1'b1;	y37 = 1'b1;	y43 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s1530;
						end
					else nx_state = s1287;
				s1288 : if( x18 && x22 && x23 && x4 && x3 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x18 && x22 && x23 && x4 && x3 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x18 && x22 && x23 && x4 && x3 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( x18 && x22 && x23 && x4 && x3 && ~x21 )
						nx_state = s1;
					else if( x18 && x22 && x23 && x4 && ~x3 && x5 && x15 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x18 && x22 && x23 && x4 && ~x3 && x5 && ~x15 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x18 && x22 && x23 && x4 && ~x3 && x5 && ~x15 && x21 && ~x16 )
						nx_state = s1;
					else if( x18 && x22 && x23 && x4 && ~x3 && x5 && ~x15 && ~x21 )
						nx_state = s1;
					else if( x18 && x22 && x23 && x4 && ~x3 && ~x5 && x16 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x18 && x22 && x23 && x4 && ~x3 && ~x5 && ~x16 && x21 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x18 && x22 && x23 && x4 && ~x3 && ~x5 && ~x16 && x21 && ~x15 )
						nx_state = s1;
					else if( x18 && x22 && x23 && x4 && ~x3 && ~x5 && ~x16 && ~x21 )
						nx_state = s1;
					else if( x18 && x22 && x23 && ~x4 && x5 && x3 )
						begin
							y25 = 1'b1;	y26 = 1'b1;	
							nx_state = s1;
						end
					else if( x18 && x22 && x23 && ~x4 && x5 && ~x3 )
						begin
							y1 = 1'b1;	y20 = 1'b1;	y47 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s535;
						end
					else if( x18 && x22 && x23 && ~x4 && ~x5 && x3 )
						begin
							y51 = 1'b1;	y52 = 1'b1;	
							nx_state = s1;
						end
					else if( x18 && x22 && x23 && ~x4 && ~x5 && ~x3 )
						begin
							y1 = 1'b1;	y19 = 1'b1;	y49 = 1'b1;	
							y50 = 1'b1;	
							nx_state = s535;
						end
					else if( x18 && x22 && ~x23 && x9 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y36 = 1'b1;	
							nx_state = s535;
						end
					else if( x18 && x22 && ~x23 && ~x9 && x3 && x5 && x4 )
						begin
							y42 = 1'b1;	
							nx_state = s754;
						end
					else if( x18 && x22 && ~x23 && ~x9 && x3 && x5 && ~x4 )
						begin
							y40 = 1'b1;	
							nx_state = s751;
						end
					else if( x18 && x22 && ~x23 && ~x9 && x3 && ~x5 && x4 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x18 && x22 && ~x23 && ~x9 && x3 && ~x5 && ~x4 )
						begin
							y39 = 1'b1;	
							nx_state = s277;
						end
					else if( x18 && x22 && ~x23 && ~x9 && ~x3 && x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y11 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s535;
						end
					else if( x18 && x22 && ~x23 && ~x9 && ~x3 && ~x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y8 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s1531;
						end
					else if( x18 && ~x22 && x23 && x9 )
						begin
							y46 = 1'b1;	
							nx_state = s1030;
						end
					else if( x18 && ~x22 && x23 && ~x9 && x10 && x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y11 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s1532;
						end
					else if( x18 && ~x22 && x23 && ~x9 && x10 && ~x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y8 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s1531;
						end
					else if( x18 && ~x22 && x23 && ~x9 && ~x10 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y8 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s1531;
						end
					else if( x18 && ~x22 && ~x23 && x3 && x5 && x4 )
						begin
							y31 = 1'b1;	y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s535;
						end
					else if( x18 && ~x22 && ~x23 && x3 && x5 && ~x4 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x18 && ~x22 && ~x23 && x3 && ~x5 && x4 )
						begin
							y30 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							nx_state = s535;
						end
					else if( x18 && ~x22 && ~x23 && x3 && ~x5 && ~x4 )
						begin
							y30 = 1'b1;	
							nx_state = s291;
						end
					else if( x18 && ~x22 && ~x23 && ~x3 && x8 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	y44 = 1'b1;	
							nx_state = s535;
						end
					else if( x18 && ~x22 && ~x23 && ~x3 && ~x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y8 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s1531;
						end
					else if( ~x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y11 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s1533;
						end
					else nx_state = s1288;
				s1289 : if( 1'b1 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s1534;
						end
					else nx_state = s1289;
				s1290 : if( x11 && x19 && x20 && x2 && x1 && x4 && x3 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x11 && x19 && x20 && x2 && x1 && x4 && x3 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x11 && x19 && x20 && x2 && x1 && x4 && x3 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( x11 && x19 && x20 && x2 && x1 && x4 && x3 && ~x22 )
						nx_state = s1;
					else if( x11 && x19 && x20 && x2 && x1 && x4 && ~x3 && x5 && x18 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x11 && x19 && x20 && x2 && x1 && x4 && ~x3 && x5 && ~x18 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x11 && x19 && x20 && x2 && x1 && x4 && ~x3 && x5 && ~x18 && x22 && ~x21 )
						nx_state = s1;
					else if( x11 && x19 && x20 && x2 && x1 && x4 && ~x3 && x5 && ~x18 && ~x22 )
						nx_state = s1;
					else if( x11 && x19 && x20 && x2 && x1 && x4 && ~x3 && ~x5 && x21 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x11 && x19 && x20 && x2 && x1 && x4 && ~x3 && ~x5 && ~x21 && x22 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x11 && x19 && x20 && x2 && x1 && x4 && ~x3 && ~x5 && ~x21 && x22 && ~x18 )
						nx_state = s1;
					else if( x11 && x19 && x20 && x2 && x1 && x4 && ~x3 && ~x5 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x11 && x19 && x20 && x2 && x1 && ~x4 && x5 && x3 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x11 && x19 && x20 && x2 && x1 && ~x4 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	y36 = 1'b1;	
							nx_state = s654;
						end
					else if( x11 && x19 && x20 && x2 && x1 && ~x4 && ~x5 && x3 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x11 && x19 && x20 && x2 && x1 && ~x4 && ~x5 && ~x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y34 = 1'b1;	y37 = 1'b1;	
							nx_state = s654;
						end
					else if( x11 && x19 && x20 && x2 && ~x1 )
						begin
							y26 = 1'b1;	
							nx_state = s413;
						end
					else if( x11 && x19 && x20 && ~x2 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s715;
						end
					else if( x11 && x19 && x20 && ~x2 && ~x8 )
						begin
							y26 = 1'b1;	
							nx_state = s413;
						end
					else if( x11 && x19 && ~x20 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s716;
						end
					else if( x11 && ~x19 )
						begin
							y28 = 1'b1;	
							nx_state = s717;
						end
					else if( ~x11 )
						begin
							y29 = 1'b1;	
							nx_state = s771;
						end
					else nx_state = s1290;
				s1291 : if( 1'b1 )
						begin
							y55 = 1'b1;	
							nx_state = s282;
						end
					else nx_state = s1291;
				s1292 : if( x21 && x20 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( x21 && ~x20 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else if( ~x21 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s58;
						end
					else nx_state = s1292;
				s1293 : if( x64 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s591;
						end
					else if( ~x64 && x30 )
						begin
							y47 = 1'b1;	y52 = 1'b1;	y61 = 1'b1;	
							y66 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x64 && ~x30 )
						begin
							y47 = 1'b1;	y50 = 1'b1;	y61 = 1'b1;	
							y65 = 1'b1;	
							nx_state = s1148;
						end
					else nx_state = s1293;
				s1294 : if( 1'b1 )
						begin
							y6 = 1'b1;	
							nx_state = s239;
						end
					else nx_state = s1294;
				s1295 : if( x64 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1535;
						end
					else if( ~x64 )
						begin
							y48 = 1'b1;	y55 = 1'b1;	y61 = 1'b1;	
							nx_state = s1536;
						end
					else nx_state = s1295;
				s1296 : if( 1'b1 )
						begin
							y6 = 1'b1;	
							nx_state = s659;
						end
					else nx_state = s1296;
				s1297 : if( 1'b1 )
						begin
							y39 = 1'b1;	
							nx_state = s1537;
						end
					else nx_state = s1297;
				s1298 : if( x14 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x14 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x14 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x14 && ~x23 )
						nx_state = s1;
					else if( ~x14 )
						begin
							y39 = 1'b1;	
							nx_state = s277;
						end
					else nx_state = s1298;
				s1299 : if( 1'b1 )
						begin
							y9 = 1'b1;	
							nx_state = s892;
						end
					else nx_state = s1299;
				s1300 : if( 1'b1 )
						begin
							y13 = 1'b1;	
							nx_state = s1281;
						end
					else nx_state = s1300;
				s1301 : if( 1'b1 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1131;
						end
					else nx_state = s1301;
				s1302 : if( 1'b1 )
						begin
							y37 = 1'b1;	
							nx_state = s1173;
						end
					else nx_state = s1302;
				s1303 : if( 1'b1 )
						begin
							y22 = 1'b1;	
							nx_state = s823;
						end
					else nx_state = s1303;
				s1304 : if( 1'b1 )
						begin
							y8 = 1'b1;	
							nx_state = s568;
						end
					else nx_state = s1304;
				s1305 : if( x21 && x18 && x13 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( x21 && x18 && ~x13 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else if( x21 && ~x18 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x21 && x22 && x18 && x19 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x21 && x22 && x18 && ~x19 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x21 && x22 && ~x18 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x21 && ~x22 && x19 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x21 && ~x22 && ~x19 && x13 && x20 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x21 && ~x22 && ~x19 && x13 && ~x20 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x21 && ~x22 && ~x19 && ~x13 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s1305;
				s1306 : if( 1'b1 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1094;
						end
					else nx_state = s1306;
				s1307 : if( 1'b1 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else nx_state = s1307;
				s1308 : if( x4 && x22 && x30 && x9 && x10 && x8 )
						begin
							y11 = 1'b1;	
							nx_state = s34;
						end
					else if( x4 && x22 && x30 && x9 && x10 && ~x8 )
						begin
							y8 = 1'b1;	
							nx_state = s784;
						end
					else if( x4 && x22 && x30 && x9 && ~x10 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x4 && x22 && x30 && x9 && ~x10 && ~x8 )
						begin
							y8 = 1'b1;	
							nx_state = s785;
						end
					else if( x4 && x22 && x30 && ~x9 && x10 && x8 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( x4 && x22 && x30 && ~x9 && x10 && ~x8 && x27 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( x4 && x22 && x30 && ~x9 && x10 && ~x8 && ~x27 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else if( x4 && x22 && x30 && ~x9 && ~x10 && x8 )
						begin
							y8 = 1'b1;	
							nx_state = s786;
						end
					else if( x4 && x22 && x30 && ~x9 && ~x10 && ~x8 && x26 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x4 && x22 && x30 && ~x9 && ~x10 && ~x8 && ~x26 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( x4 && x22 && ~x30 && x31 && x9 && x10 && x8 )
						begin
							y9 = 1'b1;	
							nx_state = s790;
						end
					else if( x4 && x22 && ~x30 && x31 && x9 && x10 && ~x8 && x21 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( x4 && x22 && ~x30 && x31 && x9 && x10 && ~x8 && ~x21 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x4 && x22 && ~x30 && x31 && x9 && x10 && ~x8 && ~x21 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x4 && x22 && ~x30 && x31 && x9 && x10 && ~x8 && ~x21 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x4 && x22 && ~x30 && x31 && x9 && x10 && ~x8 && ~x21 && ~x23 )
						nx_state = s1;
					else if( x4 && x22 && ~x30 && x31 && x9 && ~x10 && x8 )
						begin
							y3 = 1'b1;	
							nx_state = s789;
						end
					else if( x4 && x22 && ~x30 && x31 && x9 && ~x10 && ~x8 && x18 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( x4 && x22 && ~x30 && x31 && x9 && ~x10 && ~x8 && ~x18 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x4 && x22 && ~x30 && x31 && x9 && ~x10 && ~x8 && ~x18 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x4 && x22 && ~x30 && x31 && x9 && ~x10 && ~x8 && ~x18 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x4 && x22 && ~x30 && x31 && x9 && ~x10 && ~x8 && ~x18 && ~x23 )
						nx_state = s1;
					else if( x4 && x22 && ~x30 && x31 && ~x9 && x8 && x10 && x19 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( x4 && x22 && ~x30 && x31 && ~x9 && x8 && x10 && ~x19 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x4 && x22 && ~x30 && x31 && ~x9 && x8 && x10 && ~x19 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x4 && x22 && ~x30 && x31 && ~x9 && x8 && x10 && ~x19 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x4 && x22 && ~x30 && x31 && ~x9 && x8 && x10 && ~x19 && ~x23 )
						nx_state = s1;
					else if( x4 && x22 && ~x30 && x31 && ~x9 && x8 && ~x10 && x20 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( x4 && x22 && ~x30 && x31 && ~x9 && x8 && ~x10 && ~x20 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x4 && x22 && ~x30 && x31 && ~x9 && x8 && ~x10 && ~x20 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x4 && x22 && ~x30 && x31 && ~x9 && x8 && ~x10 && ~x20 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x4 && x22 && ~x30 && x31 && ~x9 && x8 && ~x10 && ~x20 && ~x23 )
						nx_state = s1;
					else if( x4 && x22 && ~x30 && x31 && ~x9 && ~x8 )
						begin
							y3 = 1'b1;	
							nx_state = s711;
						end
					else if( x4 && x22 && ~x30 && ~x31 )
						begin
							y9 = 1'b1;	
							nx_state = s790;
						end
					else if( x4 && ~x22 )
						begin
							y45 = 1'b1;	y47 = 1'b1;	y50 = 1'b1;	
							y60 = 1'b1;	y62 = 1'b1;	y64 = 1'b1;	
							nx_state = s787;
						end
					else if( ~x4 && x30 )
						begin
							y37 = 1'b1;	
							nx_state = s1356;
						end
					else if( ~x4 && ~x30 && x31 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x4 && ~x30 && ~x31 )
						begin
							y37 = 1'b1;	
							nx_state = s1173;
						end
					else nx_state = s1308;
				s1309 : if( x3 && x4 && x6 )
						begin
							y39 = 1'b1;	
							nx_state = s1295;
						end
					else if( x3 && x4 && ~x6 )
						begin
							y39 = 1'b1;	
							nx_state = s1537;
						end
					else if( x3 && ~x4 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1538;
						end
					else if( ~x3 && x5 )
						begin
							y6 = 1'b1;	y26 = 1'b1;	
							nx_state = s815;
						end
					else if( ~x3 && ~x5 )
						begin
							y20 = 1'b1;	
							nx_state = s95;
						end
					else nx_state = s1309;
				s1310 : if( x63 && x2 && x3 && x4 && x9 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x63 && x2 && x3 && x4 && x9 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x63 && x2 && x3 && x4 && x9 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x63 && x2 && x3 && x4 && x9 && ~x1 )
						nx_state = s1;
					else if( x63 && x2 && x3 && x4 && ~x9 && x8 )
						begin
							y45 = 1'b1;	
							nx_state = s286;
						end
					else if( x63 && x2 && x3 && x4 && ~x9 && ~x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x63 && x2 && x3 && ~x4 && x9 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s602;
						end
					else if( x63 && x2 && x3 && ~x4 && x9 && ~x6 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x63 && x2 && x3 && ~x4 && ~x9 && x8 )
						begin
							y44 = 1'b1;	
							nx_state = s1138;
						end
					else if( x63 && x2 && x3 && ~x4 && ~x9 && ~x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x63 && x2 && ~x3 && x4 && x9 )
						begin
							y3 = 1'b1;	y18 = 1'b1;	y21 = 1'b1;	
							nx_state = s1382;
						end
					else if( x63 && x2 && ~x3 && x4 && ~x9 && x8 )
						begin
							y46 = 1'b1;	
							nx_state = s531;
						end
					else if( x63 && x2 && ~x3 && x4 && ~x9 && ~x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x63 && x2 && ~x3 && ~x4 && x9 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( x63 && x2 && ~x3 && ~x4 && x9 && ~x13 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x63 && x2 && ~x3 && ~x4 && x9 && ~x13 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x63 && x2 && ~x3 && ~x4 && x9 && ~x13 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x63 && x2 && ~x3 && ~x4 && x9 && ~x13 && ~x1 )
						nx_state = s1;
					else if( x63 && x2 && ~x3 && ~x4 && ~x9 && x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x63 && x2 && ~x3 && ~x4 && ~x9 && ~x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x63 && ~x2 && x4 && x3 && x9 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( x63 && ~x2 && x4 && x3 && x9 && ~x14 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x63 && ~x2 && x4 && x3 && x9 && ~x14 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x63 && ~x2 && x4 && x3 && x9 && ~x14 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x63 && ~x2 && x4 && x3 && x9 && ~x14 && ~x1 )
						nx_state = s1;
					else if( x63 && ~x2 && x4 && x3 && ~x9 && x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y37 = 1'b1;	
							nx_state = s1540;
						end
					else if( x63 && ~x2 && x4 && x3 && ~x9 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x63 && ~x2 && x4 && ~x3 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( x63 && ~x2 && x4 && ~x3 && ~x9 && x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x63 && ~x2 && x4 && ~x3 && ~x9 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x63 && ~x2 && ~x4 && x9 && x3 && x12 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( x63 && ~x2 && ~x4 && x9 && x3 && ~x12 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x63 && ~x2 && ~x4 && x9 && x3 && ~x12 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x63 && ~x2 && ~x4 && x9 && x3 && ~x12 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x63 && ~x2 && ~x4 && x9 && x3 && ~x12 && ~x1 )
						nx_state = s1;
					else if( x63 && ~x2 && ~x4 && x9 && ~x3 )
						begin
							y26 = 1'b1;	
							nx_state = s1197;
						end
					else if( x63 && ~x2 && ~x4 && ~x9 && x8 && x3 )
						begin
							y3 = 1'b1;	y18 = 1'b1;	y42 = 1'b1;	
							nx_state = s1539;
						end
					else if( x63 && ~x2 && ~x4 && ~x9 && x8 && ~x3 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x63 && ~x2 && ~x4 && ~x9 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x63 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x63 && ~x15 )
						nx_state = s1;
					else nx_state = s1310;
				s1311 : if( 1'b1 )
						begin
							y7 = 1'b1;	
							nx_state = s222;
						end
					else nx_state = s1311;
				s1312 : if( x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y29 = 1'b1;	y36 = 1'b1;	
							nx_state = s1541;
						end
					else if( ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1089;
						end
					else nx_state = s1312;
				s1313 : if( x22 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s1092;
						end
					else if( x22 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1340;
						end
					else if( ~x22 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s1339;
						end
					else if( ~x22 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1089;
						end
					else nx_state = s1313;
				s1314 : if( x21 && x22 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( x21 && ~x22 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( x21 && ~x22 && ~x23 )
						nx_state = s1;
					else if( ~x21 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x21 && ~x23 )
						nx_state = s1;
					else nx_state = s1314;
				s1315 : if( 1'b1 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s604;
						end
					else nx_state = s1315;
				s1316 : if( 1'b1 )
						begin
							y48 = 1'b1;	y53 = 1'b1;	y61 = 1'b1;	
							nx_state = s1536;
						end
					else nx_state = s1316;
				s1317 : if( x63 )
						begin
							y25 = 1'b1;	
							nx_state = s838;
						end
					else if( ~x63 && x66 && x30 )
						begin
							y25 = 1'b1;	
							nx_state = s238;
						end
					else if( ~x63 && x66 && ~x30 )
						begin
							y47 = 1'b1;	y49 = 1'b1;	y58 = 1'b1;	
							y61 = 1'b1;	y68 = 1'b1;	
							nx_state = s831;
						end
					else if( ~x63 && ~x66 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s328;
						end
					else nx_state = s1317;
				s1318 : if( x20 )
						begin
							y8 = 1'b1;	
							nx_state = s568;
						end
					else if( ~x20 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s168;
						end
					else nx_state = s1318;
				s1319 : if( 1'b1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s150;
						end
					else nx_state = s1319;
				s1320 : if( 1'b1 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y21 = 1'b1;	
							nx_state = s820;
						end
					else nx_state = s1320;
				s1321 : if( 1'b1 )
						begin
							y21 = 1'b1;	y29 = 1'b1;	y48 = 1'b1;	
							nx_state = s1542;
						end
					else nx_state = s1321;
				s1322 : if( x15 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	
							nx_state = s1280;
						end
					else if( ~x15 && x3 && x2 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s764;
						end
					else if( ~x15 && x3 && ~x2 )
						nx_state = s1322;
					else if( ~x15 && ~x3 && x4 && x2 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s1284;
						end
					else if( ~x15 && ~x3 && x4 && ~x2 )
						nx_state = s1322;
					else if( ~x15 && ~x3 && ~x4 && x2 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s761;
						end
					else if( ~x15 && ~x3 && ~x4 && ~x2 )
						nx_state = s1322;
					else nx_state = s1322;
				s1323 : if( x20 )
						begin
							y6 = 1'b1;	y11 = 1'b1;	y42 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1028;
						end
					else if( ~x20 )
						begin
							y22 = 1'b1;	
							nx_state = s130;
						end
					else nx_state = s1323;
				s1324 : if( 1'b1 )
						begin
							y2 = 1'b1;	
							nx_state = s768;
						end
					else nx_state = s1324;
				s1325 : if( 1'b1 )
						begin
							y24 = 1'b1;	
							nx_state = s1262;
						end
					else nx_state = s1325;
				s1326 : if( x65 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y14 = 1'b1;	y15 = 1'b1;	y21 = 1'b1;	
							nx_state = s1543;
						end
					else if( ~x65 && x9 )
						begin
							y15 = 1'b1;	
							nx_state = s1544;
						end
					else if( ~x65 && ~x9 && x20 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y45 = 1'b1;	
							y49 = 1'b1;	
							nx_state = s1065;
						end
					else if( ~x65 && ~x9 && ~x20 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1066;
						end
					else nx_state = s1326;
				s1327 : if( x32 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s341;
						end
					else if( ~x32 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x32 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x32 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x32 && ~x10 )
						nx_state = s1;
					else nx_state = s1327;
				s1328 : if( 1'b1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1545;
						end
					else nx_state = s1328;
				s1329 : if( 1'b1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s1044;
						end
					else nx_state = s1329;
				s1330 : if( 1'b1 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s318;
						end
					else nx_state = s1330;
				s1331 : if( x8 && x21 && x16 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x8 && x21 && x16 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s261;
						end
					else if( x8 && x21 && ~x16 && x17 && x18 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s810;
						end
					else if( x8 && x21 && ~x16 && x17 && x18 && ~x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( x8 && x21 && ~x16 && x17 && ~x18 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( x8 && x21 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s252;
						end
					else if( x8 && ~x21 && x22 && x16 && x19 && x18 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( x8 && ~x21 && x22 && x16 && x19 && x18 && ~x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s264;
						end
					else if( x8 && ~x21 && x22 && x16 && x19 && ~x18 && x13 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x8 && ~x21 && x22 && x16 && x19 && ~x18 && ~x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x8 && ~x21 && x22 && x16 && ~x19 && x13 )
						begin
							y3 = 1'b1;	y16 = 1'b1;	
							nx_state = s252;
						end
					else if( x8 && ~x21 && x22 && x16 && ~x19 && ~x13 && x18 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s252;
						end
					else if( x8 && ~x21 && x22 && x16 && ~x19 && ~x13 && ~x18 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x8 && ~x21 && x22 && ~x16 && x17 && x19 && x18 && x10 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else if( x8 && ~x21 && x22 && ~x16 && x17 && x19 && x18 && ~x10 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s252;
						end
					else if( x8 && ~x21 && x22 && ~x16 && x17 && x19 && ~x18 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else if( x8 && ~x21 && x22 && ~x16 && x17 && x19 && ~x18 && ~x13 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( x8 && ~x21 && x22 && ~x16 && x17 && ~x19 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else if( x8 && ~x21 && x22 && ~x16 && x17 && ~x19 && ~x13 && x18 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x8 && ~x21 && x22 && ~x16 && x17 && ~x19 && ~x13 && ~x18 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( x8 && ~x21 && x22 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s252;
						end
					else if( x8 && ~x21 && ~x22 && x19 && x17 && x13 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x8 && ~x21 && ~x22 && x19 && x17 && ~x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x8 && ~x21 && ~x22 && x19 && ~x17 && x18 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else if( x8 && ~x21 && ~x22 && x19 && ~x17 && x18 && ~x13 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( x8 && ~x21 && ~x22 && x19 && ~x17 && ~x18 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s252;
						end
					else if( x8 && ~x21 && ~x22 && ~x19 && x16 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x8 && ~x21 && ~x22 && ~x19 && x16 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s261;
						end
					else if( x8 && ~x21 && ~x22 && ~x19 && ~x16 && x17 && x20 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( x8 && ~x21 && ~x22 && ~x19 && ~x16 && x17 && ~x20 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s810;
						end
					else if( x8 && ~x21 && ~x22 && ~x19 && ~x16 && x17 && ~x20 && ~x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( x8 && ~x21 && ~x22 && ~x19 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x8 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s1332;
						end
					else nx_state = s1331;
				s1332 : if( x21 && x16 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x21 && x16 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s261;
						end
					else if( x21 && ~x16 && x17 && x18 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s810;
						end
					else if( x21 && ~x16 && x17 && x18 && ~x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( x21 && ~x16 && x17 && ~x18 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( x21 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x21 && x22 && x16 && x19 && x18 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x21 && x22 && x16 && x19 && x18 && ~x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s264;
						end
					else if( ~x21 && x22 && x16 && x19 && ~x18 && x13 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && x16 && x19 && ~x18 && ~x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x21 && x22 && x16 && ~x19 && x13 )
						begin
							y3 = 1'b1;	y16 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x21 && x22 && x16 && ~x19 && ~x13 && x18 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x21 && x22 && x16 && ~x19 && ~x13 && ~x18 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x21 && x22 && ~x16 && x17 && x18 && x19 && x10 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else if( ~x21 && x22 && ~x16 && x17 && x18 && x19 && ~x10 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x21 && x22 && ~x16 && x17 && x18 && ~x19 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else if( ~x21 && x22 && ~x16 && x17 && x18 && ~x19 && ~x13 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x21 && x22 && ~x16 && x17 && ~x18 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else if( ~x21 && x22 && ~x16 && x17 && ~x18 && ~x13 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x21 && x22 && ~x16 && x17 && ~x18 && ~x13 && ~x19 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x21 && x22 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x21 && ~x22 && x19 && x17 && x13 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && ~x22 && x19 && x17 && ~x13 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x21 && ~x22 && x19 && ~x17 && x18 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s809;
						end
					else if( ~x21 && ~x22 && x19 && ~x17 && x18 && ~x13 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x21 && ~x22 && x19 && ~x17 && ~x18 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x21 && ~x22 && ~x19 && x16 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x21 && ~x22 && ~x19 && x16 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s261;
						end
					else if( ~x21 && ~x22 && ~x19 && ~x16 && x17 && x20 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( ~x21 && ~x22 && ~x19 && ~x16 && x17 && ~x20 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s810;
						end
					else if( ~x21 && ~x22 && ~x19 && ~x16 && x17 && ~x20 && ~x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s1004;
						end
					else if( ~x21 && ~x22 && ~x19 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s252;
						end
					else nx_state = s1332;
				s1333 : if( x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s1230;
						end
					else nx_state = s1333;
				s1334 : if( x37 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s1230;
						end
					else if( ~x37 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s542;
						end
					else nx_state = s1334;
				s1335 : if( x64 && x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s545;
						end
					else if( x64 && ~x6 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s542;
						end
					else if( ~x64 && x6 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y20 = 1'b1;	
							nx_state = s1230;
						end
					else if( ~x64 && ~x6 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y22 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s801;
						end
					else nx_state = s1335;
				s1336 : if( x64 )
						begin
							y1 = 1'b1;	
							nx_state = s611;
						end
					else if( ~x64 )
						begin
							y7 = 1'b1;	y13 = 1'b1;	y28 = 1'b1;	
							nx_state = s917;
						end
					else nx_state = s1336;
				s1337 : if( x16 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x16 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x16 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x16 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x16 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x16 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y65 = 1'b1;	
							y66 = 1'b1;	
							nx_state = s1041;
						end
					else nx_state = s1337;
				s1338 : if( 1'b1 )
						begin
							y17 = 1'b1;	y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s925;
						end
					else nx_state = s1338;
				s1339 : if( x16 && x22 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1100;
						end
					else if( x16 && x22 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y30 = 1'b1;	
							y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s523;
						end
					else if( x16 && ~x22 )
						begin
							y50 = 1'b1;	
							nx_state = s658;
						end
					else if( ~x16 && x22 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s524;
						end
					else if( ~x16 && ~x22 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s657;
						end
					else nx_state = s1339;
				s1340 : if( 1'b1 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1546;
						end
					else nx_state = s1340;
				s1341 : if( x46 )
						begin
							y9 = 1'b1;	y32 = 1'b1;	y34 = 1'b1;	
							nx_state = s322;
						end
					else if( ~x46 && x14 && x44 )
						begin
							y3 = 1'b1;	y22 = 1'b1;	y24 = 1'b1;	
							nx_state = s1032;
						end
					else if( ~x46 && x14 && ~x44 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( ~x46 && ~x14 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s441;
						end
					else nx_state = s1341;
				s1342 : if( x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s326;
						end
					else if( ~x15 && x14 && x64 && x13 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s498;
						end
					else if( ~x15 && x14 && x64 && ~x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s324;
						end
					else if( ~x15 && x14 && ~x64 && x13 )
						begin
							y19 = 1'b1;	y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s1032;
						end
					else if( ~x15 && x14 && ~x64 && ~x13 )
						begin
							y7 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							nx_state = s1143;
						end
					else if( ~x15 && ~x14 && x64 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s441;
						end
					else if( ~x15 && ~x14 && ~x64 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s1045;
						end
					else nx_state = s1342;
				s1343 : if( x38 && x39 && x41 && x42 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y40 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s1154;
						end
					else if( x38 && x39 && x41 && ~x42 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y40 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s584;
						end
					else if( x38 && x39 && ~x41 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y37 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s939;
						end
					else if( x38 && ~x39 && x40 && x55 && x56 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( x38 && ~x39 && x40 && x55 && ~x56 && x58 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( x38 && ~x39 && x40 && x55 && ~x56 && ~x58 && x59 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s584;
						end
					else if( x38 && ~x39 && x40 && x55 && ~x56 && ~x58 && ~x59 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x38 && ~x39 && x40 && x55 && ~x56 && ~x58 && ~x59 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x38 && ~x39 && x40 && x55 && ~x56 && ~x58 && ~x59 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( x38 && ~x39 && x40 && x55 && ~x56 && ~x58 && ~x59 && ~x27 )
						nx_state = s1;
					else if( x38 && ~x39 && x40 && ~x55 && x54 && x57 && x28 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s584;
						end
					else if( x38 && ~x39 && x40 && ~x55 && x54 && x57 && ~x28 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x38 && ~x39 && x40 && ~x55 && x54 && x57 && ~x28 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x38 && ~x39 && x40 && ~x55 && x54 && x57 && ~x28 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( x38 && ~x39 && x40 && ~x55 && x54 && x57 && ~x28 && ~x27 )
						nx_state = s1;
					else if( x38 && ~x39 && x40 && ~x55 && x54 && ~x57 && x29 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s584;
						end
					else if( x38 && ~x39 && x40 && ~x55 && x54 && ~x57 && ~x29 && x27 && x37 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x38 && ~x39 && x40 && ~x55 && x54 && ~x57 && ~x29 && x27 && ~x37 && x3 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x38 && ~x39 && x40 && ~x55 && x54 && ~x57 && ~x29 && x27 && ~x37 && ~x3 )
						nx_state = s1;
					else if( x38 && ~x39 && x40 && ~x55 && x54 && ~x57 && ~x29 && ~x27 )
						nx_state = s1;
					else if( x38 && ~x39 && x40 && ~x55 && ~x54 && x53 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s584;
						end
					else if( x38 && ~x39 && x40 && ~x55 && ~x54 && ~x53 )
						begin
							y30 = 1'b1;	
							nx_state = s291;
						end
					else if( x38 && ~x39 && ~x40 )
						begin
							y1 = 1'b1;	y13 = 1'b1;	y37 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s1155;
						end
					else if( ~x38 )
						begin
							y2 = 1'b1;	y35 = 1'b1;	y37 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s1156;
						end
					else nx_state = s1343;
				s1344 : if( x3 && x4 && x6 && x8 && x9 && x12 )
						begin
							y47 = 1'b1;	
							nx_state = s287;
						end
					else if( x3 && x4 && x6 && x8 && x9 && ~x12 )
						begin
							y53 = 1'b1;	
							nx_state = s344;
						end
					else if( x3 && x4 && x6 && x8 && ~x9 && x10 && x11 && x16 )
						begin
							y48 = 1'b1;	
							nx_state = s676;
						end
					else if( x3 && x4 && x6 && x8 && ~x9 && x10 && x11 && ~x16 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x3 && x4 && x6 && x8 && ~x9 && x10 && x11 && ~x16 && x14 && ~x15 )
						nx_state = s1;
					else if( x3 && x4 && x6 && x8 && ~x9 && x10 && x11 && ~x16 && ~x14 )
						nx_state = s1;
					else if( x3 && x4 && x6 && x8 && ~x9 && x10 && ~x11 && x15 )
						begin
							y48 = 1'b1;	
							nx_state = s676;
						end
					else if( x3 && x4 && x6 && x8 && ~x9 && x10 && ~x11 && ~x15 && x14 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x3 && x4 && x6 && x8 && ~x9 && x10 && ~x11 && ~x15 && x14 && ~x16 )
						nx_state = s1;
					else if( x3 && x4 && x6 && x8 && ~x9 && x10 && ~x11 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x3 && x4 && x6 && x8 && ~x9 && ~x10 && x11 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y21 = 1'b1;	
							y51 = 1'b1;	y52 = 1'b1;	
							nx_state = s1430;
						end
					else if( x3 && x4 && x6 && x8 && ~x9 && ~x10 && ~x11 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y49 = 1'b1;	y50 = 1'b1;	
							nx_state = s1430;
						end
					else if( x3 && x4 && x6 && ~x8 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s1547;
						end
					else if( x3 && x4 && ~x6 && x12 && x9 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x3 && x4 && ~x6 && x12 && x9 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x3 && x4 && ~x6 && x12 && x9 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x3 && x4 && ~x6 && x12 && x9 && ~x14 )
						nx_state = s1;
					else if( x3 && x4 && ~x6 && x12 && ~x9 && x10 && x8 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x3 && x4 && ~x6 && x12 && ~x9 && x10 && x8 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x3 && x4 && ~x6 && x12 && ~x9 && x10 && x8 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x3 && x4 && ~x6 && x12 && ~x9 && x10 && x8 && ~x14 )
						nx_state = s1;
					else if( x3 && x4 && ~x6 && x12 && ~x9 && x10 && ~x8 && x11 )
						begin
							y5 = 1'b1;	y11 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y29 = 1'b1;	
							nx_state = s1430;
						end
					else if( x3 && x4 && ~x6 && x12 && ~x9 && x10 && ~x8 && ~x11 )
						begin
							y5 = 1'b1;	y11 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y28 = 1'b1;	
							nx_state = s1430;
						end
					else if( x3 && x4 && ~x6 && x12 && ~x9 && ~x10 && x8 && x11 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s1430;
						end
					else if( x3 && x4 && ~x6 && x12 && ~x9 && ~x10 && x8 && ~x11 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x3 && x4 && ~x6 && x12 && ~x9 && ~x10 && x8 && ~x11 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x3 && x4 && ~x6 && x12 && ~x9 && ~x10 && x8 && ~x11 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x3 && x4 && ~x6 && x12 && ~x9 && ~x10 && x8 && ~x11 && ~x14 )
						nx_state = s1;
					else if( x3 && x4 && ~x6 && x12 && ~x9 && ~x10 && ~x8 )
						begin
							y5 = 1'b1;	y11 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s1430;
						end
					else if( x3 && x4 && ~x6 && ~x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s1547;
						end
					else if( x3 && ~x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1548;
						end
					else if( ~x3 )
						begin
							y14 = 1'b1;	
							nx_state = s366;
						end
					else nx_state = s1344;
				s1345 : if( x7 )
						begin
							y31 = 1'b1;	y32 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x7 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x7 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x7 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x7 && ~x17 )
						nx_state = s1;
					else nx_state = s1345;
				s1346 : if( x66 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x66 && ~x8 )
						nx_state = s1;
					else if( ~x66 && x67 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x66 && x67 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x66 && x67 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x17 )
						nx_state = s1;
					else if( ~x66 && ~x67 && x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x66 && ~x67 && x26 && ~x25 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x66 && ~x67 && x26 && ~x25 && ~x24 )
						nx_state = s1;
					else if( ~x66 && ~x67 && ~x26 )
						nx_state = s1;
					else nx_state = s1346;
				s1347 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else nx_state = s1347;
				s1348 : if( x20 && x5 && x6 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y23 = 1'b1;	
							nx_state = s1225;
						end
					else if( x20 && x5 && ~x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y25 = 1'b1;	
							nx_state = s1225;
						end
					else if( x20 && ~x5 )
						begin
							y3 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y30 = 1'b1;	y43 = 1'b1;	
							nx_state = s1345;
						end
					else if( ~x20 && x4 && x21 && x6 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s1270;
						end
					else if( ~x20 && x4 && x21 && x6 && ~x5 && x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x20 && x4 && x21 && x6 && ~x5 && ~x11 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x20 && x4 && x21 && x6 && ~x5 && ~x11 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x20 && x4 && x21 && x6 && ~x5 && ~x11 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x20 && x4 && x21 && x6 && ~x5 && ~x11 && ~x17 )
						nx_state = s1;
					else if( ~x20 && x4 && x21 && ~x6 && x5 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y15 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1347;
						end
					else if( ~x20 && x4 && x21 && ~x6 && ~x5 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x20 && x4 && x21 && ~x6 && ~x5 && ~x10 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x20 && x4 && x21 && ~x6 && ~x5 && ~x10 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x20 && x4 && x21 && ~x6 && ~x5 && ~x10 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x20 && x4 && x21 && ~x6 && ~x5 && ~x10 && ~x17 )
						nx_state = s1;
					else if( ~x20 && x4 && ~x21 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x20 && ~x4 && x21 && x6 && x5 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x20 && ~x4 && x21 && x6 && x5 && ~x13 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x20 && ~x4 && x21 && x6 && x5 && ~x13 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x20 && ~x4 && x21 && x6 && x5 && ~x13 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x20 && ~x4 && x21 && x6 && x5 && ~x13 && ~x17 )
						nx_state = s1;
					else if( ~x20 && ~x4 && x21 && x6 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x20 && ~x4 && x21 && ~x6 && x5 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x20 && ~x4 && x21 && ~x6 && x5 && ~x14 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x20 && ~x4 && x21 && ~x6 && x5 && ~x14 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x20 && ~x4 && x21 && ~x6 && x5 && ~x14 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x20 && ~x4 && x21 && ~x6 && x5 && ~x14 && ~x17 )
						nx_state = s1;
					else if( ~x20 && ~x4 && x21 && ~x6 && ~x5 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x20 && ~x4 && ~x21 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y23 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s1225;
						end
					else nx_state = s1348;
				s1349 : if( x6 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s1330;
						end
					else if( ~x6 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s1171;
						end
					else nx_state = s1349;
				s1350 : if( 1'b1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s806;
						end
					else nx_state = s1350;
				s1351 : if( x18 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x18 )
						begin
							y44 = 1'b1;	y45 = 1'b1;	
							nx_state = s392;
						end
					else nx_state = s1351;
				s1352 : if( x14 )
						begin
							y8 = 1'b1;	
							nx_state = s1549;
						end
					else if( ~x14 )
						begin
							y47 = 1'b1;	y55 = 1'b1;	y61 = 1'b1;	
							y68 = 1'b1;	
							nx_state = s1515;
						end
					else nx_state = s1352;
				s1353 : if( 1'b1 )
						begin
							y13 = 1'b1;	
							nx_state = s1528;
						end
					else nx_state = s1353;
				s1354 : if( 1'b1 )
						begin
							y60 = 1'b1;	y65 = 1'b1;	y78 = 1'b1;	
							y92 = 1'b1;	
							nx_state = s1132;
						end
					else nx_state = s1354;
				s1355 : if( 1'b1 )
						begin
							y1 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s379;
						end
					else nx_state = s1355;
				s1356 : if( x30 )
						begin
							y31 = 1'b1;	
							nx_state = s1053;
						end
					else if( ~x30 && x31 )
						begin
							y47 = 1'b1;	y51 = 1'b1;	y61 = 1'b1;	
							y68 = 1'b1;	
							nx_state = s1316;
						end
					else if( ~x30 && ~x31 )
						begin
							y5 = 1'b1;	
							nx_state = s945;
						end
					else nx_state = s1356;
				s1357 : if( x63 && x67 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s666;
						end
					else if( x63 && ~x67 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x63 && ~x67 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x63 && ~x67 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x63 && ~x67 && ~x14 )
						nx_state = s1;
					else if( ~x63 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s1550;
						end
					else nx_state = s1357;
				s1358 : if( x63 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x63 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x63 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x63 && ~x14 )
						nx_state = s1;
					else if( ~x63 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x63 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x63 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x63 && ~x18 )
						nx_state = s1;
					else nx_state = s1358;
				s1359 : if( x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x14 )
						nx_state = s1;
					else nx_state = s1359;
				s1360 : if( x63 && x14 && x10 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x63 && x14 && ~x10 && x11 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x63 && x14 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x63 && ~x14 )
						nx_state = s1;
					else if( ~x63 && x14 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x63 && x14 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x63 && x14 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x63 && x14 && ~x23 )
						nx_state = s1;
					else if( ~x63 && ~x14 )
						begin
							y47 = 1'b1;	y53 = 1'b1;	y61 = 1'b1;	
							y70 = 1'b1;	
							nx_state = s1473;
						end
					else nx_state = s1360;
				s1361 : if( x12 && x4 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s1362;
						end
					else if( x12 && ~x4 && x5 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s1363;
						end
					else if( x12 && ~x4 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y16 = 1'b1;	
							nx_state = s1359;
						end
					else if( ~x12 && x4 && x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y14 = 1'b1;	
							nx_state = s1359;
						end
					else if( ~x12 && x4 && ~x5 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s1364;
						end
					else if( ~x12 && ~x4 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s1365;
						end
					else nx_state = s1361;
				s1362 : if( 1'b1 )
						begin
							y17 = 1'b1;	
							nx_state = s3;
						end
					else nx_state = s1362;
				s1363 : if( 1'b1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y16 = 1'b1;	
							nx_state = s1359;
						end
					else nx_state = s1363;
				s1364 : if( 1'b1 )
						begin
							y3 = 1'b1;	y13 = 1'b1;	
							nx_state = s1359;
						end
					else nx_state = s1364;
				s1365 : if( x5 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x5 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else nx_state = s1365;
				s1366 : if( 1'b1 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else nx_state = s1366;
				s1367 : if( 1'b1 )
						begin
							y68 = 1'b1;	
							nx_state = s1404;
						end
					else nx_state = s1367;
				s1368 : if( 1'b1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s1551;
						end
					else nx_state = s1368;
				s1369 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y32 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s720;
						end
					else nx_state = s1369;
				s1370 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y32 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else nx_state = s1370;
				s1371 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y59 = 1'b1;	
							y67 = 1'b1;	
							nx_state = s720;
						end
					else nx_state = s1371;
				s1372 : if( x5 && x7 && x6 && x12 && x10 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x5 && x7 && x6 && x12 && ~x10 && x11 && x13 )
						begin
							y13 = 1'b1;	
							nx_state = s240;
						end
					else if( x5 && x7 && x6 && x12 && ~x10 && x11 && ~x13 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x5 && x7 && x6 && x12 && ~x10 && x11 && ~x13 && x19 && ~x14 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( x5 && x7 && x6 && x12 && ~x10 && x11 && ~x13 && ~x19 )
						nx_state = s1;
					else if( x5 && x7 && x6 && x12 && ~x10 && ~x11 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y32 = 1'b1;	
							y53 = 1'b1;	
							nx_state = s954;
						end
					else if( x5 && x7 && x6 && ~x12 && x10 )
						begin
							y25 = 1'b1;	
							nx_state = s955;
						end
					else if( x5 && x7 && x6 && ~x12 && ~x10 && x11 && x14 )
						begin
							y13 = 1'b1;	
							nx_state = s240;
						end
					else if( x5 && x7 && x6 && ~x12 && ~x10 && x11 && ~x14 && x19 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x5 && x7 && x6 && ~x12 && ~x10 && x11 && ~x14 && x19 && ~x13 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( x5 && x7 && x6 && ~x12 && ~x10 && x11 && ~x14 && ~x19 )
						nx_state = s1;
					else if( x5 && x7 && x6 && ~x12 && ~x10 && ~x11 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y54 = 1'b1;	
							nx_state = s956;
						end
					else if( x5 && x7 && ~x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s957;
						end
					else if( x5 && ~x7 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s957;
						end
					else if( x5 && ~x7 && ~x9 && x10 && x11 && x12 && x6 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( x5 && ~x7 && ~x9 && x10 && x11 && x12 && ~x6 )
						begin
							y4 = 1'b1;	y33 = 1'b1;	y34 = 1'b1;	
							y38 = 1'b1;	y42 = 1'b1;	
							nx_state = s720;
						end
					else if( x5 && ~x7 && ~x9 && x10 && x11 && ~x12 && x6 )
						begin
							y29 = 1'b1;	
							nx_state = s771;
						end
					else if( x5 && ~x7 && ~x9 && x10 && x11 && ~x12 && ~x6 )
						begin
							y4 = 1'b1;	y33 = 1'b1;	y34 = 1'b1;	
							y38 = 1'b1;	y41 = 1'b1;	
							nx_state = s720;
						end
					else if( x5 && ~x7 && ~x9 && x10 && ~x11 && x6 && x12 )
						begin
							y30 = 1'b1;	
							nx_state = s291;
						end
					else if( x5 && ~x7 && ~x9 && x10 && ~x11 && x6 && ~x12 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x5 && ~x7 && ~x9 && x10 && ~x11 && ~x6 )
						begin
							y4 = 1'b1;	y33 = 1'b1;	y34 = 1'b1;	
							y38 = 1'b1;	y40 = 1'b1;	
							nx_state = s720;
						end
					else if( x5 && ~x7 && ~x9 && ~x10 && x11 && x12 && x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s959;
						end
					else if( x5 && ~x7 && ~x9 && ~x10 && x11 && x12 && ~x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y59 = 1'b1;	
							y60 = 1'b1;	
							nx_state = s960;
						end
					else if( x5 && ~x7 && ~x9 && ~x10 && x11 && ~x12 && x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y31 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s720;
						end
					else if( x5 && ~x7 && ~x9 && ~x10 && x11 && ~x12 && ~x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y63 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s961;
						end
					else if( x5 && ~x7 && ~x9 && ~x10 && ~x11 && x12 && x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( x5 && ~x7 && ~x9 && ~x10 && ~x11 && x12 && ~x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y61 = 1'b1;	
							y62 = 1'b1;	
							nx_state = s962;
						end
					else if( x5 && ~x7 && ~x9 && ~x10 && ~x11 && ~x12 && x6 )
						begin
							y36 = 1'b1;	
							nx_state = s963;
						end
					else if( x5 && ~x7 && ~x9 && ~x10 && ~x11 && ~x12 && ~x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y65 = 1'b1;	
							y66 = 1'b1;	
							nx_state = s646;
						end
					else if( ~x5 )
						begin
							y17 = 1'b1;	
							nx_state = s3;
						end
					else nx_state = s1372;
				s1373 : if( 1'b1 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else nx_state = s1373;
				s1374 : if( 1'b1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s353;
						end
					else nx_state = s1374;
				s1375 : if( 1'b1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y12 = 1'b1;	
							y37 = 1'b1;	y38 = 1'b1;	
							nx_state = s1552;
						end
					else nx_state = s1375;
				s1376 : if( x8 )
						begin
							y6 = 1'b1;	y47 = 1'b1;	
							nx_state = s1553;
						end
					else if( ~x8 && x32 )
						begin
							y6 = 1'b1;	y47 = 1'b1;	
							nx_state = s1553;
						end
					else if( ~x8 && ~x32 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s340;
						end
					else nx_state = s1376;
				s1377 : if( x15 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x15 )
						nx_state = s1;
					else nx_state = s1377;
				s1378 : if( x10 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s1554;
						end
					else if( ~x10 && x14 && x6 && x5 )
						nx_state = s1;
					else if( ~x10 && x14 && x6 && ~x5 && x7 && x8 )
						begin
							y46 = 1'b1;	
							nx_state = s1428;
						end
					else if( ~x10 && x14 && x6 && ~x5 && x7 && ~x8 && x9 )
						begin
							y3 = 1'b1;	y19 = 1'b1;	y42 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s1555;
						end
					else if( ~x10 && x14 && x6 && ~x5 && x7 && ~x8 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( ~x10 && x14 && x6 && ~x5 && ~x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( ~x10 && x14 && ~x6 )
						begin
							y46 = 1'b1;	
							nx_state = s1428;
						end
					else if( ~x10 && ~x14 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y40 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s1556;
						end
					else nx_state = s1378;
				s1379 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y47 = 1'b1;	
							nx_state = s1557;
						end
					else nx_state = s1379;
				s1380 : if( x5 && x7 && x9 && x6 )
						begin
							y22 = 1'b1;	
							nx_state = s130;
						end
					else if( x5 && x7 && x9 && ~x6 && x8 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x5 && x7 && x9 && ~x6 && ~x8 )
						begin
							y29 = 1'b1;	
							nx_state = s771;
						end
					else if( x5 && x7 && ~x9 && x6 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x5 && x7 && ~x9 && ~x6 && x8 )
						begin
							y30 = 1'b1;	
							nx_state = s291;
						end
					else if( x5 && x7 && ~x9 && ~x6 && ~x8 )
						begin
							y28 = 1'b1;	
							nx_state = s1427;
						end
					else if( x5 && ~x7 && x9 && x6 && x8 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x5 && ~x7 && x9 && x6 && x8 && ~x12 )
						nx_state = s1;
					else if( x5 && ~x7 && x9 && x6 && ~x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1558;
						end
					else if( x5 && ~x7 && x9 && ~x6 && x10 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1556;
						end
					else if( x5 && ~x7 && x9 && ~x6 && ~x10 && x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s1559;
						end
					else if( x5 && ~x7 && x9 && ~x6 && ~x10 && ~x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y15 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1314;
						end
					else if( x5 && ~x7 && ~x9 && x8 && x6 && x13 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x5 && ~x7 && ~x9 && x8 && x6 && ~x13 )
						nx_state = s1;
					else if( x5 && ~x7 && ~x9 && x8 && ~x6 && x10 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s1556;
						end
					else if( x5 && ~x7 && ~x9 && x8 && ~x6 && ~x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y24 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1314;
						end
					else if( x5 && ~x7 && ~x9 && ~x8 && x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s872;
						end
					else if( x5 && ~x7 && ~x9 && ~x8 && ~x6 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x5 && x6 && x8 && x7 && x10 && x3 && x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y17 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1379;
						end
					else if( ~x5 && x6 && x8 && x7 && x10 && x3 && ~x11 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1378;
						end
					else if( ~x5 && x6 && x8 && x7 && x10 && ~x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1556;
						end
					else if( ~x5 && x6 && x8 && x7 && ~x10 )
						begin
							y72 = 1'b1;	
							nx_state = s1377;
						end
					else if( ~x5 && x6 && x8 && ~x7 && x9 && x18 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1378;
						end
					else if( ~x5 && x6 && x8 && ~x7 && x9 && x18 && ~x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1556;
						end
					else if( ~x5 && x6 && x8 && ~x7 && x9 && ~x18 )
						nx_state = s1;
					else if( ~x5 && x6 && x8 && ~x7 && ~x9 && x17 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1378;
						end
					else if( ~x5 && x6 && x8 && ~x7 && ~x9 && x17 && ~x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1556;
						end
					else if( ~x5 && x6 && x8 && ~x7 && ~x9 && ~x17 )
						nx_state = s1;
					else if( ~x5 && x6 && ~x8 && x9 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1378;
						end
					else if( ~x5 && x6 && ~x8 && x9 && ~x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1556;
						end
					else if( ~x5 && x6 && ~x8 && ~x9 && x7 && x16 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1378;
						end
					else if( ~x5 && x6 && ~x8 && ~x9 && x7 && x16 && ~x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1556;
						end
					else if( ~x5 && x6 && ~x8 && ~x9 && x7 && ~x16 )
						nx_state = s1;
					else if( ~x5 && x6 && ~x8 && ~x9 && ~x7 )
						begin
							y71 = 1'b1;	
							nx_state = s394;
						end
					else if( ~x5 && ~x6 && x10 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1556;
						end
					else if( ~x5 && ~x6 && ~x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y15 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s1557;
						end
					else nx_state = s1380;
				s1381 : if( x62 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y23 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s535;
						end
					else if( ~x62 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							nx_state = s1323;
						end
					else nx_state = s1381;
				s1382 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1560;
						end
					else nx_state = s1382;
				s1383 : if( x10 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s1478;
						end
					else if( ~x10 && x11 )
						begin
							y28 = 1'b1;	
							nx_state = s991;
						end
					else if( ~x10 && ~x11 )
						begin
							y29 = 1'b1;	
							nx_state = s1109;
						end
					else nx_state = s1383;
				s1384 : if( 1'b1 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s1561;
						end
					else nx_state = s1384;
				s1385 : if( x65 )
						begin
							y8 = 1'b1;	
							nx_state = s1172;
						end
					else if( ~x65 )
						begin
							y7 = 1'b1;	
							nx_state = s1200;
						end
					else nx_state = s1385;
				s1386 : if( x20 && x26 && x27 && x7 && x8 && x6 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s1220;
						end
					else if( x20 && x26 && x27 && x7 && x8 && ~x6 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y42 = 1'b1;	y44 = 1'b1;	
							nx_state = s1220;
						end
					else if( x20 && x26 && x27 && x7 && ~x8 && x6 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y47 = 1'b1;	
							nx_state = s1220;
						end
					else if( x20 && x26 && x27 && x7 && ~x8 && ~x6 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y42 = 1'b1;	y44 = 1'b1;	
							nx_state = s1220;
						end
					else if( x20 && x26 && x27 && ~x7 && x6 && x8 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1220;
						end
					else if( x20 && x26 && x27 && ~x7 && x6 && ~x8 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y46 = 1'b1;	
							nx_state = s1220;
						end
					else if( x20 && x26 && x27 && ~x7 && ~x6 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y42 = 1'b1;	y44 = 1'b1;	
							nx_state = s1220;
						end
					else if( x20 && x26 && ~x27 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s1562;
						end
					else if( x20 && ~x26 )
						begin
							y58 = 1'b1;	
							nx_state = s1508;
						end
					else if( ~x20 )
						begin
							y26 = 1'b1;	
							nx_state = s262;
						end
					else nx_state = s1386;
				s1387 : if( 1'b1 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s1563;
						end
					else nx_state = s1387;
				s1388 : if( 1'b1 )
						begin
							y6 = 1'b1;	y42 = 1'b1;	y43 = 1'b1;	
							nx_state = s1028;
						end
					else nx_state = s1388;
				s1389 : if( x11 && x19 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1564;
						end
					else if( x11 && ~x19 )
						begin
							y28 = 1'b1;	
							nx_state = s1565;
						end
					else if( ~x11 )
						begin
							y29 = 1'b1;	
							nx_state = s1017;
						end
					else nx_state = s1389;
				s1390 : if( 1'b1 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else nx_state = s1390;
				s1391 : if( 1'b1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y13 = 1'b1;	y34 = 1'b1;	
							nx_state = s1566;
						end
					else nx_state = s1391;
				s1392 : if( x21 )
						begin
							y80 = 1'b1;	
							nx_state = s1567;
						end
					else if( ~x21 )
						begin
							y80 = 1'b1;	
							nx_state = s1568;
						end
					else nx_state = s1392;
				s1393 : if( 1'b1 )
						begin
							y80 = 1'b1;	
							nx_state = s1567;
						end
					else nx_state = s1393;
				s1394 : if( x15 && x17 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x15 && ~x17 && x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x15 && ~x17 && x10 && ~x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x15 && ~x17 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x15 && ~x17 && ~x10 )
						nx_state = s1;
					else if( ~x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else nx_state = s1394;
				s1395 : if( x3 && x5 && x30 && x31 && x9 && x8 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x3 && x5 && x30 && x31 && x9 && x8 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x3 && x5 && x30 && x31 && x9 && x8 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x3 && x5 && x30 && x31 && x9 && x8 && ~x23 )
						nx_state = s1;
					else if( x3 && x5 && x30 && x31 && x9 && ~x8 && x10 && x25 )
						begin
							y29 = 1'b1;	
							nx_state = s771;
						end
					else if( x3 && x5 && x30 && x31 && x9 && ~x8 && x10 && ~x25 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x3 && x5 && x30 && x31 && x9 && ~x8 && x10 && ~x25 && x23 && ~x24 )
						nx_state = s1;
					else if( x3 && x5 && x30 && x31 && x9 && ~x8 && x10 && ~x25 && ~x23 )
						nx_state = s1;
					else if( x3 && x5 && x30 && x31 && x9 && ~x8 && ~x10 && x24 )
						begin
							y29 = 1'b1;	
							nx_state = s771;
						end
					else if( x3 && x5 && x30 && x31 && x9 && ~x8 && ~x10 && ~x24 && x23 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x3 && x5 && x30 && x31 && x9 && ~x8 && ~x10 && ~x24 && x23 && ~x25 )
						nx_state = s1;
					else if( x3 && x5 && x30 && x31 && x9 && ~x8 && ~x10 && ~x24 && ~x23 )
						nx_state = s1;
					else if( x3 && x5 && x30 && x31 && ~x9 && x10 && x8 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s253;
						end
					else if( x3 && x5 && x30 && x31 && ~x9 && x10 && ~x8 )
						begin
							y8 = 1'b1;	
							nx_state = s783;
						end
					else if( x3 && x5 && x30 && x31 && ~x9 && ~x10 && x8 )
						begin
							y10 = 1'b1;	y23 = 1'b1;	
							nx_state = s1;
						end
					else if( x3 && x5 && x30 && x31 && ~x9 && ~x10 && ~x8 )
						begin
							y8 = 1'b1;	
							nx_state = s568;
						end
					else if( x3 && x5 && x30 && ~x31 && x13 )
						begin
							y35 = 1'b1;	
							nx_state = s414;
						end
					else if( x3 && x5 && x30 && ~x31 && ~x13 )
						begin
							y3 = 1'b1;	
							nx_state = s835;
						end
					else if( x3 && x5 && ~x30 && x31 && x15 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x3 && x5 && ~x30 && x31 && x15 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( x3 && x5 && ~x30 && x31 && x15 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x3 && x5 && ~x30 && x31 && x15 && ~x23 )
						nx_state = s1;
					else if( x3 && x5 && ~x30 && x31 && ~x15 && x16 && x13 )
						begin
							y3 = 1'b1;	
							nx_state = s835;
						end
					else if( x3 && x5 && ~x30 && x31 && ~x15 && x16 && ~x13 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( x3 && x5 && ~x30 && x31 && ~x15 && ~x16 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( x3 && x5 && ~x30 && ~x31 && x8 && x9 )
						begin
							y47 = 1'b1;	y55 = 1'b1;	y63 = 1'b1;	
							y70 = 1'b1;	
							nx_state = s1175;
						end
					else if( x3 && x5 && ~x30 && ~x31 && x8 && ~x9 )
						begin
							y47 = 1'b1;	y56 = 1'b1;	y63 = 1'b1;	
							y71 = 1'b1;	
							nx_state = s1175;
						end
					else if( x3 && x5 && ~x30 && ~x31 && ~x8 && x13 )
						begin
							y45 = 1'b1;	y46 = 1'b1;	y47 = 1'b1;	
							y55 = 1'b1;	y59 = 1'b1;	y63 = 1'b1;	
							y70 = 1'b1;	
							nx_state = s1175;
						end
					else if( x3 && x5 && ~x30 && ~x31 && ~x8 && ~x13 )
						begin
							y3 = 1'b1;	
							nx_state = s137;
						end
					else if( x3 && ~x5 && x31 && x30 )
						begin
							y3 = 1'b1;	
							nx_state = s835;
						end
					else if( x3 && ~x5 && x31 && ~x30 )
						begin
							y3 = 1'b1;	
							nx_state = s1569;
						end
					else if( x3 && ~x5 && ~x31 && x30 )
						begin
							y3 = 1'b1;	
							nx_state = s1293;
						end
					else if( x3 && ~x5 && ~x31 && ~x30 )
						begin
							y3 = 1'b1;	
							nx_state = s462;
						end
					else if( ~x3 )
						begin
							y34 = 1'b1;	
							nx_state = s1165;
						end
					else nx_state = s1395;
				s1396 : if( 1'b1 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s1570;
						end
					else nx_state = s1396;
				s1397 : if( x14 && x16 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x14 && x16 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x14 && x16 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x14 && ~x16 )
						nx_state = s1;
					else if( ~x14 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else nx_state = s1397;
				s1398 : if( x9 && x6 && x12 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s1273;
						end
					else if( x9 && x6 && ~x12 && x11 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s1008;
						end
					else if( x9 && x6 && ~x12 && ~x11 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x9 && x6 && ~x12 && ~x11 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x9 && x6 && ~x12 && ~x11 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x9 && x6 && ~x12 && ~x11 && ~x18 )
						nx_state = s1;
					else if( x9 && ~x6 && x8 && x11 && x12 && x10 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x9 && ~x6 && x8 && x11 && x12 && x10 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x9 && ~x6 && x8 && x11 && x12 && x10 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x9 && ~x6 && x8 && x11 && x12 && x10 && ~x18 )
						nx_state = s1;
					else if( x9 && ~x6 && x8 && x11 && x12 && ~x10 && x16 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s749;
						end
					else if( x9 && ~x6 && x8 && x11 && x12 && ~x10 && ~x16 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x9 && ~x6 && x8 && x11 && x12 && ~x10 && ~x16 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x9 && ~x6 && x8 && x11 && x12 && ~x10 && ~x16 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x9 && ~x6 && x8 && x11 && x12 && ~x10 && ~x16 && ~x18 )
						nx_state = s1;
					else if( x9 && ~x6 && x8 && x11 && ~x12 && x10 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s1274;
						end
					else if( x9 && ~x6 && x8 && x11 && ~x12 && ~x10 && x17 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s749;
						end
					else if( x9 && ~x6 && x8 && x11 && ~x12 && ~x10 && ~x17 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x9 && ~x6 && x8 && x11 && ~x12 && ~x10 && ~x17 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x9 && ~x6 && x8 && x11 && ~x12 && ~x10 && ~x17 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x9 && ~x6 && x8 && x11 && ~x12 && ~x10 && ~x17 && ~x18 )
						nx_state = s1;
					else if( x9 && ~x6 && x8 && ~x11 && x12 && x10 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y34 = 1'b1;	
							nx_state = s1275;
						end
					else if( x9 && ~x6 && x8 && ~x11 && x12 && ~x10 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s749;
						end
					else if( x9 && ~x6 && x8 && ~x11 && ~x12 && x10 && x15 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s749;
						end
					else if( x9 && ~x6 && x8 && ~x11 && ~x12 && x10 && ~x15 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x9 && ~x6 && x8 && ~x11 && ~x12 && x10 && ~x15 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( x9 && ~x6 && x8 && ~x11 && ~x12 && x10 && ~x15 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x9 && ~x6 && x8 && ~x11 && ~x12 && x10 && ~x15 && ~x18 )
						nx_state = s1;
					else if( x9 && ~x6 && x8 && ~x11 && ~x12 && ~x10 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x9 && ~x6 && ~x8 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s1273;
						end
					else if( ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y28 = 1'b1;	y33 = 1'b1;	
							nx_state = s750;
						end
					else nx_state = s1398;
				s1399 : if( x63 && x6 && x4 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && x6 && ~x4 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && x6 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x63 && ~x6 && x5 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x63 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x63 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y54 = 1'b1;	
							nx_state = s1400;
						end
					else nx_state = s1399;
				s1400 : if( x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x15 )
						nx_state = s1;
					else nx_state = s1400;
				s1401 : if( x18 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s1249;
						end
					else if( ~x18 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s1401;
						end
					else nx_state = s1401;
				s1402 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s1414;
						end
					else nx_state = s1402;
				s1403 : if( x15 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x15 && x3 && x6 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s1571;
						end
					else if( ~x15 && x3 && x6 && ~x10 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s1439;
						end
					else if( ~x15 && x3 && ~x6 && x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s1439;
						end
					else if( ~x15 && x3 && ~x6 && ~x5 && x10 )
						begin
							y5 = 1'b1;	y23 = 1'b1;	y32 = 1'b1;	
							y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s1571;
						end
					else if( ~x15 && x3 && ~x6 && ~x5 && ~x10 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s1439;
						end
					else if( ~x15 && ~x3 && x4 && x1 && x7 && x6 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x15 && ~x3 && x4 && x1 && x7 && ~x6 && x13 && x8 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x15 && ~x3 && x4 && x1 && x7 && ~x6 && x13 && ~x8 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x15 && ~x3 && x4 && x1 && x7 && ~x6 && x13 && ~x8 && ~x12 && x16 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x15 && ~x3 && x4 && x1 && x7 && ~x6 && x13 && ~x8 && ~x12 && ~x16 )
						nx_state = s1;
					else if( ~x15 && ~x3 && x4 && x1 && x7 && ~x6 && ~x13 && x16 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x15 && ~x3 && x4 && x1 && x7 && ~x6 && ~x13 && x16 && ~x12 )
						nx_state = s1;
					else if( ~x15 && ~x3 && x4 && x1 && x7 && ~x6 && ~x13 && ~x16 )
						nx_state = s1;
					else if( ~x15 && ~x3 && x4 && x1 && ~x7 && x6 )
						begin
							y44 = 1'b1;	
							nx_state = s1138;
						end
					else if( ~x15 && ~x3 && x4 && x1 && ~x7 && ~x6 && x8 )
						begin
							y23 = 1'b1;	y42 = 1'b1;	y43 = 1'b1;	
							nx_state = s1571;
						end
					else if( ~x15 && ~x3 && x4 && x1 && ~x7 && ~x6 && ~x8 )
						begin
							y11 = 1'b1;	y15 = 1'b1;	y41 = 1'b1;	
							nx_state = s1571;
						end
					else if( ~x15 && ~x3 && x4 && ~x1 && x9 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1572;
						end
					else if( ~x15 && ~x3 && x4 && ~x1 && ~x9 && x6 && x8 && x7 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x15 && ~x3 && x4 && ~x1 && ~x9 && x6 && x8 && ~x7 )
						begin
							y39 = 1'b1;	
							nx_state = s277;
						end
					else if( ~x15 && ~x3 && x4 && ~x1 && ~x9 && x6 && ~x8 && x7 )
						begin
							y40 = 1'b1;	
							nx_state = s751;
						end
					else if( ~x15 && ~x3 && x4 && ~x1 && ~x9 && x6 && ~x8 && ~x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y33 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s1571;
						end
					else if( ~x15 && ~x3 && x4 && ~x1 && ~x9 && ~x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y33 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s1571;
						end
					else if( ~x15 && ~x3 && ~x4 && x5 && x7 && x6 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1573;
						end
					else if( ~x15 && ~x3 && ~x4 && x5 && x7 && ~x6 && x11 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x15 && ~x3 && ~x4 && x5 && x7 && ~x6 && ~x11 && x16 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x15 && ~x3 && ~x4 && x5 && x7 && ~x6 && ~x11 && x16 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x15 && ~x3 && ~x4 && x5 && x7 && ~x6 && ~x11 && x16 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x15 && ~x3 && ~x4 && x5 && x7 && ~x6 && ~x11 && ~x16 )
						nx_state = s1;
					else if( ~x15 && ~x3 && ~x4 && x5 && ~x7 && x8 && x6 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1574;
						end
					else if( ~x15 && ~x3 && ~x4 && x5 && ~x7 && x8 && ~x6 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1575;
						end
					else if( ~x15 && ~x3 && ~x4 && x5 && ~x7 && ~x8 && x6 && x11 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x15 && ~x3 && ~x4 && x5 && ~x7 && ~x8 && x6 && ~x11 && x16 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x15 && ~x3 && ~x4 && x5 && ~x7 && ~x8 && x6 && ~x11 && x16 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x15 && ~x3 && ~x4 && x5 && ~x7 && ~x8 && x6 && ~x11 && x16 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x15 && ~x3 && ~x4 && x5 && ~x7 && ~x8 && x6 && ~x11 && ~x16 )
						nx_state = s1;
					else if( ~x15 && ~x3 && ~x4 && x5 && ~x7 && ~x8 && ~x6 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x15 && ~x3 && ~x4 && ~x5 && x9 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1572;
						end
					else if( ~x15 && ~x3 && ~x4 && ~x5 && ~x9 && x6 )
						begin
							y5 = 1'b1;	y34 = 1'b1;	y35 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1405;
						end
					else if( ~x15 && ~x3 && ~x4 && ~x5 && ~x9 && ~x6 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s1571;
						end
					else nx_state = s1403;
				s1404 : if( x63 && x66 )
						begin
							y69 = 1'b1;	
							nx_state = s1123;
						end
					else if( x63 && ~x66 && x11 && x6 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( x63 && ~x66 && x11 && x6 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( x63 && ~x66 && x11 && ~x6 && x7 && x10 )
						begin
							y48 = 1'b1;	
							nx_state = s1009;
						end
					else if( x63 && ~x66 && x11 && ~x6 && x7 && ~x10 && x12 && x18 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y47 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s720;
						end
					else if( x63 && ~x66 && x11 && ~x6 && x7 && ~x10 && x12 && ~x18 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x63 && ~x66 && x11 && ~x6 && x7 && ~x10 && x12 && ~x18 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x63 && ~x66 && x11 && ~x6 && x7 && ~x10 && x12 && ~x18 && x19 && ~x14 && ~x13 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( x63 && ~x66 && x11 && ~x6 && x7 && ~x10 && x12 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x63 && ~x66 && x11 && ~x6 && x7 && ~x10 && ~x12 && x17 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y47 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s720;
						end
					else if( x63 && ~x66 && x11 && ~x6 && x7 && ~x10 && ~x12 && ~x17 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x63 && ~x66 && x11 && ~x6 && x7 && ~x10 && ~x12 && ~x17 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x63 && ~x66 && x11 && ~x6 && x7 && ~x10 && ~x12 && ~x17 && x19 && ~x14 && ~x13 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( x63 && ~x66 && x11 && ~x6 && x7 && ~x10 && ~x12 && ~x17 && ~x19 )
						nx_state = s1;
					else if( x63 && ~x66 && x11 && ~x6 && ~x7 && x12 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	y38 = 1'b1;	y40 = 1'b1;	
							nx_state = s720;
						end
					else if( x63 && ~x66 && x11 && ~x6 && ~x7 && ~x12 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	y38 = 1'b1;	y41 = 1'b1;	
							nx_state = s720;
						end
					else if( x63 && ~x66 && ~x11 && x6 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( x63 && ~x66 && ~x11 && ~x6 && x7 && x12 && x10 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y45 = 1'b1;	
							y49 = 1'b1;	
							nx_state = s1576;
						end
					else if( x63 && ~x66 && ~x11 && ~x6 && x7 && x12 && ~x10 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y47 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s720;
						end
					else if( x63 && ~x66 && ~x11 && ~x6 && x7 && ~x12 && x10 && x16 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y47 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s720;
						end
					else if( x63 && ~x66 && ~x11 && ~x6 && x7 && ~x12 && x10 && ~x16 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x63 && ~x66 && ~x11 && ~x6 && x7 && ~x12 && x10 && ~x16 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x63 && ~x66 && ~x11 && ~x6 && x7 && ~x12 && x10 && ~x16 && x19 && ~x14 && ~x13 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( x63 && ~x66 && ~x11 && ~x6 && x7 && ~x12 && x10 && ~x16 && ~x19 )
						nx_state = s1;
					else if( x63 && ~x66 && ~x11 && ~x6 && x7 && ~x12 && ~x10 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x63 && ~x66 && ~x11 && ~x6 && ~x7 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	y38 = 1'b1;	y42 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x63 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x63 && ~x15 )
						nx_state = s1;
					else nx_state = s1404;
				s1405 : if( x63 && x16 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x63 && x16 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x63 && x16 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x63 && ~x16 )
						nx_state = s1;
					else if( ~x63 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x63 && ~x15 )
						nx_state = s1;
					else nx_state = s1405;
				s1406 : if( x65 && x10 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1577;
						end
					else if( x65 && ~x10 && x18 && x8 && x7 )
						begin
							y5 = 1'b1;	y19 = 1'b1;	y25 = 1'b1;	
							y27 = 1'b1;	y30 = 1'b1;	
							nx_state = s1578;
						end
					else if( x65 && ~x10 && x18 && x8 && ~x7 && x9 && x14 )
						begin
							y61 = 1'b1;	
							nx_state = s1098;
						end
					else if( x65 && ~x10 && x18 && x8 && ~x7 && x9 && ~x14 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x65 && ~x10 && x18 && x8 && ~x7 && x9 && ~x14 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x65 && ~x10 && x18 && x8 && ~x7 && x9 && ~x14 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x10 && x18 && x8 && ~x7 && x9 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x65 && ~x10 && x18 && x8 && ~x7 && ~x9 && x12 )
						begin
							y61 = 1'b1;	
							nx_state = s1098;
						end
					else if( x65 && ~x10 && x18 && x8 && ~x7 && ~x9 && ~x12 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x65 && ~x10 && x18 && x8 && ~x7 && ~x9 && ~x12 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x65 && ~x10 && x18 && x8 && ~x7 && ~x9 && ~x12 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x10 && x18 && x8 && ~x7 && ~x9 && ~x12 && ~x15 )
						nx_state = s1;
					else if( x65 && ~x10 && x18 && ~x8 && x9 && x7 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y26 = 1'b1;	
							nx_state = s1579;
						end
					else if( x65 && ~x10 && x18 && ~x8 && x9 && ~x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s1580;
						end
					else if( x65 && ~x10 && x18 && ~x8 && ~x9 && x7 && x13 )
						begin
							y61 = 1'b1;	
							nx_state = s1098;
						end
					else if( x65 && ~x10 && x18 && ~x8 && ~x9 && x7 && ~x13 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x65 && ~x10 && x18 && ~x8 && ~x9 && x7 && ~x13 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x65 && ~x10 && x18 && ~x8 && ~x9 && x7 && ~x13 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x10 && x18 && ~x8 && ~x9 && x7 && ~x13 && ~x15 )
						nx_state = s1;
					else if( x65 && ~x10 && x18 && ~x8 && ~x9 && ~x7 )
						begin
							y69 = 1'b1;	
							nx_state = s1123;
						end
					else if( x65 && ~x10 && ~x18 )
						begin
							y5 = 1'b1;	y19 = 1'b1;	y23 = 1'b1;	
							y25 = 1'b1;	y27 = 1'b1;	
							nx_state = s1581;
						end
					else if( ~x65 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x17 )
						nx_state = s1;
					else nx_state = s1406;
				s1407 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s1582;
						end
					else nx_state = s1407;
				s1408 : if( x10 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1583;
						end
					else if( ~x10 && x18 && x8 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s1584;
						end
					else if( ~x10 && x18 && x8 && ~x9 )
						begin
							y3 = 1'b1;	y26 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1400;
						end
					else if( ~x10 && x18 && ~x8 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1400;
						end
					else if( ~x10 && ~x18 )
						begin
							y5 = 1'b1;	y19 = 1'b1;	y23 = 1'b1;	
							y25 = 1'b1;	y27 = 1'b1;	
							nx_state = s1585;
						end
					else nx_state = s1408;
				s1409 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y50 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s1586;
						end
					else nx_state = s1409;
				s1410 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y40 = 1'b1;	
							y59 = 1'b1;	
							nx_state = s1587;
						end
					else nx_state = s1410;
				s1411 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y52 = 1'b1;	
							nx_state = s1400;
						end
					else nx_state = s1411;
				s1412 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y41 = 1'b1;	
							nx_state = s1400;
						end
					else nx_state = s1412;
				s1413 : if( x10 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1588;
						end
					else if( ~x10 && x18 && x8 && x9 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y55 = 1'b1;	y65 = 1'b1;	
							nx_state = s1589;
						end
					else if( ~x10 && x18 && x8 && x9 && ~x7 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1400;
						end
					else if( ~x10 && x18 && x8 && ~x9 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y47 = 1'b1;	y49 = 1'b1;	
							nx_state = s1590;
						end
					else if( ~x10 && x18 && x8 && ~x9 && ~x7 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							y20 = 1'b1;	y22 = 1'b1;	
							nx_state = s1400;
						end
					else if( ~x10 && x18 && ~x8 && x7 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y66 = 1'b1;	
							y67 = 1'b1;	
							nx_state = s1591;
						end
					else if( ~x10 && x18 && ~x8 && x7 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y56 = 1'b1;	
							y57 = 1'b1;	
							nx_state = s1592;
						end
					else if( ~x10 && x18 && ~x8 && ~x7 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	y22 = 1'b1;	
							nx_state = s1400;
						end
					else if( ~x10 && ~x18 )
						begin
							y5 = 1'b1;	y19 = 1'b1;	y23 = 1'b1;	
							y25 = 1'b1;	y27 = 1'b1;	
							nx_state = s1593;
						end
					else nx_state = s1413;
				s1414 : if( x65 && x4 )
						begin
							y24 = 1'b1;	
							nx_state = s1317;
						end
					else if( x65 && ~x4 && x5 && x6 && x9 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s11;
						end
					else if( x65 && ~x4 && x5 && x6 && x9 && ~x7 && x8 && x17 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x65 && ~x4 && x5 && x6 && x9 && ~x7 && x8 && ~x17 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x65 && ~x4 && x5 && x6 && x9 && ~x7 && x8 && ~x17 && x15 && ~x16 )
						nx_state = s1;
					else if( x65 && ~x4 && x5 && x6 && x9 && ~x7 && x8 && ~x17 && ~x15 )
						nx_state = s1;
					else if( x65 && ~x4 && x5 && x6 && x9 && ~x7 && ~x8 )
						begin
							y5 = 1'b1;	y31 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1400;
						end
					else if( x65 && ~x4 && x5 && x6 && ~x9 && x7 )
						begin
							y68 = 1'b1;	
							nx_state = s1404;
						end
					else if( x65 && ~x4 && x5 && x6 && ~x9 && ~x7 && x8 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( x65 && ~x4 && x5 && x6 && ~x9 && ~x7 && x8 && ~x18 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x65 && ~x4 && x5 && x6 && ~x9 && ~x7 && x8 && ~x18 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x65 && ~x4 && x5 && x6 && ~x9 && ~x7 && x8 && ~x18 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x4 && x5 && x6 && ~x9 && ~x7 && x8 && ~x18 && ~x15 )
						nx_state = s1;
					else if( x65 && ~x4 && x5 && x6 && ~x9 && ~x7 && ~x8 )
						begin
							y5 = 1'b1;	y34 = 1'b1;	y35 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1405;
						end
					else if( x65 && ~x4 && x5 && ~x6 && x7 && x9 && x8 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( x65 && ~x4 && x5 && ~x6 && x7 && x9 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s98;
						end
					else if( x65 && ~x4 && x5 && ~x6 && x7 && ~x9 && x8 )
						begin
							y18 = 1'b1;	
							nx_state = s530;
						end
					else if( x65 && ~x4 && x5 && ~x6 && x7 && ~x9 && ~x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x65 && ~x4 && x5 && ~x6 && ~x7 && x8 && x3 && x11 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s1407;
						end
					else if( x65 && ~x4 && x5 && ~x6 && ~x7 && x8 && x3 && x11 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y28 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s1400;
						end
					else if( x65 && ~x4 && x5 && ~x6 && ~x7 && x8 && x3 && ~x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1408;
						end
					else if( x65 && ~x4 && x5 && ~x6 && ~x7 && x8 && ~x3 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y23 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1585;
						end
					else if( x65 && ~x4 && x5 && ~x6 && ~x7 && x8 && ~x3 && ~x10 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y35 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s1594;
						end
					else if( x65 && ~x4 && x5 && ~x6 && ~x7 && x8 && ~x3 && ~x10 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y37 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s1595;
						end
					else if( x65 && ~x4 && x5 && ~x6 && ~x7 && ~x8 && x9 && x3 && x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1400;
						end
					else if( x65 && ~x4 && x5 && ~x6 && ~x7 && ~x8 && x9 && x3 && ~x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1408;
						end
					else if( x65 && ~x4 && x5 && ~x6 && ~x7 && ~x8 && x9 && ~x3 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y23 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1585;
						end
					else if( x65 && ~x4 && x5 && ~x6 && ~x7 && ~x8 && x9 && ~x3 && ~x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y22 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s1310;
						end
					else if( x65 && ~x4 && x5 && ~x6 && ~x7 && ~x8 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y22 = 1'b1;	
							nx_state = s1400;
						end
					else if( x65 && ~x4 && ~x5 && x6 && x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1406;
						end
					else if( x65 && ~x4 && ~x5 && x6 && ~x3 && x8 && x7 )
						begin
							y5 = 1'b1;	y19 = 1'b1;	y30 = 1'b1;	
							y39 = 1'b1;	y60 = 1'b1;	
							nx_state = s1596;
						end
					else if( x65 && ~x4 && ~x5 && x6 && ~x3 && x8 && ~x7 && x9 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s1580;
						end
					else if( x65 && ~x4 && ~x5 && x6 && ~x3 && x8 && ~x7 && x9 && ~x14 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x65 && ~x4 && ~x5 && x6 && ~x3 && x8 && ~x7 && x9 && ~x14 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x65 && ~x4 && ~x5 && x6 && ~x3 && x8 && ~x7 && x9 && ~x14 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x4 && ~x5 && x6 && ~x3 && x8 && ~x7 && x9 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x65 && ~x4 && ~x5 && x6 && ~x3 && x8 && ~x7 && ~x9 && x12 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s1580;
						end
					else if( x65 && ~x4 && ~x5 && x6 && ~x3 && x8 && ~x7 && ~x9 && ~x12 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x65 && ~x4 && ~x5 && x6 && ~x3 && x8 && ~x7 && ~x9 && ~x12 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x65 && ~x4 && ~x5 && x6 && ~x3 && x8 && ~x7 && ~x9 && ~x12 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x4 && ~x5 && x6 && ~x3 && x8 && ~x7 && ~x9 && ~x12 && ~x15 )
						nx_state = s1;
					else if( x65 && ~x4 && ~x5 && x6 && ~x3 && ~x8 && x9 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y22 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s1597;
						end
					else if( x65 && ~x4 && ~x5 && x6 && ~x3 && ~x8 && x9 && ~x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y23 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1598;
						end
					else if( x65 && ~x4 && ~x5 && x6 && ~x3 && ~x8 && ~x9 && x7 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s1580;
						end
					else if( x65 && ~x4 && ~x5 && x6 && ~x3 && ~x8 && ~x9 && x7 && ~x13 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x65 && ~x4 && ~x5 && x6 && ~x3 && ~x8 && ~x9 && x7 && ~x13 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x65 && ~x4 && ~x5 && x6 && ~x3 && ~x8 && ~x9 && x7 && ~x13 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x4 && ~x5 && x6 && ~x3 && ~x8 && ~x9 && x7 && ~x13 && ~x15 )
						nx_state = s1;
					else if( x65 && ~x4 && ~x5 && x6 && ~x3 && ~x8 && ~x9 && ~x7 )
						begin
							y69 = 1'b1;	
							nx_state = s1123;
						end
					else if( x65 && ~x4 && ~x5 && ~x6 && x3 && x11 && x8 && x9 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y47 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s1409;
						end
					else if( x65 && ~x4 && ~x5 && ~x6 && x3 && x11 && x8 && x9 && ~x7 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1400;
						end
					else if( x65 && ~x4 && ~x5 && ~x6 && x3 && x11 && x8 && ~x9 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y47 = 1'b1;	
							y58 = 1'b1;	
							nx_state = s1410;
						end
					else if( x65 && ~x4 && ~x5 && ~x6 && x3 && x11 && x8 && ~x9 && ~x7 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	y14 = 1'b1;	
							y20 = 1'b1;	y22 = 1'b1;	
							nx_state = s1400;
						end
					else if( x65 && ~x4 && ~x5 && ~x6 && x3 && x11 && ~x8 && x7 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y50 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s1411;
						end
					else if( x65 && ~x4 && ~x5 && ~x6 && x3 && x11 && ~x8 && x7 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y40 = 1'b1;	
							y59 = 1'b1;	
							nx_state = s1412;
						end
					else if( x65 && ~x4 && ~x5 && ~x6 && x3 && x11 && ~x8 && ~x7 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	y22 = 1'b1;	
							nx_state = s1400;
						end
					else if( x65 && ~x4 && ~x5 && ~x6 && x3 && ~x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1413;
						end
					else if( x65 && ~x4 && ~x5 && ~x6 && ~x3 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y23 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1593;
						end
					else if( x65 && ~x4 && ~x5 && ~x6 && ~x3 && ~x10 && x8 && x9 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y47 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s1599;
						end
					else if( x65 && ~x4 && ~x5 && ~x6 && ~x3 && ~x10 && x8 && x9 && ~x7 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	y23 = 1'b1;	
							nx_state = s1400;
						end
					else if( x65 && ~x4 && ~x5 && ~x6 && ~x3 && ~x10 && x8 && ~x9 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y46 = 1'b1;	
							y47 = 1'b1;	
							nx_state = s1600;
						end
					else if( x65 && ~x4 && ~x5 && ~x6 && ~x3 && ~x10 && x8 && ~x9 && ~x7 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y20 = 1'b1;	
							y22 = 1'b1;	y23 = 1'b1;	
							nx_state = s1400;
						end
					else if( x65 && ~x4 && ~x5 && ~x6 && ~x3 && ~x10 && ~x8 && x7 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y44 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1399;
						end
					else if( x65 && ~x4 && ~x5 && ~x6 && ~x3 && ~x10 && ~x8 && x7 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y42 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s1042;
						end
					else if( x65 && ~x4 && ~x5 && ~x6 && ~x3 && ~x10 && ~x8 && ~x7 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y19 = 1'b1;	
							y22 = 1'b1;	y23 = 1'b1;	
							nx_state = s1400;
						end
					else if( ~x65 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s1249;
						end
					else nx_state = s1414;
				s1415 : if( x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s938;
						end
					else if( ~x3 && x19 && x20 && x5 && x6 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y23 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x3 && x19 && x20 && x5 && ~x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y25 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x3 && x19 && x20 && ~x5 )
						begin
							y3 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y30 = 1'b1;	y43 = 1'b1;	
							nx_state = s1345;
						end
					else if( ~x3 && x19 && ~x20 && x4 && x21 && x6 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s1270;
						end
					else if( ~x3 && x19 && ~x20 && x4 && x21 && x6 && ~x5 && x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x3 && x19 && ~x20 && x4 && x21 && x6 && ~x5 && ~x11 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x3 && x19 && ~x20 && x4 && x21 && x6 && ~x5 && ~x11 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x3 && x19 && ~x20 && x4 && x21 && x6 && ~x5 && ~x11 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x3 && x19 && ~x20 && x4 && x21 && x6 && ~x5 && ~x11 && ~x17 )
						nx_state = s1;
					else if( ~x3 && x19 && ~x20 && x4 && x21 && ~x6 && x5 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y15 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1347;
						end
					else if( ~x3 && x19 && ~x20 && x4 && x21 && ~x6 && ~x5 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x3 && x19 && ~x20 && x4 && x21 && ~x6 && ~x5 && ~x10 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x3 && x19 && ~x20 && x4 && x21 && ~x6 && ~x5 && ~x10 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x3 && x19 && ~x20 && x4 && x21 && ~x6 && ~x5 && ~x10 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x3 && x19 && ~x20 && x4 && x21 && ~x6 && ~x5 && ~x10 && ~x17 )
						nx_state = s1;
					else if( ~x3 && x19 && ~x20 && x4 && ~x21 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x3 && x19 && ~x20 && ~x4 && x21 && x6 && x5 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x3 && x19 && ~x20 && ~x4 && x21 && x6 && x5 && ~x13 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x3 && x19 && ~x20 && ~x4 && x21 && x6 && x5 && ~x13 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x3 && x19 && ~x20 && ~x4 && x21 && x6 && x5 && ~x13 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x3 && x19 && ~x20 && ~x4 && x21 && x6 && x5 && ~x13 && ~x17 )
						nx_state = s1;
					else if( ~x3 && x19 && ~x20 && ~x4 && x21 && x6 && ~x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x3 && x19 && ~x20 && ~x4 && x21 && ~x6 && x5 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x3 && x19 && ~x20 && ~x4 && x21 && ~x6 && x5 && ~x14 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x3 && x19 && ~x20 && ~x4 && x21 && ~x6 && x5 && ~x14 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x3 && x19 && ~x20 && ~x4 && x21 && ~x6 && x5 && ~x14 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x3 && x19 && ~x20 && ~x4 && x21 && ~x6 && x5 && ~x14 && ~x17 )
						nx_state = s1;
					else if( ~x3 && x19 && ~x20 && ~x4 && x21 && ~x6 && ~x5 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x3 && x19 && ~x20 && ~x4 && ~x21 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y23 = 1'b1;	y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x3 && ~x19 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s1348;
						end
					else nx_state = s1415;
				s1416 : if( x7 )
						begin
							y31 = 1'b1;	y32 = 1'b1;	
							nx_state = s1225;
						end
					else if( ~x7 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x7 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x7 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x7 && ~x17 )
						nx_state = s1;
					else nx_state = s1416;
				s1417 : if( x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x26 && ~x25 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x26 && ~x25 && ~x24 )
						nx_state = s1;
					else if( ~x26 )
						nx_state = s1;
					else nx_state = s1417;
				s1418 : if( x14 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s1417;
						end
					else if( x14 && ~x5 && x6 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x14 && ~x5 && ~x6 )
						begin
							y25 = 1'b1;	y26 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s1417;
						end
					else if( ~x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s743;
						end
					else nx_state = s1418;
				s1419 : if( x4 )
						begin
							y10 = 1'b1;	
							nx_state = s841;
						end
					else if( ~x4 && x6 && x5 && x21 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y13 = 1'b1;	
							y31 = 1'b1;	y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s1417;
						end
					else if( ~x4 && x6 && x5 && x21 && ~x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y13 = 1'b1;	
							y34 = 1'b1;	y36 = 1'b1;	
							nx_state = s1417;
						end
					else if( ~x4 && x6 && x5 && ~x21 && x22 && x10 && x24 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( ~x4 && x6 && x5 && ~x21 && x22 && x10 && ~x24 && x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x4 && x6 && x5 && ~x21 && x22 && x10 && ~x24 && x26 && ~x25 )
						nx_state = s1;
					else if( ~x4 && x6 && x5 && ~x21 && x22 && x10 && ~x24 && ~x26 )
						nx_state = s1;
					else if( ~x4 && x6 && x5 && ~x21 && x22 && ~x10 && x25 )
						begin
							y9 = 1'b1;	
							nx_state = s400;
						end
					else if( ~x4 && x6 && x5 && ~x21 && x22 && ~x10 && ~x25 && x26 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x4 && x6 && x5 && ~x21 && x22 && ~x10 && ~x25 && x26 && ~x24 )
						nx_state = s1;
					else if( ~x4 && x6 && x5 && ~x21 && x22 && ~x10 && ~x25 && ~x26 )
						nx_state = s1;
					else if( ~x4 && x6 && x5 && ~x21 && ~x22 && x23 && x10 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( ~x4 && x6 && x5 && ~x21 && ~x22 && x23 && ~x10 )
						begin
							y22 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x4 && x6 && x5 && ~x21 && ~x22 && ~x23 && x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x4 && x6 && x5 && ~x21 && ~x22 && ~x23 && x26 && ~x25 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x4 && x6 && x5 && ~x21 && ~x22 && ~x23 && x26 && ~x25 && ~x24 )
						nx_state = s1;
					else if( ~x4 && x6 && x5 && ~x21 && ~x22 && ~x23 && ~x26 )
						nx_state = s1;
					else if( ~x4 && x6 && ~x5 && x9 && x8 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1269;
						end
					else if( ~x4 && x6 && ~x5 && x9 && x8 && ~x15 && x17 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x4 && x6 && ~x5 && x9 && x8 && ~x15 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x4 && x6 && ~x5 && x9 && ~x8 && x10 && x11 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1269;
						end
					else if( ~x4 && x6 && ~x5 && x9 && ~x8 && x10 && x11 && ~x15 && x17 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x4 && x6 && ~x5 && x9 && ~x8 && x10 && x11 && ~x15 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x4 && x6 && ~x5 && x9 && ~x8 && x10 && ~x11 && x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x4 && x6 && ~x5 && x9 && ~x8 && x10 && ~x11 && x26 && ~x25 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x4 && x6 && ~x5 && x9 && ~x8 && x10 && ~x11 && x26 && ~x25 && ~x24 )
						nx_state = s1;
					else if( ~x4 && x6 && ~x5 && x9 && ~x8 && x10 && ~x11 && ~x26 )
						nx_state = s1;
					else if( ~x4 && x6 && ~x5 && x9 && ~x8 && ~x10 && x12 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1269;
						end
					else if( ~x4 && x6 && ~x5 && x9 && ~x8 && ~x10 && x12 && ~x15 && x17 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x4 && x6 && ~x5 && x9 && ~x8 && ~x10 && x12 && ~x15 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x4 && x6 && ~x5 && x9 && ~x8 && ~x10 && ~x12 && x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x4 && x6 && ~x5 && x9 && ~x8 && ~x10 && ~x12 && x26 && ~x25 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x4 && x6 && ~x5 && x9 && ~x8 && ~x10 && ~x12 && x26 && ~x25 && ~x24 )
						nx_state = s1;
					else if( ~x4 && x6 && ~x5 && x9 && ~x8 && ~x10 && ~x12 && ~x26 )
						nx_state = s1;
					else if( ~x4 && x6 && ~x5 && ~x9 && x10 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s1601;
						end
					else if( ~x4 && x6 && ~x5 && ~x9 && x10 && ~x8 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1269;
						end
					else if( ~x4 && x6 && ~x5 && ~x9 && x10 && ~x8 && ~x15 && x17 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x4 && x6 && ~x5 && ~x9 && x10 && ~x8 && ~x15 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x4 && x6 && ~x5 && ~x9 && ~x10 && x8 && x13 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1269;
						end
					else if( ~x4 && x6 && ~x5 && ~x9 && ~x10 && x8 && x13 && ~x15 && x17 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x4 && x6 && ~x5 && ~x9 && ~x10 && x8 && x13 && ~x15 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x4 && x6 && ~x5 && ~x9 && ~x10 && x8 && ~x13 && x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x4 && x6 && ~x5 && ~x9 && ~x10 && x8 && ~x13 && x26 && ~x25 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x4 && x6 && ~x5 && ~x9 && ~x10 && x8 && ~x13 && x26 && ~x25 && ~x24 )
						nx_state = s1;
					else if( ~x4 && x6 && ~x5 && ~x9 && ~x10 && x8 && ~x13 && ~x26 )
						nx_state = s1;
					else if( ~x4 && x6 && ~x5 && ~x9 && ~x10 && ~x8 )
						begin
							y30 = 1'b1;	
							nx_state = s291;
						end
					else if( ~x4 && ~x6 && x5 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y26 = 1'b1;	
							y37 = 1'b1;	y38 = 1'b1;	
							nx_state = s1417;
						end
					else if( ~x4 && ~x6 && x5 && ~x7 && x8 )
						begin
							y5 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s1417;
						end
					else if( ~x4 && ~x6 && x5 && ~x7 && ~x8 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1269;
						end
					else if( ~x4 && ~x6 && x5 && ~x7 && ~x8 && ~x15 && x9 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1602;
						end
					else if( ~x4 && ~x6 && x5 && ~x7 && ~x8 && ~x15 && x9 && ~x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s1580;
						end
					else if( ~x4 && ~x6 && x5 && ~x7 && ~x8 && ~x15 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s1417;
						end
					else if( ~x4 && ~x6 && ~x5 && x8 )
						begin
							y5 = 1'b1;	y23 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1417;
						end
					else if( ~x4 && ~x6 && ~x5 && ~x8 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1269;
						end
					else if( ~x4 && ~x6 && ~x5 && ~x8 && ~x15 )
						begin
							y5 = 1'b1;	y23 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	y39 = 1'b1;	
							nx_state = s1417;
						end
					else nx_state = s1419;
				s1420 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s1603;
						end
					else nx_state = s1420;
				s1421 : if( 1'b1 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s81;
						end
					else nx_state = s1421;
				s1422 : if( x15 )
						begin
							y5 = 1'b1;	y42 = 1'b1;	y43 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s1604;
						end
					else if( ~x15 )
						begin
							y5 = 1'b1;	y42 = 1'b1;	y43 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s1057;
						end
					else nx_state = s1422;
				s1423 : if( x62 )
						begin
							y53 = 1'b1;	
							nx_state = s285;
						end
					else if( ~x62 )
						begin
							y25 = 1'b1;	
							nx_state = s1605;
						end
					else nx_state = s1423;
				s1424 : if( x62 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x62 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x62 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x62 && ~x10 )
						nx_state = s1;
					else if( ~x62 )
						begin
							y2 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1606;
						end
					else nx_state = s1424;
				s1425 : if( x33 && x32 )
						begin
							y53 = 1'b1;	
							nx_state = s344;
						end
					else if( x33 && ~x32 && x30 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	
							nx_state = s1061;
						end
					else if( x33 && ~x32 && ~x30 && x10 && x11 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x33 && ~x32 && ~x30 && x10 && ~x11 && x12 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( x33 && ~x32 && ~x30 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x33 && ~x32 && ~x30 && ~x10 )
						nx_state = s1;
					else if( ~x33 )
						begin
							y53 = 1'b1;	
							nx_state = s344;
						end
					else nx_state = s1425;
				s1426 : if( 1'b1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	y45 = 1'b1;	
							nx_state = s1607;
						end
					else nx_state = s1426;
				s1427 : if( x63 && x20 && x9 )
						begin
							y15 = 1'b1;	
							nx_state = s243;
						end
					else if( x63 && x20 && ~x9 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							nx_state = s1323;
						end
					else if( x63 && ~x20 && x9 )
						begin
							y15 = 1'b1;	
							nx_state = s1115;
						end
					else if( x63 && ~x20 && ~x9 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( ~x63 && x21 && x22 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x63 && x21 && ~x22 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x63 && x21 && ~x22 && ~x23 )
						nx_state = s1;
					else if( ~x63 && ~x21 && x23 )
						begin
							y70 = 1'b1;	
							nx_state = s533;
						end
					else if( ~x63 && ~x21 && ~x23 )
						nx_state = s1;
					else nx_state = s1427;
				s1428 : if( x64 && x9 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x64 && x9 && ~x10 && x11 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x64 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x64 && ~x9 )
						nx_state = s1;
					else if( ~x64 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s604;
						end
					else nx_state = s1428;
				s1429 : if( x62 )
						begin
							y18 = 1'b1;	y48 = 1'b1;	
							nx_state = s1608;
						end
					else if( ~x62 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y56 = 1'b1;	
							nx_state = s1609;
						end
					else nx_state = s1429;
				s1430 : if( x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( ~x14 )
						nx_state = s1;
					else nx_state = s1430;
				s1431 : if( x7 && x19 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1564;
						end
					else if( x7 && ~x19 )
						begin
							y28 = 1'b1;	
							nx_state = s1565;
						end
					else if( ~x7 && x9 && x1 && x3 )
						begin
							y26 = 1'b1;	
							nx_state = s1197;
						end
					else if( ~x7 && x9 && x1 && ~x3 && x4 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s656;
						end
					else if( ~x7 && x9 && x1 && ~x3 && x4 && ~x5 && x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s653;
						end
					else if( ~x7 && x9 && x1 && ~x3 && x4 && ~x5 && ~x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x7 && x9 && x1 && ~x3 && ~x4 )
						begin
							y26 = 1'b1;	
							nx_state = s1197;
						end
					else if( ~x7 && x9 && ~x1 && x2 && x4 && x3 )
						begin
							y26 = 1'b1;	
							nx_state = s1468;
						end
					else if( ~x7 && x9 && ~x1 && x2 && x4 && ~x3 && x5 && x15 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x7 && x9 && ~x1 && x2 && x4 && ~x3 && x5 && ~x15 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x7 && x9 && ~x1 && x2 && x4 && ~x3 && x5 && ~x15 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x7 && x9 && ~x1 && x2 && x4 && ~x3 && x5 && ~x15 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( ~x7 && x9 && ~x1 && x2 && x4 && ~x3 && x5 && ~x15 && ~x22 )
						nx_state = s1;
					else if( ~x7 && x9 && ~x1 && x2 && x4 && ~x3 && ~x5 && x17 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x7 && x9 && ~x1 && x2 && x4 && ~x3 && ~x5 && ~x17 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x7 && x9 && ~x1 && x2 && x4 && ~x3 && ~x5 && ~x17 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x7 && x9 && ~x1 && x2 && x4 && ~x3 && ~x5 && ~x17 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( ~x7 && x9 && ~x1 && x2 && x4 && ~x3 && ~x5 && ~x17 && ~x22 )
						nx_state = s1;
					else if( ~x7 && x9 && ~x1 && x2 && ~x4 && x5 && x3 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1509;
						end
					else if( ~x7 && x9 && ~x1 && x2 && ~x4 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x7 && x9 && ~x1 && x2 && ~x4 && ~x5 && x3 && x16 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x7 && x9 && ~x1 && x2 && ~x4 && ~x5 && x3 && ~x16 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x7 && x9 && ~x1 && x2 && ~x4 && ~x5 && x3 && ~x16 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x7 && x9 && ~x1 && x2 && ~x4 && ~x5 && x3 && ~x16 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( ~x7 && x9 && ~x1 && x2 && ~x4 && ~x5 && x3 && ~x16 && ~x22 )
						nx_state = s1;
					else if( ~x7 && x9 && ~x1 && x2 && ~x4 && ~x5 && ~x3 )
						begin
							y38 = 1'b1;	
							nx_state = s845;
						end
					else if( ~x7 && x9 && ~x1 && ~x2 )
						begin
							y26 = 1'b1;	
							nx_state = s1197;
						end
					else if( ~x7 && ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y8 = 1'b1;	y32 = 1'b1;	
							nx_state = s1610;
						end
					else nx_state = s1431;
				s1432 : if( x20 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1611;
						end
					else if( ~x20 )
						begin
							y26 = 1'b1;	
							nx_state = s413;
						end
					else nx_state = s1432;
				s1433 : if( x22 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y29 = 1'b1;	y36 = 1'b1;	
							nx_state = s1541;
						end
					else if( x22 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1089;
						end
					else if( ~x22 && x23 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s1339;
						end
					else if( ~x22 && x23 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1089;
						end
					else if( ~x22 && ~x23 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s1092;
						end
					else if( ~x22 && ~x23 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1088;
						end
					else nx_state = s1433;
				s1434 : if( x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s1086;
						end
					else if( ~x17 && x22 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1090;
						end
					else if( ~x17 && ~x22 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1091;
						end
					else nx_state = s1434;
				s1435 : if( x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s1339;
						end
					else if( ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1091;
						end
					else nx_state = s1435;
				s1436 : if( x10 && x18 && x2 && x19 && x4 && x3 && x5 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1612;
						end
					else if( x10 && x18 && x2 && x19 && x4 && x3 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1612;
						end
					else if( x10 && x18 && x2 && x19 && x4 && x3 && ~x5 && ~x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y21 = 1'b1;	
							y32 = 1'b1;	y35 = 1'b1;	
							nx_state = s1500;
						end
					else if( x10 && x18 && x2 && x19 && x4 && ~x3 && x17 && x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s820;
						end
					else if( x10 && x18 && x2 && x19 && x4 && ~x3 && x17 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s821;
						end
					else if( x10 && x18 && x2 && x19 && x4 && ~x3 && x17 && ~x5 && ~x6 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( x10 && x18 && x2 && x19 && x4 && ~x3 && ~x17 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x10 && x18 && x2 && x19 && x4 && ~x3 && ~x17 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x10 && x18 && x2 && x19 && x4 && ~x3 && ~x17 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x10 && x18 && x2 && x19 && x4 && ~x3 && ~x17 && ~x11 )
						nx_state = s1;
					else if( x10 && x18 && x2 && x19 && ~x4 && x3 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y19 = 1'b1;	
							nx_state = s872;
						end
					else if( x10 && x18 && x2 && x19 && ~x4 && ~x3 && x16 && x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s820;
						end
					else if( x10 && x18 && x2 && x19 && ~x4 && ~x3 && x16 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s821;
						end
					else if( x10 && x18 && x2 && x19 && ~x4 && ~x3 && x16 && ~x5 && ~x6 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( x10 && x18 && x2 && x19 && ~x4 && ~x3 && ~x16 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x10 && x18 && x2 && x19 && ~x4 && ~x3 && ~x16 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x10 && x18 && x2 && x19 && ~x4 && ~x3 && ~x16 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x10 && x18 && x2 && x19 && ~x4 && ~x3 && ~x16 && ~x11 )
						nx_state = s1;
					else if( x10 && x18 && x2 && ~x19 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x10 && x18 && x2 && ~x19 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x10 && x18 && x2 && ~x19 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x10 && x18 && x2 && ~x19 && ~x11 )
						nx_state = s1;
					else if( x10 && x18 && ~x2 && x3 && x19 && x4 && x15 && x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s820;
						end
					else if( x10 && x18 && ~x2 && x3 && x19 && x4 && x15 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s821;
						end
					else if( x10 && x18 && ~x2 && x3 && x19 && x4 && x15 && ~x5 && ~x6 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( x10 && x18 && ~x2 && x3 && x19 && x4 && ~x15 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x10 && x18 && ~x2 && x3 && x19 && x4 && ~x15 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x10 && x18 && ~x2 && x3 && x19 && x4 && ~x15 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x10 && x18 && ~x2 && x3 && x19 && x4 && ~x15 && ~x11 )
						nx_state = s1;
					else if( x10 && x18 && ~x2 && x3 && x19 && ~x4 && x14 && x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s820;
						end
					else if( x10 && x18 && ~x2 && x3 && x19 && ~x4 && x14 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s821;
						end
					else if( x10 && x18 && ~x2 && x3 && x19 && ~x4 && x14 && ~x5 && ~x6 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( x10 && x18 && ~x2 && x3 && x19 && ~x4 && ~x14 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x10 && x18 && ~x2 && x3 && x19 && ~x4 && ~x14 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x10 && x18 && ~x2 && x3 && x19 && ~x4 && ~x14 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x10 && x18 && ~x2 && x3 && x19 && ~x4 && ~x14 && ~x11 )
						nx_state = s1;
					else if( x10 && x18 && ~x2 && x3 && ~x19 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x10 && x18 && ~x2 && x3 && ~x19 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x10 && x18 && ~x2 && x3 && ~x19 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x10 && x18 && ~x2 && x3 && ~x19 && ~x11 )
						nx_state = s1;
					else if( x10 && x18 && ~x2 && ~x3 && x19 && x4 && x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s820;
						end
					else if( x10 && x18 && ~x2 && ~x3 && x19 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s821;
						end
					else if( x10 && x18 && ~x2 && ~x3 && x19 && x4 && ~x5 && ~x6 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( x10 && x18 && ~x2 && ~x3 && x19 && ~x4 )
						begin
							y47 = 1'b1;	
							nx_state = s287;
						end
					else if( x10 && x18 && ~x2 && ~x3 && ~x19 && x4 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1612;
						end
					else if( x10 && x18 && ~x2 && ~x3 && ~x19 && ~x4 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s1321;
						end
					else if( x10 && ~x18 && x19 && x2 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1612;
						end
					else if( x10 && ~x18 && x19 && ~x2 && x4 && x3 )
						begin
							y23 = 1'b1;	y27 = 1'b1;	y48 = 1'b1;	
							nx_state = s1613;
						end
					else if( x10 && ~x18 && x19 && ~x2 && x4 && ~x3 )
						begin
							y37 = 1'b1;	
							nx_state = s888;
						end
					else if( x10 && ~x18 && x19 && ~x2 && ~x4 && x3 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s79;
						end
					else if( x10 && ~x18 && x19 && ~x2 && ~x4 && ~x3 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1093;
						end
					else if( x10 && ~x18 && ~x19 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1612;
						end
					else if( ~x10 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							y30 = 1'b1;	y35 = 1'b1;	y51 = 1'b1;	
							nx_state = s1499;
						end
					else nx_state = s1436;
				s1437 : if( 1'b1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y20 = 1'b1;	
							nx_state = s1095;
						end
					else nx_state = s1437;
				s1438 : if( x63 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s1614;
						end
					else if( ~x63 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x63 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x63 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x63 && ~x8 )
						nx_state = s1;
					else nx_state = s1438;
				s1439 : if( x66 && x9 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s1615;
						end
					else if( x66 && ~x9 && x19 && x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s1616;
						end
					else if( x66 && ~x9 && x19 && ~x4 && x5 && x6 && x7 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s1617;
						end
					else if( x66 && ~x9 && x19 && ~x4 && x5 && x6 && ~x7 )
						begin
							y3 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	y30 = 1'b1;	
							nx_state = s1618;
						end
					else if( x66 && ~x9 && x19 && ~x4 && x5 && ~x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1571;
						end
					else if( x66 && ~x9 && x19 && ~x4 && ~x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s1619;
						end
					else if( x66 && ~x9 && ~x19 )
						begin
							y4 = 1'b1;	y20 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s1620;
						end
					else if( ~x66 )
						begin
							y6 = 1'b1;	
							nx_state = s310;
						end
					else nx_state = s1439;
				s1440 : if( 1'b1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y5 = 1'b1;	
							y22 = 1'b1;	y23 = 1'b1;	
							nx_state = s72;
						end
					else nx_state = s1440;
				s1441 : if( x64 && x3 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1263;
						end
					else if( x64 && ~x3 )
						begin
							y3 = 1'b1;	y6 = 1'b1;	y12 = 1'b1;	
							y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s1621;
						end
					else if( ~x64 && x14 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x64 && x14 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x64 && x14 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x64 && x14 && ~x23 )
						nx_state = s1;
					else if( ~x64 && ~x14 )
						begin
							y47 = 1'b1;	y56 = 1'b1;	y61 = 1'b1;	
							y70 = 1'b1;	
							nx_state = s1514;
						end
					else nx_state = s1441;
				s1442 : if( 1'b1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y8 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1622;
						end
					else nx_state = s1442;
				s1443 : if( x11 && x10 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s1478;
						end
					else if( x11 && ~x10 )
						begin
							y28 = 1'b1;	
							nx_state = s991;
						end
					else if( ~x11 )
						begin
							y29 = 1'b1;	
							nx_state = s1109;
						end
					else nx_state = s1443;
				s1444 : if( x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1623;
						end
					else if( ~x3 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y25 = 1'b1;	
							y30 = 1'b1;	y31 = 1'b1;	y32 = 1'b1;	
							nx_state = s1624;
						end
					else nx_state = s1444;
				s1445 : if( x62 )
						begin
							y29 = 1'b1;	
							nx_state = s771;
						end
					else if( ~x62 )
						begin
							y15 = 1'b1;	
							nx_state = s1625;
						end
					else nx_state = s1445;
				s1446 : if( 1'b1 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s1626;
						end
					else nx_state = s1446;
				s1447 : if( x3 && x21 && x26 && x27 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x3 && x21 && x26 && x27 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x3 && x21 && x26 && x27 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x3 && x21 && x26 && x27 && x22 && ~x23 )
						nx_state = s1;
					else if( x3 && x21 && x26 && x27 && ~x22 )
						nx_state = s1;
					else if( x3 && x21 && x26 && ~x27 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1627;
						end
					else if( x3 && x21 && ~x26 && x7 && x8 && x6 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x3 && x21 && ~x26 && x7 && x8 && x6 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x3 && x21 && ~x26 && x7 && x8 && x6 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x3 && x21 && ~x26 && x7 && x8 && x6 && x22 && ~x23 )
						nx_state = s1;
					else if( x3 && x21 && ~x26 && x7 && x8 && x6 && ~x22 )
						nx_state = s1;
					else if( x3 && x21 && ~x26 && x7 && x8 && ~x6 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( x3 && x21 && ~x26 && x7 && x8 && ~x6 && ~x9 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x3 && x21 && ~x26 && x7 && x8 && ~x6 && ~x9 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x3 && x21 && ~x26 && x7 && x8 && ~x6 && ~x9 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x3 && x21 && ~x26 && x7 && x8 && ~x6 && ~x9 && x22 && ~x23 )
						nx_state = s1;
					else if( x3 && x21 && ~x26 && x7 && x8 && ~x6 && ~x9 && ~x22 )
						nx_state = s1;
					else if( x3 && x21 && ~x26 && x7 && ~x8 && x6 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( x3 && x21 && ~x26 && x7 && ~x8 && ~x6 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( x3 && x21 && ~x26 && x7 && ~x8 && ~x6 && ~x10 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x3 && x21 && ~x26 && x7 && ~x8 && ~x6 && ~x10 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x3 && x21 && ~x26 && x7 && ~x8 && ~x6 && ~x10 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x3 && x21 && ~x26 && x7 && ~x8 && ~x6 && ~x10 && x22 && ~x23 )
						nx_state = s1;
					else if( x3 && x21 && ~x26 && x7 && ~x8 && ~x6 && ~x10 && ~x22 )
						nx_state = s1;
					else if( x3 && x21 && ~x26 && ~x7 && x8 && x6 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y42 = 1'b1;	
							nx_state = s1628;
						end
					else if( x3 && x21 && ~x26 && ~x7 && x8 && ~x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( x3 && x21 && ~x26 && ~x7 && ~x8 && x6 && x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( x3 && x21 && ~x26 && ~x7 && ~x8 && x6 && ~x11 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x3 && x21 && ~x26 && ~x7 && ~x8 && x6 && ~x11 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x3 && x21 && ~x26 && ~x7 && ~x8 && x6 && ~x11 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x3 && x21 && ~x26 && ~x7 && ~x8 && x6 && ~x11 && x22 && ~x23 )
						nx_state = s1;
					else if( x3 && x21 && ~x26 && ~x7 && ~x8 && x6 && ~x11 && ~x22 )
						nx_state = s1;
					else if( x3 && x21 && ~x26 && ~x7 && ~x8 && ~x6 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( x3 && ~x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y28 = 1'b1;	y29 = 1'b1;	
							nx_state = s1629;
						end
					else if( ~x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y16 = 1'b1;	y24 = 1'b1;	
							nx_state = s1630;
						end
					else nx_state = s1447;
				s1448 : if( x26 && x27 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s1631;
						end
					else if( x26 && ~x27 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1627;
						end
					else if( ~x26 && x12 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x26 && ~x12 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x26 && ~x12 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x26 && ~x12 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x26 && ~x12 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x26 && ~x12 && ~x22 )
						nx_state = s1;
					else nx_state = s1448;
				s1449 : if( x13 )
						begin
							y61 = 1'b1;	
							nx_state = s1098;
						end
					else if( ~x13 && x26 && x14 && x27 && x6 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s1448;
						end
					else if( ~x13 && x26 && x14 && x27 && x6 && ~x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s677;
						end
					else if( ~x13 && x26 && x14 && x27 && ~x6 && x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s1447;
						end
					else if( ~x13 && x26 && x14 && x27 && ~x6 && ~x5 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							nx_state = s1199;
						end
					else if( ~x13 && x26 && x14 && ~x27 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s1220;
						end
					else if( ~x13 && x26 && x14 && ~x27 && ~x5 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							nx_state = s1199;
						end
					else if( ~x13 && x26 && ~x14 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s1448;
						end
					else if( ~x13 && x26 && ~x14 && ~x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s677;
						end
					else if( ~x13 && ~x26 && x27 && x14 && x5 )
						begin
							y50 = 1'b1;	
							nx_state = s658;
						end
					else if( ~x13 && ~x26 && x27 && x14 && ~x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s1447;
						end
					else if( ~x13 && ~x26 && x27 && ~x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s1448;
						end
					else if( ~x13 && ~x26 && ~x27 && x7 && x6 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x13 && ~x26 && ~x27 && x7 && x6 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x13 && ~x26 && ~x27 && x7 && x6 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x13 && ~x26 && ~x27 && x7 && x6 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x13 && ~x26 && ~x27 && x7 && x6 && ~x22 )
						nx_state = s1;
					else if( ~x13 && ~x26 && ~x27 && x7 && ~x6 && x8 && x15 )
						begin
							y10 = 1'b1;	
							nx_state = s405;
						end
					else if( ~x13 && ~x26 && ~x27 && x7 && ~x6 && x8 && ~x15 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x13 && ~x26 && ~x27 && x7 && ~x6 && x8 && ~x15 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x13 && ~x26 && ~x27 && x7 && ~x6 && x8 && ~x15 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x13 && ~x26 && ~x27 && x7 && ~x6 && x8 && ~x15 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x13 && ~x26 && ~x27 && x7 && ~x6 && x8 && ~x15 && ~x22 )
						nx_state = s1;
					else if( ~x13 && ~x26 && ~x27 && x7 && ~x6 && ~x8 && x16 )
						begin
							y10 = 1'b1;	
							nx_state = s405;
						end
					else if( ~x13 && ~x26 && ~x27 && x7 && ~x6 && ~x8 && ~x16 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x13 && ~x26 && ~x27 && x7 && ~x6 && ~x8 && ~x16 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x13 && ~x26 && ~x27 && x7 && ~x6 && ~x8 && ~x16 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x13 && ~x26 && ~x27 && x7 && ~x6 && ~x8 && ~x16 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x13 && ~x26 && ~x27 && x7 && ~x6 && ~x8 && ~x16 && ~x22 )
						nx_state = s1;
					else if( ~x13 && ~x26 && ~x27 && ~x7 && x8 && x6 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x13 && ~x26 && ~x27 && ~x7 && x8 && ~x6 )
						begin
							y5 = 1'b1;	y44 = 1'b1;	y55 = 1'b1;	
							y60 = 1'b1;	
							nx_state = s1220;
						end
					else if( ~x13 && ~x26 && ~x27 && ~x7 && ~x8 && x6 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x13 && ~x26 && ~x27 && ~x7 && ~x8 && ~x6 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y53 = 1'b1;	
							y54 = 1'b1;	
							nx_state = s1220;
						end
					else nx_state = s1449;
				s1450 : if( 1'b1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y23 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s1632;
						end
					else nx_state = s1450;
				s1451 : if( 1'b1 )
						begin
							y80 = 1'b1;	
							nx_state = s1568;
						end
					else nx_state = s1451;
				s1452 : if( 1'b1 )
						begin
							y80 = 1'b1;	
							nx_state = s1633;
						end
					else nx_state = s1452;
				s1453 : if( x15 )
						begin
							y44 = 1'b1;	y45 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x15 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x15 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x15 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x15 && ~x6 )
						nx_state = s1;
					else nx_state = s1453;
				s1454 : if( 1'b1 )
						begin
							y19 = 1'b1;	y24 = 1'b1;	y26 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s1454;
				s1455 : if( x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x19 )
						nx_state = s1;
					else nx_state = s1455;
				s1456 : if( x6 )
						begin
							y4 = 1'b1;	y12 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1634;
						end
					else if( ~x6 && x14 && x7 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1635;
						end
					else if( ~x6 && x14 && ~x7 && x5 && x10 && x9 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1636;
						end
					else if( ~x6 && x14 && ~x7 && x5 && x10 && ~x9 && x11 && x16 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1455;
						end
					else if( ~x6 && x14 && ~x7 && x5 && x10 && ~x9 && x11 && ~x16 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x6 && x14 && ~x7 && x5 && x10 && ~x9 && x11 && ~x16 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x6 && x14 && ~x7 && x5 && x10 && ~x9 && x11 && ~x16 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x6 && x14 && ~x7 && x5 && x10 && ~x9 && x11 && ~x16 && ~x19 )
						nx_state = s1;
					else if( ~x6 && x14 && ~x7 && x5 && x10 && ~x9 && ~x11 && x17 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1455;
						end
					else if( ~x6 && x14 && ~x7 && x5 && x10 && ~x9 && ~x11 && ~x17 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x6 && x14 && ~x7 && x5 && x10 && ~x9 && ~x11 && ~x17 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x6 && x14 && ~x7 && x5 && x10 && ~x9 && ~x11 && ~x17 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x6 && x14 && ~x7 && x5 && x10 && ~x9 && ~x11 && ~x17 && ~x19 )
						nx_state = s1;
					else if( ~x6 && x14 && ~x7 && x5 && ~x10 && x11 && x9 )
						begin
							y6 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s80;
						end
					else if( ~x6 && x14 && ~x7 && x5 && ~x10 && x11 && ~x9 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1455;
						end
					else if( ~x6 && x14 && ~x7 && x5 && ~x10 && ~x11 && x9 && x15 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1455;
						end
					else if( ~x6 && x14 && ~x7 && x5 && ~x10 && ~x11 && x9 && ~x15 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x6 && x14 && ~x7 && x5 && ~x10 && ~x11 && x9 && ~x15 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x6 && x14 && ~x7 && x5 && ~x10 && ~x11 && x9 && ~x15 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x6 && x14 && ~x7 && x5 && ~x10 && ~x11 && x9 && ~x15 && ~x19 )
						nx_state = s1;
					else if( ~x6 && x14 && ~x7 && x5 && ~x10 && ~x11 && ~x9 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x6 && x14 && ~x7 && ~x5 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1637;
						end
					else if( ~x6 && ~x14 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s1638;
						end
					else nx_state = s1456;
				s1457 : if( x4 )
						begin
							y23 = 1'b1;	
							nx_state = s588;
						end
					else if( ~x4 && x5 && x7 && x9 && x11 )
						begin
							y26 = 1'b1;	
							nx_state = s262;
						end
					else if( ~x4 && x5 && x7 && x9 && ~x11 )
						begin
							y28 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x4 && x5 && x7 && ~x9 && x10 && x11 && x12 )
						begin
							y19 = 1'b1;	
							nx_state = s404;
						end
					else if( ~x4 && x5 && x7 && ~x9 && x10 && x11 && ~x12 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x4 && x5 && x7 && ~x9 && x10 && x11 && ~x12 && x19 && ~x13 )
						nx_state = s1;
					else if( ~x4 && x5 && x7 && ~x9 && x10 && x11 && ~x12 && ~x19 )
						nx_state = s1;
					else if( ~x4 && x5 && x7 && ~x9 && x10 && ~x11 && x13 )
						begin
							y19 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x4 && x5 && x7 && ~x9 && x10 && ~x11 && ~x13 && x19 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x4 && x5 && x7 && ~x9 && x10 && ~x11 && ~x13 && x19 && ~x12 )
						nx_state = s1;
					else if( ~x4 && x5 && x7 && ~x9 && x10 && ~x11 && ~x13 && ~x19 )
						nx_state = s1;
					else if( ~x4 && x5 && x7 && ~x9 && ~x10 && x11 )
						begin
							y5 = 1'b1;	y18 = 1'b1;	y27 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s1455;
						end
					else if( ~x4 && x5 && x7 && ~x9 && ~x10 && ~x11 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1455;
						end
					else if( ~x4 && x5 && ~x7 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1638;
						end
					else if( ~x4 && ~x5 && x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1638;
						end
					else if( ~x4 && ~x5 && ~x6 && x9 && x10 && x11 && x7 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x4 && ~x5 && ~x6 && x9 && x10 && x11 && ~x7 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	y16 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1639;
						end
					else if( ~x4 && ~x5 && ~x6 && x9 && x10 && ~x11 && x7 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x4 && ~x5 && ~x6 && x9 && x10 && ~x11 && ~x7 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y50 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s1640;
						end
					else if( ~x4 && ~x5 && ~x6 && x9 && ~x10 && x11 && x7 )
						begin
							y25 = 1'b1;	
							nx_state = s1641;
						end
					else if( ~x4 && ~x5 && ~x6 && x9 && ~x10 && x11 && ~x7 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y46 = 1'b1;	
							y47 = 1'b1;	
							nx_state = s1642;
						end
					else if( ~x4 && ~x5 && ~x6 && x9 && ~x10 && ~x11 && x7 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1455;
						end
					else if( ~x4 && ~x5 && ~x6 && x9 && ~x10 && ~x11 && ~x7 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y52 = 1'b1;	
							y53 = 1'b1;	
							nx_state = s1643;
						end
					else if( ~x4 && ~x5 && ~x6 && ~x9 && x10 && x11 && x7 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s1644;
						end
					else if( ~x4 && ~x5 && ~x6 && ~x9 && x10 && x11 && ~x7 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s1455;
						end
					else if( ~x4 && ~x5 && ~x6 && ~x9 && x10 && ~x11 && x7 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y34 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s1455;
						end
					else if( ~x4 && ~x5 && ~x6 && ~x9 && x10 && ~x11 && ~x7 )
						begin
							y17 = 1'b1;	y18 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	y37 = 1'b1;	
							nx_state = s1455;
						end
					else if( ~x4 && ~x5 && ~x6 && ~x9 && ~x10 && x7 && x11 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1455;
						end
					else if( ~x4 && ~x5 && ~x6 && ~x9 && ~x10 && x7 && ~x11 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s575;
						end
					else if( ~x4 && ~x5 && ~x6 && ~x9 && ~x10 && ~x7 )
						begin
							y11 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							y33 = 1'b1;	y34 = 1'b1;	
							nx_state = s1455;
						end
					else nx_state = s1457;
				s1458 : if( 1'b1 )
						begin
							y15 = 1'b1;	
							nx_state = s1645;
						end
					else nx_state = s1458;
				s1459 : if( x9 && x17 && x19 && x20 && x14 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else if( x9 && x17 && x19 && x20 && ~x14 )
						begin
							y4 = 1'b1;	y29 = 1'b1;	y32 = 1'b1;	
							nx_state = s863;
						end
					else if( x9 && x17 && x19 && ~x20 && x14 )
						begin
							y4 = 1'b1;	y18 = 1'b1;	y29 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s863;
						end
					else if( x9 && x17 && x19 && ~x20 && ~x14 && x16 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	y32 = 1'b1;	
							nx_state = s863;
						end
					else if( x9 && x17 && x19 && ~x20 && ~x14 && ~x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s863;
						end
					else if( x9 && x17 && ~x19 && x16 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s863;
						end
					else if( x9 && x17 && ~x19 && ~x16 && x20 )
						begin
							y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s863;
						end
					else if( x9 && x17 && ~x19 && ~x16 && ~x20 && x15 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s364;
						end
					else if( x9 && x17 && ~x19 && ~x16 && ~x20 && ~x15 )
						begin
							y25 = 1'b1;	
							nx_state = s148;
						end
					else if( x9 && ~x17 && x18 && x19 && x14 && x16 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	y19 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s861;
						end
					else if( x9 && ~x17 && x18 && x19 && x14 && ~x16 )
						begin
							y2 = 1'b1;	y21 = 1'b1;	
							nx_state = s1318;
						end
					else if( x9 && ~x17 && x18 && x19 && ~x14 )
						begin
							y7 = 1'b1;	
							nx_state = s747;
						end
					else if( x9 && ~x17 && x18 && ~x19 )
						begin
							y7 = 1'b1;	
							nx_state = s747;
						end
					else if( x9 && ~x17 && ~x18 )
						begin
							y4 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x9 && x19 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s868;
						end
					else if( ~x9 && ~x19 && x20 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s868;
						end
					else if( ~x9 && ~x19 && ~x20 && x17 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s868;
						end
					else if( ~x9 && ~x19 && ~x20 && ~x17 && x18 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s548;
						end
					else if( ~x9 && ~x19 && ~x20 && ~x17 && ~x18 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s868;
						end
					else nx_state = s1459;
				s1460 : if( 1'b1 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y39 = 1'b1;	
							nx_state = s584;
						end
					else nx_state = s1460;
				s1461 : if( 1'b1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y37 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s1646;
						end
					else nx_state = s1461;
				s1462 : if( 1'b1 )
						begin
							y47 = 1'b1;	y53 = 1'b1;	y61 = 1'b1;	
							y71 = 1'b1;	
							nx_state = s1554;
						end
					else nx_state = s1462;
				s1463 : if( 1'b1 )
						begin
							y40 = 1'b1;	
							nx_state = s1647;
						end
					else nx_state = s1463;
				s1464 : if( 1'b1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y37 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s584;
						end
					else nx_state = s1464;
				s1465 : if( 1'b1 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y39 = 1'b1;	
							nx_state = s584;
						end
					else nx_state = s1465;
				s1466 : if( 1'b1 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y39 = 1'b1;	
							nx_state = s584;
						end
					else nx_state = s1466;
				s1467 : if( x30 )
						begin
							y5 = 1'b1;	
							nx_state = s560;
						end
					else if( ~x30 )
						begin
							y5 = 1'b1;	
							nx_state = s66;
						end
					else nx_state = s1467;
				s1468 : if( x63 )
						begin
							y27 = 1'b1;	
							nx_state = s648;
						end
					else if( ~x63 && x64 )
						begin
							y5 = 1'b1;	y13 = 1'b1;	y17 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1648;
						end
					else if( ~x63 && ~x64 )
						begin
							y41 = 1'b1;	
							nx_state = s1649;
						end
					else nx_state = s1468;
				s1469 : if( 1'b1 )
						begin
							y6 = 1'b1;	y19 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1650;
						end
					else nx_state = s1469;
				s1470 : if( x4 )
						begin
							y15 = 1'b1;	
							nx_state = s1544;
						end
					else if( ~x4 )
						begin
							y6 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s1651;
						end
					else nx_state = s1470;
				s1471 : if( 1'b1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s597;
						end
					else nx_state = s1471;
				s1472 : if( 1'b1 )
						begin
							y6 = 1'b1;	
							nx_state = s1049;
						end
					else nx_state = s1472;
				s1473 : if( 1'b1 )
						begin
							y38 = 1'b1;	
							nx_state = s1503;
						end
					else nx_state = s1473;
				s1474 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1627;
						end
					else nx_state = s1474;
				s1475 : if( 1'b1 )
						begin
							y6 = 1'b1;	y11 = 1'b1;	y40 = 1'b1;	
							y41 = 1'b1;	y42 = 1'b1;	y45 = 1'b1;	
							nx_state = s1652;
						end
					else nx_state = s1475;
				s1476 : if( 1'b1 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s1014;
						end
					else nx_state = s1476;
				s1477 : if( 1'b1 )
						begin
							y3 = 1'b1;	y77 = 1'b1;	
							nx_state = s1133;
						end
					else nx_state = s1477;
				s1478 : if( 1'b1 )
						begin
							y53 = 1'b1;	
							nx_state = s1424;
						end
					else nx_state = s1478;
				s1479 : if( 1'b1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							nx_state = s1653;
						end
					else nx_state = s1479;
				s1480 : if( x3 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1654;
						end
					else if( ~x3 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							y16 = 1'b1;	y18 = 1'b1;	y25 = 1'b1;	
							nx_state = s662;
						end
					else nx_state = s1480;
				s1481 : if( x8 && x20 && x14 && x15 )
						begin
							y6 = 1'b1;	y11 = 1'b1;	y26 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1307;
						end
					else if( x8 && x20 && x14 && ~x15 )
						begin
							y6 = 1'b1;	y11 = 1'b1;	y42 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1068;
						end
					else if( x8 && x20 && ~x14 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y44 = 1'b1;	
							y45 = 1'b1;	y49 = 1'b1;	
							nx_state = s1482;
						end
					else if( x8 && ~x20 && x13 && x21 && x14 && x15 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else if( x8 && ~x20 && x13 && x21 && x14 && ~x15 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( x8 && ~x20 && x13 && x21 && x14 && ~x15 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( x8 && ~x20 && x13 && x21 && ~x14 && x15 && x17 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( x8 && ~x20 && x13 && x21 && ~x14 && x15 && x17 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( x8 && ~x20 && x13 && x21 && ~x14 && x15 && ~x17 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x8 && ~x20 && x13 && x21 && ~x14 && x15 && ~x17 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x8 && ~x20 && x13 && x21 && ~x14 && x15 && ~x17 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x8 && ~x20 && x13 && x21 && ~x14 && x15 && ~x17 && ~x10 )
						nx_state = s1;
					else if( x8 && ~x20 && x13 && x21 && ~x14 && ~x15 && x9 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( x8 && ~x20 && x13 && x21 && ~x14 && ~x15 && x9 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( x8 && ~x20 && x13 && x21 && ~x14 && ~x15 && ~x9 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x8 && ~x20 && x13 && x21 && ~x14 && ~x15 && ~x9 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x8 && ~x20 && x13 && x21 && ~x14 && ~x15 && ~x9 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x8 && ~x20 && x13 && x21 && ~x14 && ~x15 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x8 && ~x20 && x13 && ~x21 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							nx_state = s1213;
						end
					else if( x8 && ~x20 && ~x13 && x14 && x21 && x15 && x18 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( x8 && ~x20 && ~x13 && x14 && x21 && x15 && x18 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( x8 && ~x20 && ~x13 && x14 && x21 && x15 && ~x18 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x8 && ~x20 && ~x13 && x14 && x21 && x15 && ~x18 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x8 && ~x20 && ~x13 && x14 && x21 && x15 && ~x18 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x8 && ~x20 && ~x13 && x14 && x21 && x15 && ~x18 && ~x10 )
						nx_state = s1;
					else if( x8 && ~x20 && ~x13 && x14 && x21 && ~x15 && x19 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( x8 && ~x20 && ~x13 && x14 && x21 && ~x15 && x19 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( x8 && ~x20 && ~x13 && x14 && x21 && ~x15 && ~x19 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x8 && ~x20 && ~x13 && x14 && x21 && ~x15 && ~x19 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x8 && ~x20 && ~x13 && x14 && x21 && ~x15 && ~x19 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x8 && ~x20 && ~x13 && x14 && x21 && ~x15 && ~x19 && ~x10 )
						nx_state = s1;
					else if( x8 && ~x20 && ~x13 && x14 && ~x21 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y22 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s722;
						end
					else if( x8 && ~x20 && ~x13 && ~x14 && x21 && x15 && x5 )
						begin
							y14 = 1'b1;	
							nx_state = s5;
						end
					else if( x8 && ~x20 && ~x13 && ~x14 && x21 && x15 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1207;
						end
					else if( x8 && ~x20 && ~x13 && ~x14 && x21 && ~x15 && x7 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1208;
						end
					else if( x8 && ~x20 && ~x13 && ~x14 && x21 && ~x15 && ~x7 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1209;
						end
					else if( x8 && ~x20 && ~x13 && ~x14 && ~x21 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x8 && ~x20 && ~x13 && ~x14 && ~x21 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x8 && ~x20 && ~x13 && ~x14 && ~x21 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x8 && ~x20 && ~x13 && ~x14 && ~x21 && ~x10 )
						nx_state = s1;
					else if( ~x8 )
						begin
							y6 = 1'b1;	y9 = 1'b1;	y25 = 1'b1;	
							y56 = 1'b1;	
							nx_state = s1483;
						end
					else nx_state = s1481;
				s1482 : if( 1'b1 )
						begin
							y11 = 1'b1;	y41 = 1'b1;	y45 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s1655;
						end
					else nx_state = s1482;
				s1483 : if( x9 )
						begin
							y15 = 1'b1;	
							nx_state = s1141;
						end
					else if( ~x9 && x20 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s1656;
						end
					else if( ~x9 && ~x20 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s1484;
						end
					else nx_state = s1483;
				s1484 : if( x20 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1657;
						end
					else if( ~x20 )
						begin
							y6 = 1'b1;	y9 = 1'b1;	y25 = 1'b1;	
							y56 = 1'b1;	
							nx_state = s1512;
						end
					else nx_state = s1484;
				s1485 : if( x20 && x14 && x15 )
						begin
							y6 = 1'b1;	y11 = 1'b1;	y26 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1307;
						end
					else if( x20 && x14 && ~x15 )
						begin
							y6 = 1'b1;	y11 = 1'b1;	y42 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1068;
						end
					else if( x20 && ~x14 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y44 = 1'b1;	
							y45 = 1'b1;	y49 = 1'b1;	
							nx_state = s1482;
						end
					else if( ~x20 && x21 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1658;
						end
					else if( ~x20 && ~x21 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1657;
						end
					else nx_state = s1485;
				s1486 : if( 1'b1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s1659;
						end
					else nx_state = s1486;
				s1487 : if( 1'b1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s1660;
						end
					else nx_state = s1487;
				s1488 : if( 1'b1 )
						begin
							y29 = 1'b1;	
							nx_state = s1661;
						end
					else nx_state = s1488;
				s1489 : if( 1'b1 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							nx_state = s1213;
						end
					else nx_state = s1489;
				s1490 : if( 1'b1 )
						begin
							y7 = 1'b1;	y39 = 1'b1;	y49 = 1'b1;	
							nx_state = s1662;
						end
					else nx_state = s1490;
				s1491 : if( 1'b1 )
						begin
							y5 = 1'b1;	y42 = 1'b1;	y43 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s1663;
						end
					else nx_state = s1491;
				s1492 : if( 1'b1 )
						begin
							y33 = 1'b1;	
							nx_state = s1033;
						end
					else nx_state = s1492;
				s1493 : if( 1'b1 )
						begin
							y9 = 1'b1;	
							nx_state = s967;
						end
					else nx_state = s1493;
				s1494 : if( 1'b1 )
						begin
							y9 = 1'b1;	
							nx_state = s790;
						end
					else nx_state = s1494;
				s1495 : if( 1'b1 )
						begin
							y9 = 1'b1;	
							nx_state = s1664;
						end
					else nx_state = s1495;
				s1496 : if( 1'b1 )
						begin
							y9 = 1'b1;	
							nx_state = s1665;
						end
					else nx_state = s1496;
				s1497 : if( 1'b1 )
						begin
							y9 = 1'b1;	
							nx_state = s1666;
						end
					else nx_state = s1497;
				s1498 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s1225;
						end
					else nx_state = s1498;
				s1499 : if( x18 && x2 && x19 && x4 && x3 && x5 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1612;
						end
					else if( x18 && x2 && x19 && x4 && x3 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1612;
						end
					else if( x18 && x2 && x19 && x4 && x3 && ~x5 && ~x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y21 = 1'b1;	
							y32 = 1'b1;	y35 = 1'b1;	
							nx_state = s1500;
						end
					else if( x18 && x2 && x19 && x4 && ~x3 && x17 && x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s820;
						end
					else if( x18 && x2 && x19 && x4 && ~x3 && x17 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s821;
						end
					else if( x18 && x2 && x19 && x4 && ~x3 && x17 && ~x5 && ~x6 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( x18 && x2 && x19 && x4 && ~x3 && ~x17 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x18 && x2 && x19 && x4 && ~x3 && ~x17 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x18 && x2 && x19 && x4 && ~x3 && ~x17 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x18 && x2 && x19 && x4 && ~x3 && ~x17 && ~x11 )
						nx_state = s1;
					else if( x18 && x2 && x19 && ~x4 && x3 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y19 = 1'b1;	
							nx_state = s872;
						end
					else if( x18 && x2 && x19 && ~x4 && ~x3 && x16 && x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s820;
						end
					else if( x18 && x2 && x19 && ~x4 && ~x3 && x16 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s821;
						end
					else if( x18 && x2 && x19 && ~x4 && ~x3 && x16 && ~x5 && ~x6 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( x18 && x2 && x19 && ~x4 && ~x3 && ~x16 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x18 && x2 && x19 && ~x4 && ~x3 && ~x16 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x18 && x2 && x19 && ~x4 && ~x3 && ~x16 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x18 && x2 && x19 && ~x4 && ~x3 && ~x16 && ~x11 )
						nx_state = s1;
					else if( x18 && x2 && ~x19 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x18 && x2 && ~x19 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x18 && x2 && ~x19 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x18 && x2 && ~x19 && ~x11 )
						nx_state = s1;
					else if( x18 && ~x2 && x3 && x19 && x4 && x15 && x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s820;
						end
					else if( x18 && ~x2 && x3 && x19 && x4 && x15 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s821;
						end
					else if( x18 && ~x2 && x3 && x19 && x4 && x15 && ~x5 && ~x6 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( x18 && ~x2 && x3 && x19 && x4 && ~x15 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x18 && ~x2 && x3 && x19 && x4 && ~x15 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x18 && ~x2 && x3 && x19 && x4 && ~x15 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x18 && ~x2 && x3 && x19 && x4 && ~x15 && ~x11 )
						nx_state = s1;
					else if( x18 && ~x2 && x3 && x19 && ~x4 && x14 && x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s820;
						end
					else if( x18 && ~x2 && x3 && x19 && ~x4 && x14 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s821;
						end
					else if( x18 && ~x2 && x3 && x19 && ~x4 && x14 && ~x5 && ~x6 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( x18 && ~x2 && x3 && x19 && ~x4 && ~x14 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x18 && ~x2 && x3 && x19 && ~x4 && ~x14 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x18 && ~x2 && x3 && x19 && ~x4 && ~x14 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x18 && ~x2 && x3 && x19 && ~x4 && ~x14 && ~x11 )
						nx_state = s1;
					else if( x18 && ~x2 && x3 && ~x19 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x18 && ~x2 && x3 && ~x19 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x18 && ~x2 && x3 && ~x19 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( x18 && ~x2 && x3 && ~x19 && ~x11 )
						nx_state = s1;
					else if( x18 && ~x2 && ~x3 && x19 && x4 && x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s820;
						end
					else if( x18 && ~x2 && ~x3 && x19 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s821;
						end
					else if( x18 && ~x2 && ~x3 && x19 && x4 && ~x5 && ~x6 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( x18 && ~x2 && ~x3 && x19 && ~x4 )
						begin
							y47 = 1'b1;	
							nx_state = s287;
						end
					else if( x18 && ~x2 && ~x3 && ~x19 && x4 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1612;
						end
					else if( x18 && ~x2 && ~x3 && ~x19 && ~x4 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s1321;
						end
					else if( ~x18 && x19 && x2 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1612;
						end
					else if( ~x18 && x19 && ~x2 && x4 && x3 )
						begin
							y23 = 1'b1;	y27 = 1'b1;	y48 = 1'b1;	
							nx_state = s1613;
						end
					else if( ~x18 && x19 && ~x2 && x4 && ~x3 )
						begin
							y37 = 1'b1;	
							nx_state = s888;
						end
					else if( ~x18 && x19 && ~x2 && ~x4 && x3 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s79;
						end
					else if( ~x18 && x19 && ~x2 && ~x4 && ~x3 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1093;
						end
					else if( ~x18 && ~x19 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1612;
						end
					else nx_state = s1499;
				s1500 : if( x14 )
						begin
							y1 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x14 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x14 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x14 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x14 && ~x11 )
						nx_state = s1;
					else nx_state = s1500;
				s1501 : if( 1'b1 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s1667;
						end
					else nx_state = s1501;
				s1502 : if( 1'b1 )
						begin
							y36 = 1'b1;	
							nx_state = s963;
						end
					else nx_state = s1502;
				s1503 : if( x64 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s1668;
						end
					else if( ~x64 )
						begin
							y40 = 1'b1;	
							nx_state = s1669;
						end
					else nx_state = s1503;
				s1504 : if( 1'b1 )
						begin
							y4 = 1'b1;	y31 = 1'b1;	y39 = 1'b1;	
							nx_state = s1240;
						end
					else nx_state = s1504;
				s1505 : if( 1'b1 )
						begin
							y9 = 1'b1;	
							nx_state = s1429;
						end
					else nx_state = s1505;
				s1506 : if( x62 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s561;
						end
					else if( ~x62 && x64 )
						begin
							y7 = 1'b1;	
							nx_state = s1272;
						end
					else if( ~x62 && ~x64 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s328;
						end
					else nx_state = s1506;
				s1507 : if( 1'b1 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else nx_state = s1507;
				s1508 : if( x64 )
						begin
							y3 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s1670;
						end
					else if( ~x64 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s1671;
						end
					else nx_state = s1508;
				s1509 : if( 1'b1 )
						begin
							y2 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							y53 = 1'b1;	
							nx_state = s1672;
						end
					else nx_state = s1509;
				s1510 : if( x7 && x9 && x8 && x3 && x2 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x7 && x9 && x8 && x3 && x2 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x7 && x9 && x8 && x3 && x2 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x7 && x9 && x8 && x3 && x2 && ~x1 )
						nx_state = s1;
					else if( x7 && x9 && x8 && x3 && ~x2 && x4 && x17 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x7 && x9 && x8 && x3 && ~x2 && x4 && ~x17 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x7 && x9 && x8 && x3 && ~x2 && x4 && ~x17 && x1 && ~x16 )
						nx_state = s1;
					else if( x7 && x9 && x8 && x3 && ~x2 && x4 && ~x17 && ~x1 )
						nx_state = s1;
					else if( x7 && x9 && x8 && x3 && ~x2 && ~x4 && x16 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( x7 && x9 && x8 && x3 && ~x2 && ~x4 && ~x16 && x1 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x7 && x9 && x8 && x3 && ~x2 && ~x4 && ~x16 && x1 && ~x17 )
						nx_state = s1;
					else if( x7 && x9 && x8 && x3 && ~x2 && ~x4 && ~x16 && ~x1 )
						nx_state = s1;
					else if( x7 && x9 && x8 && ~x3 && x4 && x2 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( x7 && x9 && x8 && ~x3 && x4 && ~x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	y29 = 1'b1;	
							nx_state = s673;
						end
					else if( x7 && x9 && x8 && ~x3 && ~x4 && x2 )
						begin
							y33 = 1'b1;	
							nx_state = s589;
						end
					else if( x7 && x9 && x8 && ~x3 && ~x4 && ~x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y29 = 1'b1;	
							y30 = 1'b1;	y31 = 1'b1;	
							nx_state = s1539;
						end
					else if( x7 && x9 && ~x8 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y13 = 1'b1;	y34 = 1'b1;	
							nx_state = s1673;
						end
					else if( x7 && ~x9 && x11 && x2 && x4 && x8 && x3 )
						begin
							y45 = 1'b1;	
							nx_state = s286;
						end
					else if( x7 && ~x9 && x11 && x2 && x4 && x8 && ~x3 )
						begin
							y46 = 1'b1;	
							nx_state = s531;
						end
					else if( x7 && ~x9 && x11 && x2 && x4 && ~x8 && x3 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x7 && ~x9 && x11 && x2 && x4 && ~x8 && ~x3 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x7 && ~x9 && x11 && x2 && ~x4 && x8 && x3 )
						begin
							y44 = 1'b1;	
							nx_state = s1138;
						end
					else if( x7 && ~x9 && x11 && x2 && ~x4 && x8 && ~x3 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x7 && ~x9 && x11 && x2 && ~x4 && ~x8 && x3 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x7 && ~x9 && x11 && x2 && ~x4 && ~x8 && ~x3 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x7 && ~x9 && x11 && ~x2 && x8 && x3 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x7 && ~x9 && x11 && ~x2 && x8 && x3 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x7 && ~x9 && x11 && ~x2 && x8 && x3 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x7 && ~x9 && x11 && ~x2 && x8 && x3 && ~x1 )
						nx_state = s1;
					else if( x7 && ~x9 && x11 && ~x2 && x8 && ~x3 && x4 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x7 && ~x9 && x11 && ~x2 && x8 && ~x3 && ~x4 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x7 && ~x9 && x11 && ~x2 && ~x8 && x4 && x3 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y38 = 1'b1;	
							y50 = 1'b1;	y51 = 1'b1;	
							nx_state = s1539;
						end
					else if( x7 && ~x9 && x11 && ~x2 && ~x8 && x4 && ~x3 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y38 = 1'b1;	
							y50 = 1'b1;	y51 = 1'b1;	
							nx_state = s1539;
						end
					else if( x7 && ~x9 && x11 && ~x2 && ~x8 && ~x4 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y38 = 1'b1;	
							y50 = 1'b1;	y51 = 1'b1;	
							nx_state = s1539;
						end
					else if( x7 && ~x9 && ~x11 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y13 = 1'b1;	y34 = 1'b1;	
							nx_state = s1673;
						end
					else if( ~x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s1674;
						end
					else nx_state = s1510;
				s1511 : if( x19 && x20 && x2 && x1 && x4 && x3 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x19 && x20 && x2 && x1 && x4 && x3 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x19 && x20 && x2 && x1 && x4 && x3 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( x19 && x20 && x2 && x1 && x4 && x3 && ~x22 )
						nx_state = s1;
					else if( x19 && x20 && x2 && x1 && x4 && ~x3 && x5 && x18 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x19 && x20 && x2 && x1 && x4 && ~x3 && x5 && ~x18 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x19 && x20 && x2 && x1 && x4 && ~x3 && x5 && ~x18 && x22 && ~x21 )
						nx_state = s1;
					else if( x19 && x20 && x2 && x1 && x4 && ~x3 && x5 && ~x18 && ~x22 )
						nx_state = s1;
					else if( x19 && x20 && x2 && x1 && x4 && ~x3 && ~x5 && x21 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x19 && x20 && x2 && x1 && x4 && ~x3 && ~x5 && ~x21 && x22 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x19 && x20 && x2 && x1 && x4 && ~x3 && ~x5 && ~x21 && x22 && ~x18 )
						nx_state = s1;
					else if( x19 && x20 && x2 && x1 && x4 && ~x3 && ~x5 && ~x21 && ~x22 )
						nx_state = s1;
					else if( x19 && x20 && x2 && x1 && ~x4 && x5 && x3 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x19 && x20 && x2 && x1 && ~x4 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y35 = 1'b1;	y36 = 1'b1;	
							nx_state = s654;
						end
					else if( x19 && x20 && x2 && x1 && ~x4 && ~x5 && x3 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x19 && x20 && x2 && x1 && ~x4 && ~x5 && ~x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y34 = 1'b1;	y37 = 1'b1;	
							nx_state = s654;
						end
					else if( x19 && x20 && x2 && ~x1 )
						begin
							y26 = 1'b1;	
							nx_state = s413;
						end
					else if( x19 && x20 && ~x2 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s715;
						end
					else if( x19 && x20 && ~x2 && ~x8 )
						begin
							y26 = 1'b1;	
							nx_state = s413;
						end
					else if( x19 && ~x20 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s716;
						end
					else if( ~x19 && x11 )
						begin
							y28 = 1'b1;	
							nx_state = s717;
						end
					else if( ~x19 && ~x11 )
						begin
							y29 = 1'b1;	
							nx_state = s771;
						end
					else nx_state = s1511;
				s1512 : if( x20 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s1485;
						end
					else if( ~x20 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s1656;
						end
					else nx_state = s1512;
				s1513 : if( 1'b1 )
						begin
							y40 = 1'b1;	
							nx_state = s1675;
						end
					else nx_state = s1513;
				s1514 : if( 1'b1 )
						begin
							y40 = 1'b1;	
							nx_state = s1676;
						end
					else nx_state = s1514;
				s1515 : if( 1'b1 )
						begin
							y38 = 1'b1;	
							nx_state = s845;
						end
					else nx_state = s1515;
				s1516 : if( 1'b1 )
						begin
							y54 = 1'b1;	
							nx_state = s281;
						end
					else nx_state = s1516;
				s1517 : if( x20 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x20 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x20 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x20 && x22 && ~x23 )
						nx_state = s1;
					else if( x20 && ~x22 )
						nx_state = s1;
					else if( ~x20 )
						begin
							y11 = 1'b1;	
							nx_state = s91;
						end
					else nx_state = s1517;
				s1518 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y59 = 1'b1;	
							y69 = 1'b1;	y70 = 1'b1;	y71 = 1'b1;	
							nx_state = s1677;
						end
					else nx_state = s1518;
				s1519 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y26 = 1'b1;	
							y63 = 1'b1;	
							nx_state = s741;
						end
					else nx_state = s1519;
				s1520 : if( x12 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x12 && x17 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x12 && x17 && ~x8 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x12 && x17 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x12 && ~x17 )
						nx_state = s1;
					else nx_state = s1520;
				s1521 : if( 1'b1 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s1678;
						end
					else nx_state = s1521;
				s1522 : if( 1'b1 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s1679;
						end
					else nx_state = s1522;
				s1523 : if( 1'b1 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y34 = 1'b1;	
							nx_state = s1680;
						end
					else nx_state = s1523;
				s1524 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y70 = 1'b1;	
							y71 = 1'b1;	y72 = 1'b1;	
							nx_state = s1681;
						end
					else nx_state = s1524;
				s1525 : if( 1'b1 )
						begin
							y4 = 1'b1;	y20 = 1'b1;	y27 = 1'b1;	
							nx_state = s1682;
						end
					else nx_state = s1525;
				s1526 : if( 1'b1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							nx_state = s1279;
						end
					else nx_state = s1526;
				s1527 : if( 1'b1 )
						begin
							y14 = 1'b1;	
							nx_state = s5;
						end
					else nx_state = s1527;
				s1528 : if( x62 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s683;
						end
					else if( x62 && ~x17 )
						begin
							y1 = 1'b1;	y12 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1353;
						end
					else if( ~x62 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else nx_state = s1528;
				s1529 : if( x6 && x19 && x18 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1683;
						end
					else if( x6 && x19 && ~x18 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s821;
						end
					else if( x6 && ~x19 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1683;
						end
					else if( ~x6 && x10 && x18 && x2 && x19 && x4 && x3 && x5 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1612;
						end
					else if( ~x6 && x10 && x18 && x2 && x19 && x4 && x3 && ~x5 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y21 = 1'b1;	
							y32 = 1'b1;	y35 = 1'b1;	
							nx_state = s1500;
						end
					else if( ~x6 && x10 && x18 && x2 && x19 && x4 && ~x3 && x17 && x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x6 && x10 && x18 && x2 && x19 && x4 && ~x3 && x17 && ~x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x6 && x10 && x18 && x2 && x19 && x4 && ~x3 && ~x17 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x6 && x10 && x18 && x2 && x19 && x4 && ~x3 && ~x17 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x6 && x10 && x18 && x2 && x19 && x4 && ~x3 && ~x17 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x6 && x10 && x18 && x2 && x19 && x4 && ~x3 && ~x17 && ~x11 )
						nx_state = s1;
					else if( ~x6 && x10 && x18 && x2 && x19 && ~x4 && x3 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y19 = 1'b1;	
							nx_state = s872;
						end
					else if( ~x6 && x10 && x18 && x2 && x19 && ~x4 && ~x3 && x16 && x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x6 && x10 && x18 && x2 && x19 && ~x4 && ~x3 && x16 && ~x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x6 && x10 && x18 && x2 && x19 && ~x4 && ~x3 && ~x16 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x6 && x10 && x18 && x2 && x19 && ~x4 && ~x3 && ~x16 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x6 && x10 && x18 && x2 && x19 && ~x4 && ~x3 && ~x16 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x6 && x10 && x18 && x2 && x19 && ~x4 && ~x3 && ~x16 && ~x11 )
						nx_state = s1;
					else if( ~x6 && x10 && x18 && x2 && ~x19 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x6 && x10 && x18 && x2 && ~x19 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x6 && x10 && x18 && x2 && ~x19 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x6 && x10 && x18 && x2 && ~x19 && ~x11 )
						nx_state = s1;
					else if( ~x6 && x10 && x18 && ~x2 && x3 && x19 && x4 && x15 && x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x6 && x10 && x18 && ~x2 && x3 && x19 && x4 && x15 && ~x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x6 && x10 && x18 && ~x2 && x3 && x19 && x4 && ~x15 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x6 && x10 && x18 && ~x2 && x3 && x19 && x4 && ~x15 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x6 && x10 && x18 && ~x2 && x3 && x19 && x4 && ~x15 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x6 && x10 && x18 && ~x2 && x3 && x19 && x4 && ~x15 && ~x11 )
						nx_state = s1;
					else if( ~x6 && x10 && x18 && ~x2 && x3 && x19 && ~x4 && x14 && x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x6 && x10 && x18 && ~x2 && x3 && x19 && ~x4 && x14 && ~x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x6 && x10 && x18 && ~x2 && x3 && x19 && ~x4 && ~x14 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x6 && x10 && x18 && ~x2 && x3 && x19 && ~x4 && ~x14 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x6 && x10 && x18 && ~x2 && x3 && x19 && ~x4 && ~x14 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x6 && x10 && x18 && ~x2 && x3 && x19 && ~x4 && ~x14 && ~x11 )
						nx_state = s1;
					else if( ~x6 && x10 && x18 && ~x2 && x3 && ~x19 && x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x6 && x10 && x18 && ~x2 && x3 && ~x19 && x11 && ~x12 && x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x6 && x10 && x18 && ~x2 && x3 && ~x19 && x11 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x6 && x10 && x18 && ~x2 && x3 && ~x19 && ~x11 )
						nx_state = s1;
					else if( ~x6 && x10 && x18 && ~x2 && ~x3 && x19 && x4 && x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x6 && x10 && x18 && ~x2 && ~x3 && x19 && x4 && ~x5 )
						begin
							y6 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x6 && x10 && x18 && ~x2 && ~x3 && x19 && ~x4 )
						begin
							y47 = 1'b1;	
							nx_state = s287;
						end
					else if( ~x6 && x10 && x18 && ~x2 && ~x3 && ~x19 && x4 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1612;
						end
					else if( ~x6 && x10 && x18 && ~x2 && ~x3 && ~x19 && ~x4 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s1321;
						end
					else if( ~x6 && x10 && ~x18 && x19 && x2 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1612;
						end
					else if( ~x6 && x10 && ~x18 && x19 && ~x2 && x4 && x3 )
						begin
							y23 = 1'b1;	y27 = 1'b1;	y48 = 1'b1;	
							nx_state = s1613;
						end
					else if( ~x6 && x10 && ~x18 && x19 && ~x2 && x4 && ~x3 )
						begin
							y37 = 1'b1;	
							nx_state = s888;
						end
					else if( ~x6 && x10 && ~x18 && x19 && ~x2 && ~x4 && x3 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s79;
						end
					else if( ~x6 && x10 && ~x18 && x19 && ~x2 && ~x4 && ~x3 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1093;
						end
					else if( ~x6 && x10 && ~x18 && ~x19 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1612;
						end
					else if( ~x6 && ~x10 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							y30 = 1'b1;	y35 = 1'b1;	y51 = 1'b1;	
							nx_state = s1499;
						end
					else nx_state = s1529;
				s1530 : if( 1'b1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y20 = 1'b1;	
							nx_state = s1287;
						end
					else nx_state = s1530;
				s1531 : if( x7 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s989;
						end
					else if( ~x7 && x19 && x23 && x4 && x5 && x3 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( ~x7 && x19 && x23 && x4 && x5 && x3 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( ~x7 && x19 && x23 && x4 && x5 && x3 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( ~x7 && x19 && x23 && x4 && x5 && x3 && ~x21 )
						nx_state = s1;
					else if( ~x7 && x19 && x23 && x4 && x5 && ~x3 && x12 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y23 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s535;
						end
					else if( ~x7 && x19 && x23 && x4 && x5 && ~x3 && ~x12 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( ~x7 && x19 && x23 && x4 && x5 && ~x3 && ~x12 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( ~x7 && x19 && x23 && x4 && x5 && ~x3 && ~x12 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( ~x7 && x19 && x23 && x4 && x5 && ~x3 && ~x12 && ~x21 )
						nx_state = s1;
					else if( ~x7 && x19 && x23 && x4 && ~x5 && x3 )
						begin
							y6 = 1'b1;	
							nx_state = s1506;
						end
					else if( ~x7 && x19 && x23 && x4 && ~x5 && ~x3 && x11 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y23 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s535;
						end
					else if( ~x7 && x19 && x23 && x4 && ~x5 && ~x3 && ~x11 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( ~x7 && x19 && x23 && x4 && ~x5 && ~x3 && ~x11 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( ~x7 && x19 && x23 && x4 && ~x5 && ~x3 && ~x11 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( ~x7 && x19 && x23 && x4 && ~x5 && ~x3 && ~x11 && ~x21 )
						nx_state = s1;
					else if( ~x7 && x19 && x23 && ~x4 && x3 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s1155;
						end
					else if( ~x7 && x19 && x23 && ~x4 && x3 && ~x5 && x13 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y23 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s535;
						end
					else if( ~x7 && x19 && x23 && ~x4 && x3 && ~x5 && ~x13 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( ~x7 && x19 && x23 && ~x4 && x3 && ~x5 && ~x13 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( ~x7 && x19 && x23 && ~x4 && x3 && ~x5 && ~x13 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( ~x7 && x19 && x23 && ~x4 && x3 && ~x5 && ~x13 && ~x21 )
						nx_state = s1;
					else if( ~x7 && x19 && x23 && ~x4 && ~x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y23 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s535;
						end
					else if( ~x7 && x19 && ~x23 && x22 && x4 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y9 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s1684;
						end
					else if( ~x7 && x19 && ~x23 && x22 && x4 && ~x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x7 && x19 && ~x23 && x22 && ~x4 )
						begin
							y6 = 1'b1;	
							nx_state = s368;
						end
					else if( ~x7 && x19 && ~x23 && ~x22 )
						begin
							y6 = 1'b1;	
							nx_state = s1506;
						end
					else if( ~x7 && ~x19 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y23 = 1'b1;	
							y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s1685;
						end
					else nx_state = s1531;
				s1532 : if( 1'b1 )
						begin
							y45 = 1'b1;	
							nx_state = s286;
						end
					else nx_state = s1532;
				s1533 : if( x6 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( ~x6 && x22 && x23 && x4 && x3 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( ~x6 && x22 && x23 && x4 && x3 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( ~x6 && x22 && x23 && x4 && x3 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( ~x6 && x22 && x23 && x4 && x3 && ~x21 )
						nx_state = s1;
					else if( ~x6 && x22 && x23 && x4 && ~x3 && x5 && x15 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x6 && x22 && x23 && x4 && ~x3 && x5 && ~x15 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( ~x6 && x22 && x23 && x4 && ~x3 && x5 && ~x15 && x21 && ~x16 )
						nx_state = s1;
					else if( ~x6 && x22 && x23 && x4 && ~x3 && x5 && ~x15 && ~x21 )
						nx_state = s1;
					else if( ~x6 && x22 && x23 && x4 && ~x3 && ~x5 && x16 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x6 && x22 && x23 && x4 && ~x3 && ~x5 && ~x16 && x21 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( ~x6 && x22 && x23 && x4 && ~x3 && ~x5 && ~x16 && x21 && ~x15 )
						nx_state = s1;
					else if( ~x6 && x22 && x23 && x4 && ~x3 && ~x5 && ~x16 && ~x21 )
						nx_state = s1;
					else if( ~x6 && x22 && x23 && ~x4 && x5 && x3 )
						begin
							y25 = 1'b1;	y26 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x6 && x22 && x23 && ~x4 && x5 && ~x3 )
						begin
							y1 = 1'b1;	y20 = 1'b1;	y47 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s535;
						end
					else if( ~x6 && x22 && x23 && ~x4 && ~x5 && x3 )
						begin
							y51 = 1'b1;	y52 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x6 && x22 && x23 && ~x4 && ~x5 && ~x3 )
						begin
							y1 = 1'b1;	y19 = 1'b1;	y49 = 1'b1;	
							y50 = 1'b1;	
							nx_state = s535;
						end
					else if( ~x6 && x22 && ~x23 && x9 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y36 = 1'b1;	
							nx_state = s535;
						end
					else if( ~x6 && x22 && ~x23 && ~x9 && x3 && x5 && x4 )
						begin
							y42 = 1'b1;	
							nx_state = s754;
						end
					else if( ~x6 && x22 && ~x23 && ~x9 && x3 && x5 && ~x4 )
						begin
							y40 = 1'b1;	
							nx_state = s751;
						end
					else if( ~x6 && x22 && ~x23 && ~x9 && x3 && ~x5 && x4 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x6 && x22 && ~x23 && ~x9 && x3 && ~x5 && ~x4 )
						begin
							y39 = 1'b1;	
							nx_state = s277;
						end
					else if( ~x6 && x22 && ~x23 && ~x9 && ~x3 && x7 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y8 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1685;
						end
					else if( ~x6 && x22 && ~x23 && ~x9 && ~x3 && ~x7 && x4 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s1686;
						end
					else if( ~x6 && x22 && ~x23 && ~x9 && ~x3 && ~x7 && x4 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s535;
						end
					else if( ~x6 && x22 && ~x23 && ~x9 && ~x3 && ~x7 && ~x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y27 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s535;
						end
					else if( ~x6 && ~x22 && x23 && x9 )
						begin
							y46 = 1'b1;	
							nx_state = s1030;
						end
					else if( ~x6 && ~x22 && x23 && ~x9 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y8 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1685;
						end
					else if( ~x6 && ~x22 && ~x23 && x3 && x5 && x4 )
						begin
							y31 = 1'b1;	y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s535;
						end
					else if( ~x6 && ~x22 && ~x23 && x3 && x5 && ~x4 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x6 && ~x22 && ~x23 && x3 && ~x5 && x4 )
						begin
							y30 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							nx_state = s535;
						end
					else if( ~x6 && ~x22 && ~x23 && x3 && ~x5 && ~x4 )
						begin
							y30 = 1'b1;	
							nx_state = s291;
						end
					else if( ~x6 && ~x22 && ~x23 && ~x3 && x7 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y8 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1685;
						end
					else if( ~x6 && ~x22 && ~x23 && ~x3 && ~x7 )
						begin
							y1 = 1'b1;	y27 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	y44 = 1'b1;	
							nx_state = s535;
						end
					else nx_state = s1533;
				s1534 : if( 1'b1 )
						begin
							y6 = 1'b1;	y39 = 1'b1;	y40 = 1'b1;	
							y41 = 1'b1;	y42 = 1'b1;	
							nx_state = s1687;
						end
					else nx_state = s1534;
				s1535 : if( 1'b1 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y27 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s749;
						end
					else nx_state = s1535;
				s1536 : if( 1'b1 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else nx_state = s1536;
				s1537 : if( x64 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1688;
						end
					else if( ~x64 )
						begin
							y48 = 1'b1;	y55 = 1'b1;	y61 = 1'b1;	
							nx_state = s1631;
						end
					else nx_state = s1537;
				s1538 : if( x7 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s1689;
						end
					else if( ~x7 && x9 && x6 && x12 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s1273;
						end
					else if( ~x7 && x9 && x6 && ~x12 && x11 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s1008;
						end
					else if( ~x7 && x9 && x6 && ~x12 && ~x11 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x7 && x9 && x6 && ~x12 && ~x11 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x7 && x9 && x6 && ~x12 && ~x11 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x7 && x9 && x6 && ~x12 && ~x11 && ~x18 )
						nx_state = s1;
					else if( ~x7 && x9 && ~x6 && x8 && x11 && x12 && x10 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x7 && x9 && ~x6 && x8 && x11 && x12 && x10 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x7 && x9 && ~x6 && x8 && x11 && x12 && x10 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x7 && x9 && ~x6 && x8 && x11 && x12 && x10 && ~x18 )
						nx_state = s1;
					else if( ~x7 && x9 && ~x6 && x8 && x11 && x12 && ~x10 && x16 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s749;
						end
					else if( ~x7 && x9 && ~x6 && x8 && x11 && x12 && ~x10 && ~x16 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x7 && x9 && ~x6 && x8 && x11 && x12 && ~x10 && ~x16 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x7 && x9 && ~x6 && x8 && x11 && x12 && ~x10 && ~x16 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x7 && x9 && ~x6 && x8 && x11 && x12 && ~x10 && ~x16 && ~x18 )
						nx_state = s1;
					else if( ~x7 && x9 && ~x6 && x8 && x11 && ~x12 && x10 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s1274;
						end
					else if( ~x7 && x9 && ~x6 && x8 && x11 && ~x12 && ~x10 && x17 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s749;
						end
					else if( ~x7 && x9 && ~x6 && x8 && x11 && ~x12 && ~x10 && ~x17 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x7 && x9 && ~x6 && x8 && x11 && ~x12 && ~x10 && ~x17 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x7 && x9 && ~x6 && x8 && x11 && ~x12 && ~x10 && ~x17 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x7 && x9 && ~x6 && x8 && x11 && ~x12 && ~x10 && ~x17 && ~x18 )
						nx_state = s1;
					else if( ~x7 && x9 && ~x6 && x8 && ~x11 && x12 && x10 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y34 = 1'b1;	
							nx_state = s1275;
						end
					else if( ~x7 && x9 && ~x6 && x8 && ~x11 && x12 && ~x10 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s749;
						end
					else if( ~x7 && x9 && ~x6 && x8 && ~x11 && ~x12 && x10 && x15 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s749;
						end
					else if( ~x7 && x9 && ~x6 && x8 && ~x11 && ~x12 && x10 && ~x15 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x7 && x9 && ~x6 && x8 && ~x11 && ~x12 && x10 && ~x15 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x7 && x9 && ~x6 && x8 && ~x11 && ~x12 && x10 && ~x15 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x7 && x9 && ~x6 && x8 && ~x11 && ~x12 && x10 && ~x15 && ~x18 )
						nx_state = s1;
					else if( ~x7 && x9 && ~x6 && x8 && ~x11 && ~x12 && ~x10 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x7 && x9 && ~x6 && ~x8 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s1273;
						end
					else if( ~x7 && ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y28 = 1'b1;	y33 = 1'b1;	
							nx_state = s750;
						end
					else nx_state = s1538;
				s1539 : if( x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x1 )
						nx_state = s1;
					else nx_state = s1539;
				s1540 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y38 = 1'b1;	
							nx_state = s1690;
						end
					else nx_state = s1540;
				s1541 : if( x16 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s427;
						end
					else if( ~x16 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y67 = 1'b1;	
							y68 = 1'b1;	
							nx_state = s1691;
						end
					else nx_state = s1541;
				s1542 : if( 1'b1 )
						begin
							y3 = 1'b1;	
							nx_state = s1569;
						end
					else nx_state = s1542;
				s1543 : if( x10 && x2 )
						nx_state = s1;
					else if( x10 && ~x2 && x3 && x4 && x5 && x1 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x10 && ~x2 && x3 && x4 && x5 && ~x1 )
						begin
							y41 = 1'b1;	y45 = 1'b1;	y46 = 1'b1;	
							nx_state = s654;
						end
					else if( x10 && ~x2 && x3 && x4 && ~x5 && x1 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( x10 && ~x2 && x3 && x4 && ~x5 && ~x1 )
						begin
							y39 = 1'b1;	y43 = 1'b1;	y44 = 1'b1;	
							nx_state = s654;
						end
					else if( x10 && ~x2 && x3 && ~x4 && x5 && x1 )
						begin
							y51 = 1'b1;	
							nx_state = s655;
						end
					else if( x10 && ~x2 && x3 && ~x4 && x5 && ~x1 )
						begin
							y41 = 1'b1;	y42 = 1'b1;	
							nx_state = s654;
						end
					else if( x10 && ~x2 && x3 && ~x4 && ~x5 && x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y48 = 1'b1;	
							y50 = 1'b1;	
							nx_state = s654;
						end
					else if( x10 && ~x2 && x3 && ~x4 && ~x5 && ~x1 )
						begin
							y39 = 1'b1;	y40 = 1'b1;	
							nx_state = s654;
						end
					else if( x10 && ~x2 && ~x3 && x4 && x5 && x1 && x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s651;
						end
					else if( x10 && ~x2 && ~x3 && x4 && x5 && x1 && ~x6 && x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s651;
						end
					else if( x10 && ~x2 && ~x3 && x4 && x5 && x1 && ~x6 && ~x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s652;
						end
					else if( x10 && ~x2 && ~x3 && x4 && x5 && ~x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y47 = 1'b1;	y48 = 1'b1;	
							nx_state = s654;
						end
					else if( x10 && ~x2 && ~x3 && x4 && ~x5 && x1 && x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s653;
						end
					else if( x10 && ~x2 && ~x3 && x4 && ~x5 && x1 && ~x6 && x7 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s653;
						end
					else if( x10 && ~x2 && ~x3 && x4 && ~x5 && x1 && ~x6 && ~x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s654;
						end
					else if( x10 && ~x2 && ~x3 && x4 && ~x5 && ~x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y48 = 1'b1;	y49 = 1'b1;	
							nx_state = s654;
						end
					else if( x10 && ~x2 && ~x3 && ~x4 && x1 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s654;
						end
					else if( x10 && ~x2 && ~x3 && ~x4 && x1 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s654;
						end
					else if( x10 && ~x2 && ~x3 && ~x4 && ~x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y32 = 1'b1;	y48 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x10 && x11 )
						begin
							y28 = 1'b1;	
							nx_state = s1326;
						end
					else if( ~x10 && ~x11 )
						begin
							y29 = 1'b1;	
							nx_state = s1661;
						end
					else nx_state = s1543;
				s1544 : if( x63 )
						begin
							y28 = 1'b1;	
							nx_state = s1565;
						end
					else if( ~x63 )
						begin
							y2 = 1'b1;	
							nx_state = s51;
						end
					else nx_state = s1544;
				s1545 : if( 1'b1 )
						begin
							y28 = 1'b1;	
							nx_state = s469;
						end
					else nx_state = s1545;
				s1546 : if( x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y23 = 1'b1;	y29 = 1'b1;	
							nx_state = s1092;
						end
					else if( ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1340;
						end
					else nx_state = s1546;
				s1547 : if( x7 && x13 && x8 && x9 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x7 && x13 && x8 && x9 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x7 && x13 && x8 && x9 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x7 && x13 && x8 && x9 && ~x14 )
						nx_state = s1;
					else if( x7 && x13 && x8 && ~x9 && x11 && x10 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x7 && x13 && x8 && ~x9 && x11 && x10 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x7 && x13 && x8 && ~x9 && x11 && x10 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x7 && x13 && x8 && ~x9 && x11 && x10 && ~x14 )
						nx_state = s1;
					else if( x7 && x13 && x8 && ~x9 && x11 && ~x10 )
						begin
							y2 = 1'b1;	
							nx_state = s768;
						end
					else if( x7 && x13 && x8 && ~x9 && ~x11 && x10 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y18 = 1'b1;	y20 = 1'b1;	
							nx_state = s1692;
						end
					else if( x7 && x13 && x8 && ~x9 && ~x11 && ~x10 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x7 && x13 && x8 && ~x9 && ~x11 && ~x10 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x7 && x13 && x8 && ~x9 && ~x11 && ~x10 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x7 && x13 && x8 && ~x9 && ~x11 && ~x10 && ~x14 )
						nx_state = s1;
					else if( x7 && x13 && ~x8 && x6 && x10 && x11 && x9 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x7 && x13 && ~x8 && x6 && x10 && x11 && x9 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x7 && x13 && ~x8 && x6 && x10 && x11 && x9 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x7 && x13 && ~x8 && x6 && x10 && x11 && x9 && ~x14 )
						nx_state = s1;
					else if( x7 && x13 && ~x8 && x6 && x10 && x11 && ~x9 && x18 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s1430;
						end
					else if( x7 && x13 && ~x8 && x6 && x10 && x11 && ~x9 && ~x18 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x7 && x13 && ~x8 && x6 && x10 && x11 && ~x9 && ~x18 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x7 && x13 && ~x8 && x6 && x10 && x11 && ~x9 && ~x18 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x7 && x13 && ~x8 && x6 && x10 && x11 && ~x9 && ~x18 && ~x14 )
						nx_state = s1;
					else if( x7 && x13 && ~x8 && x6 && x10 && ~x11 && x9 )
						begin
							y44 = 1'b1;	
							nx_state = s755;
						end
					else if( x7 && x13 && ~x8 && x6 && x10 && ~x11 && ~x9 && x17 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s1430;
						end
					else if( x7 && x13 && ~x8 && x6 && x10 && ~x11 && ~x9 && ~x17 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x7 && x13 && ~x8 && x6 && x10 && ~x11 && ~x9 && ~x17 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x7 && x13 && ~x8 && x6 && x10 && ~x11 && ~x9 && ~x17 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x7 && x13 && ~x8 && x6 && x10 && ~x11 && ~x9 && ~x17 && ~x14 )
						nx_state = s1;
					else if( x7 && x13 && ~x8 && x6 && ~x10 && x11 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s1693;
						end
					else if( x7 && x13 && ~x8 && x6 && ~x10 && x11 && ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s1430;
						end
					else if( x7 && x13 && ~x8 && x6 && ~x10 && ~x11 && x9 && x19 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s1430;
						end
					else if( x7 && x13 && ~x8 && x6 && ~x10 && ~x11 && x9 && ~x19 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x7 && x13 && ~x8 && x6 && ~x10 && ~x11 && x9 && ~x19 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x7 && x13 && ~x8 && x6 && ~x10 && ~x11 && x9 && ~x19 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x7 && x13 && ~x8 && x6 && ~x10 && ~x11 && x9 && ~x19 && ~x14 )
						nx_state = s1;
					else if( x7 && x13 && ~x8 && x6 && ~x10 && ~x11 && ~x9 )
						begin
							y44 = 1'b1;	
							nx_state = s1138;
						end
					else if( x7 && x13 && ~x8 && ~x6 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( x7 && ~x13 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y17 = 1'b1;	
							y27 = 1'b1;	y45 = 1'b1;	
							nx_state = s1694;
						end
					else if( ~x7 )
						begin
							y2 = 1'b1;	
							nx_state = s1695;
						end
					else nx_state = s1547;
				s1548 : if( x5 )
						begin
							y13 = 1'b1;	
							nx_state = s897;
						end
					else if( ~x5 && x6 && x8 && x9 && x12 )
						begin
							y47 = 1'b1;	
							nx_state = s287;
						end
					else if( ~x5 && x6 && x8 && x9 && ~x12 )
						begin
							y53 = 1'b1;	
							nx_state = s344;
						end
					else if( ~x5 && x6 && x8 && ~x9 && x10 && x11 && x16 )
						begin
							y48 = 1'b1;	
							nx_state = s676;
						end
					else if( ~x5 && x6 && x8 && ~x9 && x10 && x11 && ~x16 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x5 && x6 && x8 && ~x9 && x10 && x11 && ~x16 && x14 && ~x15 )
						nx_state = s1;
					else if( ~x5 && x6 && x8 && ~x9 && x10 && x11 && ~x16 && ~x14 )
						nx_state = s1;
					else if( ~x5 && x6 && x8 && ~x9 && x10 && ~x11 && x15 )
						begin
							y48 = 1'b1;	
							nx_state = s676;
						end
					else if( ~x5 && x6 && x8 && ~x9 && x10 && ~x11 && ~x15 && x14 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x5 && x6 && x8 && ~x9 && x10 && ~x11 && ~x15 && x14 && ~x16 )
						nx_state = s1;
					else if( ~x5 && x6 && x8 && ~x9 && x10 && ~x11 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x5 && x6 && x8 && ~x9 && ~x10 && x11 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y21 = 1'b1;	
							y51 = 1'b1;	y52 = 1'b1;	
							nx_state = s1430;
						end
					else if( ~x5 && x6 && x8 && ~x9 && ~x10 && ~x11 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y49 = 1'b1;	y50 = 1'b1;	
							nx_state = s1430;
						end
					else if( ~x5 && x6 && ~x8 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1694;
						end
					else if( ~x5 && ~x6 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1694;
						end
					else if( ~x5 && ~x6 && ~x7 && x9 && x10 && x11 && x8 )
						begin
							y25 = 1'b1;	
							nx_state = s1605;
						end
					else if( ~x5 && ~x6 && ~x7 && x9 && x10 && x11 && ~x8 )
						begin
							y32 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							nx_state = s1430;
						end
					else if( ~x5 && ~x6 && ~x7 && x9 && x10 && ~x11 && x8 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x5 && ~x6 && ~x7 && x9 && x10 && ~x11 && ~x8 )
						begin
							y30 = 1'b1;	y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s1430;
						end
					else if( ~x5 && ~x6 && ~x7 && x9 && ~x10 && x11 && x8 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( ~x5 && ~x6 && ~x7 && x9 && ~x10 && x11 && ~x8 )
						begin
							y32 = 1'b1;	y33 = 1'b1;	
							nx_state = s396;
						end
					else if( ~x5 && ~x6 && ~x7 && x9 && ~x10 && ~x11 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x5 && ~x6 && ~x7 && x9 && ~x10 && ~x11 && ~x8 )
						begin
							y30 = 1'b1;	y31 = 1'b1;	
							nx_state = s1022;
						end
					else if( ~x5 && ~x6 && ~x7 && ~x9 && x10 && x11 && x8 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y17 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s389;
						end
					else if( ~x5 && ~x6 && ~x7 && ~x9 && x10 && x11 && ~x8 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							y26 = 1'b1;	y29 = 1'b1;	
							nx_state = s1430;
						end
					else if( ~x5 && ~x6 && ~x7 && ~x9 && x10 && ~x11 && x8 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s1430;
						end
					else if( ~x5 && ~x6 && ~x7 && ~x9 && x10 && ~x11 && ~x8 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							y26 = 1'b1;	y28 = 1'b1;	
							nx_state = s1430;
						end
					else if( ~x5 && ~x6 && ~x7 && ~x9 && ~x10 && x8 && x11 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1430;
						end
					else if( ~x5 && ~x6 && ~x7 && ~x9 && ~x10 && x8 && ~x11 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							nx_state = s1430;
						end
					else if( ~x5 && ~x6 && ~x7 && ~x9 && ~x10 && ~x8 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s1430;
						end
					else nx_state = s1548;
				s1549 : if( 1'b1 )
						begin
							y47 = 1'b1;	y56 = 1'b1;	y61 = 1'b1;	
							y70 = 1'b1;	
							nx_state = s1463;
						end
					else nx_state = s1549;
				s1550 : if( x5 && x9 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1696;
						end
					else if( x5 && x9 && ~x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y13 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1697;
						end
					else if( x5 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y26 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s1417;
						end
					else if( ~x5 && x6 && x17 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x5 && x6 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x5 && ~x6 )
						begin
							y5 = 1'b1;	y26 = 1'b1;	y29 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s1417;
						end
					else nx_state = s1550;
				s1551 : if( x9 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1698;
						end
					else if( ~x9 && x15 && x11 && x6 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( ~x9 && x15 && x11 && x6 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x9 && x15 && x11 && ~x6 && x7 && x10 )
						begin
							y48 = 1'b1;	
							nx_state = s1009;
						end
					else if( ~x9 && x15 && x11 && ~x6 && x7 && ~x10 && x12 && x18 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y47 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x9 && x15 && x11 && ~x6 && x7 && ~x10 && x12 && ~x18 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( ~x9 && x15 && x11 && ~x6 && x7 && ~x10 && x12 && ~x18 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( ~x9 && x15 && x11 && ~x6 && x7 && ~x10 && x12 && ~x18 && x19 && ~x14 && ~x13 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( ~x9 && x15 && x11 && ~x6 && x7 && ~x10 && x12 && ~x18 && ~x19 )
						nx_state = s1;
					else if( ~x9 && x15 && x11 && ~x6 && x7 && ~x10 && ~x12 && x17 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y47 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x9 && x15 && x11 && ~x6 && x7 && ~x10 && ~x12 && ~x17 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( ~x9 && x15 && x11 && ~x6 && x7 && ~x10 && ~x12 && ~x17 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( ~x9 && x15 && x11 && ~x6 && x7 && ~x10 && ~x12 && ~x17 && x19 && ~x14 && ~x13 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x9 && x15 && x11 && ~x6 && x7 && ~x10 && ~x12 && ~x17 && ~x19 )
						nx_state = s1;
					else if( ~x9 && x15 && x11 && ~x6 && ~x7 && x12 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	y38 = 1'b1;	y40 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x9 && x15 && x11 && ~x6 && ~x7 && ~x12 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	y38 = 1'b1;	y41 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x9 && x15 && ~x11 && x6 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x9 && x15 && ~x11 && ~x6 && x7 && x12 && x10 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y45 = 1'b1;	
							y49 = 1'b1;	
							nx_state = s1576;
						end
					else if( ~x9 && x15 && ~x11 && ~x6 && x7 && x12 && ~x10 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y47 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x9 && x15 && ~x11 && ~x6 && x7 && ~x12 && x10 && x16 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y47 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x9 && x15 && ~x11 && ~x6 && x7 && ~x12 && x10 && ~x16 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( ~x9 && x15 && ~x11 && ~x6 && x7 && ~x12 && x10 && ~x16 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( ~x9 && x15 && ~x11 && ~x6 && x7 && ~x12 && x10 && ~x16 && x19 && ~x14 && ~x13 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x9 && x15 && ~x11 && ~x6 && x7 && ~x12 && x10 && ~x16 && ~x19 )
						nx_state = s1;
					else if( ~x9 && x15 && ~x11 && ~x6 && x7 && ~x12 && ~x10 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x9 && x15 && ~x11 && ~x6 && ~x7 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	y38 = 1'b1;	y42 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x9 && ~x15 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y33 = 1'b1;	
							y40 = 1'b1;	y47 = 1'b1;	
							nx_state = s1699;
						end
					else nx_state = s1551;
				s1552 : if( 1'b1 )
						begin
							y8 = 1'b1;	y31 = 1'b1;	
							nx_state = s345;
						end
					else nx_state = s1552;
				s1553 : if( 1'b1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s1307;
						end
					else nx_state = s1553;
				s1554 : if( 1'b1 )
						begin
							y38 = 1'b1;	
							nx_state = s1700;
						end
					else nx_state = s1554;
				s1555 : if( 1'b1 )
						begin
							y3 = 1'b1;	y19 = 1'b1;	y44 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1701;
						end
					else nx_state = s1555;
				s1556 : if( x6 && x5 )
						nx_state = s1;
					else if( x6 && ~x5 && x7 && x8 )
						begin
							y46 = 1'b1;	
							nx_state = s1428;
						end
					else if( x6 && ~x5 && x7 && ~x8 && x9 )
						begin
							y3 = 1'b1;	y19 = 1'b1;	y42 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s1555;
						end
					else if( x6 && ~x5 && x7 && ~x8 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( x6 && ~x5 && ~x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( ~x6 )
						begin
							y46 = 1'b1;	
							nx_state = s1428;
						end
					else nx_state = s1556;
				s1557 : if( x6 && x5 )
						nx_state = s1;
					else if( x6 && ~x5 )
						begin
							y69 = 1'b1;	
							nx_state = s1123;
						end
					else if( ~x6 && x8 && x9 && x5 )
						begin
							y51 = 1'b1;	
							nx_state = s391;
						end
					else if( ~x6 && x8 && x9 && ~x5 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y62 = 1'b1;	
							y63 = 1'b1;	y65 = 1'b1;	y66 = 1'b1;	
							nx_state = s1314;
						end
					else if( ~x6 && x8 && x9 && ~x5 && ~x7 )
						begin
							y5 = 1'b1;	y27 = 1'b1;	y57 = 1'b1;	
							y58 = 1'b1;	
							nx_state = s1314;
						end
					else if( ~x6 && x8 && ~x9 && x5 )
						begin
							y3 = 1'b1;	y19 = 1'b1;	y53 = 1'b1;	
							nx_state = s1314;
						end
					else if( ~x6 && x8 && ~x9 && ~x5 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y59 = 1'b1;	
							y60 = 1'b1;	y67 = 1'b1;	y68 = 1'b1;	
							nx_state = s1314;
						end
					else if( ~x6 && x8 && ~x9 && ~x5 && ~x7 )
						begin
							y5 = 1'b1;	y27 = 1'b1;	y55 = 1'b1;	
							y56 = 1'b1;	
							nx_state = s1314;
						end
					else if( ~x6 && ~x8 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1314;
						end
					else if( ~x6 && ~x8 && ~x5 && x7 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y62 = 1'b1;	
							y63 = 1'b1;	y64 = 1'b1;	
							nx_state = s1314;
						end
					else if( ~x6 && ~x8 && ~x5 && x7 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y59 = 1'b1;	
							y60 = 1'b1;	y61 = 1'b1;	
							nx_state = s1314;
						end
					else if( ~x6 && ~x8 && ~x5 && ~x7 )
						begin
							y5 = 1'b1;	y27 = 1'b1;	y41 = 1'b1;	
							y54 = 1'b1;	
							nx_state = s1314;
						end
					else nx_state = s1557;
				s1558 : if( 1'b1 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else nx_state = s1558;
				s1559 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y24 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1702;
						end
					else nx_state = s1559;
				s1560 : if( x63 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x63 )
						begin
							y10 = 1'b1;	y22 = 1'b1;	y23 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s1560;
				s1561 : if( 1'b1 )
						begin
							y2 = 1'b1;	y15 = 1'b1;	y31 = 1'b1;	
							nx_state = s1703;
						end
					else nx_state = s1561;
				s1562 : if( x6 && x8 && x27 && x7 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s1220;
						end
					else if( x6 && x8 && x27 && ~x7 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1220;
						end
					else if( x6 && x8 && ~x27 && x7 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( x6 && x8 && ~x27 && ~x7 )
						begin
							y40 = 1'b1;	
							nx_state = s751;
						end
					else if( x6 && ~x8 && x27 && x7 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y47 = 1'b1;	
							nx_state = s1220;
						end
					else if( x6 && ~x8 && x27 && ~x7 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y46 = 1'b1;	
							nx_state = s1220;
						end
					else if( x6 && ~x8 && ~x27 && x7 )
						begin
							y39 = 1'b1;	
							nx_state = s277;
						end
					else if( x6 && ~x8 && ~x27 && ~x7 )
						begin
							y18 = 1'b1;	y41 = 1'b1;	y42 = 1'b1;	
							nx_state = s1221;
						end
					else if( ~x6 && x7 && x27 && x8 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y42 = 1'b1;	y44 = 1'b1;	
							nx_state = s1220;
						end
					else if( ~x6 && x7 && x27 && ~x8 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y42 = 1'b1;	y44 = 1'b1;	
							nx_state = s1220;
						end
					else if( ~x6 && x7 && ~x27 && x13 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x6 && x7 && ~x27 && x13 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x6 && x7 && ~x27 && x13 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x6 && x7 && ~x27 && x13 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x6 && x7 && ~x27 && x13 && ~x22 )
						nx_state = s1;
					else if( ~x6 && x7 && ~x27 && ~x13 && x3 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x6 && x7 && ~x27 && ~x13 && x3 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x6 && x7 && ~x27 && ~x13 && x3 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x6 && x7 && ~x27 && ~x13 && x3 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x6 && x7 && ~x27 && ~x13 && x3 && ~x22 )
						nx_state = s1;
					else if( ~x6 && x7 && ~x27 && ~x13 && ~x3 )
						begin
							y5 = 1'b1;	y34 = 1'b1;	y41 = 1'b1;	
							y42 = 1'b1;	
							nx_state = s1222;
						end
					else if( ~x6 && ~x7 && x27 )
						begin
							y5 = 1'b1;	y32 = 1'b1;	y41 = 1'b1;	
							y42 = 1'b1;	y44 = 1'b1;	
							nx_state = s1220;
						end
					else if( ~x6 && ~x7 && ~x27 && x8 )
						begin
							y5 = 1'b1;	y17 = 1'b1;	y32 = 1'b1;	
							y42 = 1'b1;	
							nx_state = s1220;
						end
					else if( ~x6 && ~x7 && ~x27 && ~x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y32 = 1'b1;	
							nx_state = s1220;
						end
					else nx_state = s1562;
				s1563 : if( 1'b1 )
						begin
							y7 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s1563;
				s1564 : if( x9 && x1 && x3 )
						begin
							y26 = 1'b1;	
							nx_state = s1197;
						end
					else if( x9 && x1 && ~x3 && x4 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s656;
						end
					else if( x9 && x1 && ~x3 && x4 && ~x5 && x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s653;
						end
					else if( x9 && x1 && ~x3 && x4 && ~x5 && ~x6 && x7 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s653;
						end
					else if( x9 && x1 && ~x3 && x4 && ~x5 && ~x6 && ~x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s654;
						end
					else if( x9 && x1 && ~x3 && ~x4 )
						begin
							y26 = 1'b1;	
							nx_state = s1197;
						end
					else if( x9 && ~x1 && x2 && x4 && x3 )
						begin
							y26 = 1'b1;	
							nx_state = s1468;
						end
					else if( x9 && ~x1 && x2 && x4 && ~x3 && x5 && x15 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s654;
						end
					else if( x9 && ~x1 && x2 && x4 && ~x3 && x5 && ~x15 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x9 && ~x1 && x2 && x4 && ~x3 && x5 && ~x15 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x9 && ~x1 && x2 && x4 && ~x3 && x5 && ~x15 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( x9 && ~x1 && x2 && x4 && ~x3 && x5 && ~x15 && ~x22 )
						nx_state = s1;
					else if( x9 && ~x1 && x2 && x4 && ~x3 && ~x5 && x17 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s654;
						end
					else if( x9 && ~x1 && x2 && x4 && ~x3 && ~x5 && ~x17 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x9 && ~x1 && x2 && x4 && ~x3 && ~x5 && ~x17 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x9 && ~x1 && x2 && x4 && ~x3 && ~x5 && ~x17 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( x9 && ~x1 && x2 && x4 && ~x3 && ~x5 && ~x17 && ~x22 )
						nx_state = s1;
					else if( x9 && ~x1 && x2 && ~x4 && x5 && x3 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1509;
						end
					else if( x9 && ~x1 && x2 && ~x4 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s654;
						end
					else if( x9 && ~x1 && x2 && ~x4 && ~x5 && x3 && x16 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s654;
						end
					else if( x9 && ~x1 && x2 && ~x4 && ~x5 && x3 && ~x16 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x9 && ~x1 && x2 && ~x4 && ~x5 && x3 && ~x16 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x9 && ~x1 && x2 && ~x4 && ~x5 && x3 && ~x16 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( x9 && ~x1 && x2 && ~x4 && ~x5 && x3 && ~x16 && ~x22 )
						nx_state = s1;
					else if( x9 && ~x1 && x2 && ~x4 && ~x5 && ~x3 )
						begin
							y38 = 1'b1;	
							nx_state = s845;
						end
					else if( x9 && ~x1 && ~x2 )
						begin
							y26 = 1'b1;	
							nx_state = s1197;
						end
					else if( ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y8 = 1'b1;	y32 = 1'b1;	
							nx_state = s1610;
						end
					else nx_state = s1564;
				s1565 : if( x65 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y14 = 1'b1;	
							y15 = 1'b1;	y21 = 1'b1;	
							nx_state = s1704;
						end
					else if( ~x65 )
						begin
							y15 = 1'b1;	
							nx_state = s356;
						end
					else nx_state = s1565;
				s1566 : if( x10 && x2 && x3 && x4 && x9 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x10 && x2 && x3 && x4 && x9 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x10 && x2 && x3 && x4 && x9 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x10 && x2 && x3 && x4 && x9 && ~x1 )
						nx_state = s1;
					else if( x10 && x2 && x3 && x4 && ~x9 && x8 )
						begin
							y45 = 1'b1;	
							nx_state = s286;
						end
					else if( x10 && x2 && x3 && x4 && ~x9 && ~x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x10 && x2 && x3 && ~x4 && x9 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s602;
						end
					else if( x10 && x2 && x3 && ~x4 && x9 && ~x6 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x10 && x2 && x3 && ~x4 && ~x9 && x8 )
						begin
							y44 = 1'b1;	
							nx_state = s1138;
						end
					else if( x10 && x2 && x3 && ~x4 && ~x9 && ~x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x10 && x2 && ~x3 && x4 && x9 )
						begin
							y3 = 1'b1;	y18 = 1'b1;	y21 = 1'b1;	
							nx_state = s1382;
						end
					else if( x10 && x2 && ~x3 && x4 && ~x9 && x8 )
						begin
							y46 = 1'b1;	
							nx_state = s531;
						end
					else if( x10 && x2 && ~x3 && x4 && ~x9 && ~x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x10 && x2 && ~x3 && ~x4 && x9 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( x10 && x2 && ~x3 && ~x4 && x9 && ~x13 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x10 && x2 && ~x3 && ~x4 && x9 && ~x13 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x10 && x2 && ~x3 && ~x4 && x9 && ~x13 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x10 && x2 && ~x3 && ~x4 && x9 && ~x13 && ~x1 )
						nx_state = s1;
					else if( x10 && x2 && ~x3 && ~x4 && ~x9 && x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x10 && x2 && ~x3 && ~x4 && ~x9 && ~x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x10 && ~x2 && x4 && x3 && x9 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( x10 && ~x2 && x4 && x3 && x9 && ~x14 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x10 && ~x2 && x4 && x3 && x9 && ~x14 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x10 && ~x2 && x4 && x3 && x9 && ~x14 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x10 && ~x2 && x4 && x3 && x9 && ~x14 && ~x1 )
						nx_state = s1;
					else if( x10 && ~x2 && x4 && x3 && ~x9 && x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y37 = 1'b1;	
							nx_state = s1540;
						end
					else if( x10 && ~x2 && x4 && x3 && ~x9 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x10 && ~x2 && x4 && ~x3 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( x10 && ~x2 && x4 && ~x3 && ~x9 && x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x10 && ~x2 && x4 && ~x3 && ~x9 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x10 && ~x2 && ~x4 && x9 && x3 && x12 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( x10 && ~x2 && ~x4 && x9 && x3 && ~x12 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x10 && ~x2 && ~x4 && x9 && x3 && ~x12 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x10 && ~x2 && ~x4 && x9 && x3 && ~x12 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x10 && ~x2 && ~x4 && x9 && x3 && ~x12 && ~x1 )
						nx_state = s1;
					else if( x10 && ~x2 && ~x4 && x9 && ~x3 )
						begin
							y26 = 1'b1;	
							nx_state = s1197;
						end
					else if( x10 && ~x2 && ~x4 && ~x9 && x8 && x3 )
						begin
							y3 = 1'b1;	y18 = 1'b1;	y42 = 1'b1;	
							nx_state = s1539;
						end
					else if( x10 && ~x2 && ~x4 && ~x9 && x8 && ~x3 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x10 && ~x2 && ~x4 && ~x9 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y36 = 1'b1;	y40 = 1'b1;	
							nx_state = s1705;
						end
					else nx_state = s1566;
				s1567 : if( x21 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x21 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x21 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x21 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 )
						begin
							y56 = 1'b1;	
							nx_state = s1007;
						end
					else if( ~x21 && ~x22 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && ~x22 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && ~x22 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x6 )
						nx_state = s1;
					else nx_state = s1567;
				s1568 : if( x21 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x21 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( x21 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( x21 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && x20 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x21 && x22 && ~x20 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && ~x20 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && x22 && ~x20 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x20 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && ~x22 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x21 && ~x22 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x6 )
						nx_state = s1;
					else nx_state = s1568;
				s1569 : if( x63 )
						begin
							y21 = 1'b1;	y28 = 1'b1;	y48 = 1'b1;	
							nx_state = s839;
						end
					else if( ~x63 )
						begin
							y47 = 1'b1;	y52 = 1'b1;	y61 = 1'b1;	
							y66 = 1'b1;	
							nx_state = s54;
						end
					else nx_state = s1569;
				s1570 : if( 1'b1 )
						begin
							y33 = 1'b1;	
							nx_state = s589;
						end
					else nx_state = s1570;
				s1571 : if( x16 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x16 && ~x12 && x13 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x16 && ~x12 && ~x13 )
						nx_state = s1;
					else if( ~x16 )
						nx_state = s1;
					else nx_state = s1571;
				s1572 : if( 1'b1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s1619;
						end
					else nx_state = s1572;
				s1573 : if( 1'b1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s1617;
						end
					else nx_state = s1573;
				s1574 : if( 1'b1 )
						begin
							y3 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	y30 = 1'b1;	
							nx_state = s1618;
						end
					else nx_state = s1574;
				s1575 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1571;
						end
					else nx_state = s1575;
				s1576 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y55 = 1'b1;	
							y58 = 1'b1;	y69 = 1'b1;	
							nx_state = s1706;
						end
					else nx_state = s1576;
				s1577 : if( x18 && x8 && x7 )
						begin
							y5 = 1'b1;	y19 = 1'b1;	y25 = 1'b1;	
							y27 = 1'b1;	y30 = 1'b1;	
							nx_state = s1578;
						end
					else if( x18 && x8 && ~x7 && x9 && x14 )
						begin
							y61 = 1'b1;	
							nx_state = s1098;
						end
					else if( x18 && x8 && ~x7 && x9 && ~x14 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x18 && x8 && ~x7 && x9 && ~x14 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x18 && x8 && ~x7 && x9 && ~x14 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x18 && x8 && ~x7 && x9 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x18 && x8 && ~x7 && ~x9 && x12 )
						begin
							y61 = 1'b1;	
							nx_state = s1098;
						end
					else if( x18 && x8 && ~x7 && ~x9 && ~x12 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x18 && x8 && ~x7 && ~x9 && ~x12 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x18 && x8 && ~x7 && ~x9 && ~x12 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x18 && x8 && ~x7 && ~x9 && ~x12 && ~x15 )
						nx_state = s1;
					else if( x18 && ~x8 && x9 && x7 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y26 = 1'b1;	
							nx_state = s1579;
						end
					else if( x18 && ~x8 && x9 && ~x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s1580;
						end
					else if( x18 && ~x8 && ~x9 && x7 && x13 )
						begin
							y61 = 1'b1;	
							nx_state = s1098;
						end
					else if( x18 && ~x8 && ~x9 && x7 && ~x13 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x18 && ~x8 && ~x9 && x7 && ~x13 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x18 && ~x8 && ~x9 && x7 && ~x13 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x18 && ~x8 && ~x9 && x7 && ~x13 && ~x15 )
						nx_state = s1;
					else if( x18 && ~x8 && ~x9 && ~x7 )
						begin
							y69 = 1'b1;	
							nx_state = s1123;
						end
					else if( ~x18 )
						begin
							y5 = 1'b1;	y19 = 1'b1;	y23 = 1'b1;	
							y25 = 1'b1;	y27 = 1'b1;	
							nx_state = s1581;
						end
					else nx_state = s1577;
				s1578 : if( 1'b1 )
						begin
							y5 = 1'b1;	y19 = 1'b1;	y25 = 1'b1;	
							y27 = 1'b1;	y30 = 1'b1;	
							nx_state = s1707;
						end
					else nx_state = s1578;
				s1579 : if( 1'b1 )
						begin
							y5 = 1'b1;	y19 = 1'b1;	y25 = 1'b1;	
							y27 = 1'b1;	y30 = 1'b1;	
							nx_state = s1708;
						end
					else nx_state = s1579;
				s1580 : if( x65 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x65 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x65 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x15 )
						nx_state = s1;
					else if( ~x65 && x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && x26 && ~x25 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && x26 && ~x25 && ~x24 )
						nx_state = s1;
					else if( ~x65 && ~x26 )
						nx_state = s1;
					else nx_state = s1580;
				s1581 : if( x8 && x7 )
						begin
							y5 = 1'b1;	y19 = 1'b1;	y25 = 1'b1;	
							y27 = 1'b1;	y30 = 1'b1;	
							nx_state = s1578;
						end
					else if( x8 && ~x7 && x9 && x14 )
						begin
							y61 = 1'b1;	
							nx_state = s1098;
						end
					else if( x8 && ~x7 && x9 && ~x14 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x8 && ~x7 && x9 && ~x14 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x8 && ~x7 && x9 && ~x14 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x8 && ~x7 && x9 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x8 && ~x7 && ~x9 && x12 )
						begin
							y61 = 1'b1;	
							nx_state = s1098;
						end
					else if( x8 && ~x7 && ~x9 && ~x12 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x8 && ~x7 && ~x9 && ~x12 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x8 && ~x7 && ~x9 && ~x12 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x8 && ~x7 && ~x9 && ~x12 && ~x15 )
						nx_state = s1;
					else if( ~x8 && x9 && x7 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y26 = 1'b1;	
							nx_state = s1579;
						end
					else if( ~x8 && x9 && ~x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s1580;
						end
					else if( ~x8 && ~x9 && x7 && x13 )
						begin
							y61 = 1'b1;	
							nx_state = s1098;
						end
					else if( ~x8 && ~x9 && x7 && ~x13 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x8 && ~x9 && x7 && ~x13 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x8 && ~x9 && x7 && ~x13 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x8 && ~x9 && x7 && ~x13 && ~x15 )
						nx_state = s1;
					else if( ~x8 && ~x9 && ~x7 )
						begin
							y69 = 1'b1;	
							nx_state = s1123;
						end
					else nx_state = s1581;
				s1582 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y22 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s1400;
						end
					else nx_state = s1582;
				s1583 : if( x65 && x18 && x8 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s1584;
						end
					else if( x65 && x18 && x8 && ~x9 )
						begin
							y3 = 1'b1;	y26 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1400;
						end
					else if( x65 && x18 && ~x8 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1400;
						end
					else if( x65 && ~x18 )
						begin
							y5 = 1'b1;	y19 = 1'b1;	y23 = 1'b1;	
							y25 = 1'b1;	y27 = 1'b1;	
							nx_state = s1585;
						end
					else if( ~x65 )
						begin
							y9 = 1'b1;	
							nx_state = s1709;
						end
					else nx_state = s1583;
				s1584 : if( 1'b1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1400;
						end
					else nx_state = s1584;
				s1585 : if( x8 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s1584;
						end
					else if( x8 && ~x9 )
						begin
							y3 = 1'b1;	y26 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1400;
						end
					else if( ~x8 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1400;
						end
					else nx_state = s1585;
				s1586 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y52 = 1'b1;	
							y55 = 1'b1;	
							nx_state = s1400;
						end
					else nx_state = s1586;
				s1587 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y41 = 1'b1;	
							y55 = 1'b1;	
							nx_state = s1400;
						end
					else nx_state = s1587;
				s1588 : if( x18 && x8 && x9 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y55 = 1'b1;	y65 = 1'b1;	
							nx_state = s1589;
						end
					else if( x18 && x8 && x9 && ~x7 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1400;
						end
					else if( x18 && x8 && ~x9 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y47 = 1'b1;	y49 = 1'b1;	
							nx_state = s1590;
						end
					else if( x18 && x8 && ~x9 && ~x7 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							y20 = 1'b1;	y22 = 1'b1;	
							nx_state = s1400;
						end
					else if( x18 && ~x8 && x7 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y66 = 1'b1;	
							y67 = 1'b1;	
							nx_state = s1591;
						end
					else if( x18 && ~x8 && x7 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y56 = 1'b1;	
							y57 = 1'b1;	
							nx_state = s1592;
						end
					else if( x18 && ~x8 && ~x7 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	y22 = 1'b1;	
							nx_state = s1400;
						end
					else if( ~x18 )
						begin
							y5 = 1'b1;	y19 = 1'b1;	y23 = 1'b1;	
							y25 = 1'b1;	y27 = 1'b1;	
							nx_state = s1593;
						end
					else nx_state = s1588;
				s1589 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y66 = 1'b1;	
							y67 = 1'b1;	
							nx_state = s1710;
						end
					else nx_state = s1589;
				s1590 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y56 = 1'b1;	
							y57 = 1'b1;	
							nx_state = s1711;
						end
					else nx_state = s1590;
				s1591 : if( 1'b1 )
						begin
							y3 = 1'b1;	y26 = 1'b1;	y63 = 1'b1;	
							nx_state = s1400;
						end
					else nx_state = s1591;
				s1592 : if( 1'b1 )
						begin
							y3 = 1'b1;	y26 = 1'b1;	y62 = 1'b1;	
							nx_state = s1400;
						end
					else nx_state = s1592;
				s1593 : if( x8 && x9 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y55 = 1'b1;	y65 = 1'b1;	
							nx_state = s1589;
						end
					else if( x8 && x9 && ~x7 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1400;
						end
					else if( x8 && ~x9 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y47 = 1'b1;	y49 = 1'b1;	
							nx_state = s1590;
						end
					else if( x8 && ~x9 && ~x7 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							y20 = 1'b1;	y22 = 1'b1;	
							nx_state = s1400;
						end
					else if( ~x8 && x7 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y66 = 1'b1;	
							y67 = 1'b1;	
							nx_state = s1591;
						end
					else if( ~x8 && x7 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y56 = 1'b1;	
							y57 = 1'b1;	
							nx_state = s1592;
						end
					else if( ~x8 && ~x7 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							y19 = 1'b1;	y22 = 1'b1;	
							nx_state = s1400;
						end
					else nx_state = s1593;
				s1594 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y22 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s1712;
						end
					else nx_state = s1594;
				s1595 : if( x63 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x63 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x63 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x63 && ~x1 )
						nx_state = s1;
					else if( ~x63 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x63 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x63 && ~x15 )
						nx_state = s1;
					else nx_state = s1595;
				s1596 : if( 1'b1 )
						begin
							y5 = 1'b1;	y19 = 1'b1;	y30 = 1'b1;	
							y39 = 1'b1;	y60 = 1'b1;	
							nx_state = s1713;
						end
					else nx_state = s1596;
				s1597 : if( 1'b1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y26 = 1'b1;	
							nx_state = s1714;
						end
					else nx_state = s1597;
				s1598 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s1580;
						end
					else nx_state = s1598;
				s1599 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y44 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1715;
						end
					else nx_state = s1599;
				s1600 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y42 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s1716;
						end
					else nx_state = s1600;
				s1601 : if( x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1269;
						end
					else if( ~x15 && x17 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x15 && ~x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else nx_state = s1601;
				s1602 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y25 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s1717;
						end
					else nx_state = s1602;
				s1603 : if( x3 && x12 && x11 && x14 && x15 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y24 = 1'b1;	
							y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s1078;
						end
					else if( x3 && x12 && x11 && x14 && x15 && ~x13 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( x3 && x12 && x11 && x14 && ~x15 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	y34 = 1'b1;	
							nx_state = s1078;
						end
					else if( x3 && x12 && x11 && x14 && ~x15 && ~x13 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( x3 && x12 && x11 && ~x14 && x13 && x15 && x9 )
						begin
							y11 = 1'b1;	
							nx_state = s91;
						end
					else if( x3 && x12 && x11 && ~x14 && x13 && x15 && ~x9 && x8 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x3 && x12 && x11 && ~x14 && x13 && x15 && ~x9 && x8 && ~x10 )
						nx_state = s1;
					else if( x3 && x12 && x11 && ~x14 && x13 && x15 && ~x9 && ~x8 )
						nx_state = s1;
					else if( x3 && x12 && x11 && ~x14 && x13 && ~x15 && x10 )
						begin
							y11 = 1'b1;	
							nx_state = s91;
						end
					else if( x3 && x12 && x11 && ~x14 && x13 && ~x15 && ~x10 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x3 && x12 && x11 && ~x14 && x13 && ~x15 && ~x10 && x8 && ~x9 )
						nx_state = s1;
					else if( x3 && x12 && x11 && ~x14 && x13 && ~x15 && ~x10 && ~x8 )
						nx_state = s1;
					else if( x3 && x12 && x11 && ~x14 && ~x13 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x3 && x12 && x11 && ~x14 && ~x13 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x3 && x12 && x11 && ~x14 && ~x13 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x3 && x12 && x11 && ~x14 && ~x13 && ~x8 )
						nx_state = s1;
					else if( x3 && x12 && ~x11 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1718;
						end
					else if( x3 && ~x12 && x6 && x11 && x13 && x15 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y42 = 1'b1;	
							nx_state = s1078;
						end
					else if( x3 && ~x12 && x6 && x11 && x13 && x15 && ~x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y42 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s1078;
						end
					else if( x3 && ~x12 && x6 && x11 && x13 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y21 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s1078;
						end
					else if( x3 && ~x12 && x6 && x11 && x13 && ~x15 && ~x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1719;
						end
					else if( x3 && ~x12 && x6 && x11 && ~x13 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x3 && ~x12 && x6 && x11 && ~x13 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x3 && ~x12 && x6 && x11 && ~x13 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x3 && ~x12 && x6 && x11 && ~x13 && ~x8 )
						nx_state = s1;
					else if( x3 && ~x12 && x6 && ~x11 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1720;
						end
					else if( x3 && ~x12 && ~x6 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1718;
						end
					else if( ~x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1721;
						end
					else nx_state = s1603;
				s1604 : if( x5 && x7 && x9 && x8 )
						begin
							y47 = 1'b1;	
							nx_state = s675;
						end
					else if( x5 && x7 && x9 && ~x8 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( x5 && x7 && ~x9 && x8 )
						begin
							y48 = 1'b1;	
							nx_state = s676;
						end
					else if( x5 && x7 && ~x9 && ~x8 )
						begin
							y50 = 1'b1;	
							nx_state = s658;
						end
					else if( x5 && ~x7 && x8 && x9 && x3 )
						begin
							y51 = 1'b1;	
							nx_state = s655;
						end
					else if( x5 && ~x7 && x8 && x9 && ~x3 && x10 )
						begin
							y51 = 1'b1;	
							nx_state = s655;
						end
					else if( x5 && ~x7 && x8 && x9 && ~x3 && ~x10 )
						begin
							y51 = 1'b1;	
							nx_state = s391;
						end
					else if( x5 && ~x7 && x8 && ~x9 && x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s677;
						end
					else if( x5 && ~x7 && x8 && ~x9 && ~x3 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s677;
						end
					else if( x5 && ~x7 && x8 && ~x9 && ~x3 && ~x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y53 = 1'b1;	
							nx_state = s672;
						end
					else if( x5 && ~x7 && ~x8 && x3 && x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y55 = 1'b1;	
							nx_state = s672;
						end
					else if( x5 && ~x7 && ~x8 && x3 && ~x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s672;
						end
					else if( x5 && ~x7 && ~x8 && ~x3 && x9 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s672;
						end
					else if( x5 && ~x7 && ~x8 && ~x3 && x9 && ~x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							y54 = 1'b1;	
							nx_state = s672;
						end
					else if( x5 && ~x7 && ~x8 && ~x3 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s672;
						end
					else if( ~x5 && x8 && x9 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	y66 = 1'b1;	
							nx_state = s672;
						end
					else if( ~x5 && x8 && ~x9 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	y66 = 1'b1;	
							nx_state = s672;
						end
					else if( ~x5 && ~x8 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y66 = 1'b1;	
							nx_state = s672;
						end
					else nx_state = s1604;
				s1605 : if( x64 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x64 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x64 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x64 && ~x14 )
						nx_state = s1;
					else if( ~x64 && x14 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x64 && x14 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x64 && x14 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x64 && x14 && ~x23 )
						nx_state = s1;
					else if( ~x64 && ~x14 )
						begin
							y47 = 1'b1;	y56 = 1'b1;	y61 = 1'b1;	
							y72 = 1'b1;	
							nx_state = s1187;
						end
					else nx_state = s1605;
				s1606 : if( 1'b1 )
						begin
							y2 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1722;
						end
					else nx_state = s1606;
				s1607 : if( 1'b1 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s237;
						end
					else nx_state = s1607;
				s1608 : if( 1'b1 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y54 = 1'b1;	
							nx_state = s1723;
						end
					else nx_state = s1608;
				s1609 : if( 1'b1 )
						begin
							y9 = 1'b1;	
							nx_state = s1724;
						end
					else nx_state = s1609;
				s1610 : if( x1 && x3 )
						begin
							y26 = 1'b1;	
							nx_state = s1197;
						end
					else if( x1 && ~x3 && x4 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s656;
						end
					else if( x1 && ~x3 && x4 && ~x5 && x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s653;
						end
					else if( x1 && ~x3 && x4 && ~x5 && ~x6 && x7 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s653;
						end
					else if( x1 && ~x3 && x4 && ~x5 && ~x6 && ~x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s654;
						end
					else if( x1 && ~x3 && ~x4 )
						begin
							y26 = 1'b1;	
							nx_state = s1197;
						end
					else if( ~x1 && x2 && x4 && x3 )
						begin
							y26 = 1'b1;	
							nx_state = s1468;
						end
					else if( ~x1 && x2 && x4 && ~x3 && x5 && x15 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x1 && x2 && x4 && ~x3 && x5 && ~x15 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x1 && x2 && x4 && ~x3 && x5 && ~x15 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x1 && x2 && x4 && ~x3 && x5 && ~x15 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( ~x1 && x2 && x4 && ~x3 && x5 && ~x15 && ~x22 )
						nx_state = s1;
					else if( ~x1 && x2 && x4 && ~x3 && ~x5 && x17 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x1 && x2 && x4 && ~x3 && ~x5 && ~x17 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x1 && x2 && x4 && ~x3 && ~x5 && ~x17 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x1 && x2 && x4 && ~x3 && ~x5 && ~x17 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( ~x1 && x2 && x4 && ~x3 && ~x5 && ~x17 && ~x22 )
						nx_state = s1;
					else if( ~x1 && x2 && ~x4 && x5 && x3 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1509;
						end
					else if( ~x1 && x2 && ~x4 && x5 && ~x3 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x1 && x2 && ~x4 && ~x5 && x3 && x16 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x1 && x2 && ~x4 && ~x5 && x3 && ~x16 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x1 && x2 && ~x4 && ~x5 && x3 && ~x16 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x1 && x2 && ~x4 && ~x5 && x3 && ~x16 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( ~x1 && x2 && ~x4 && ~x5 && x3 && ~x16 && ~x22 )
						nx_state = s1;
					else if( ~x1 && x2 && ~x4 && ~x5 && ~x3 )
						begin
							y38 = 1'b1;	
							nx_state = s845;
						end
					else if( ~x1 && ~x2 )
						begin
							y26 = 1'b1;	
							nx_state = s1197;
						end
					else nx_state = s1610;
				s1611 : if( x21 && x26 && x27 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x21 && x26 && x27 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x21 && x26 && x27 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x21 && x26 && x27 && x22 && ~x23 )
						nx_state = s1;
					else if( x21 && x26 && x27 && ~x22 )
						nx_state = s1;
					else if( x21 && x26 && ~x27 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1627;
						end
					else if( x21 && ~x26 && x7 && x8 && x6 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x21 && ~x26 && x7 && x8 && x6 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x21 && ~x26 && x7 && x8 && x6 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x21 && ~x26 && x7 && x8 && x6 && x22 && ~x23 )
						nx_state = s1;
					else if( x21 && ~x26 && x7 && x8 && x6 && ~x22 )
						nx_state = s1;
					else if( x21 && ~x26 && x7 && x8 && ~x6 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( x21 && ~x26 && x7 && x8 && ~x6 && ~x9 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x21 && ~x26 && x7 && x8 && ~x6 && ~x9 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x21 && ~x26 && x7 && x8 && ~x6 && ~x9 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x21 && ~x26 && x7 && x8 && ~x6 && ~x9 && x22 && ~x23 )
						nx_state = s1;
					else if( x21 && ~x26 && x7 && x8 && ~x6 && ~x9 && ~x22 )
						nx_state = s1;
					else if( x21 && ~x26 && x7 && ~x8 && x6 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( x21 && ~x26 && x7 && ~x8 && ~x6 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( x21 && ~x26 && x7 && ~x8 && ~x6 && ~x10 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x21 && ~x26 && x7 && ~x8 && ~x6 && ~x10 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x21 && ~x26 && x7 && ~x8 && ~x6 && ~x10 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x21 && ~x26 && x7 && ~x8 && ~x6 && ~x10 && x22 && ~x23 )
						nx_state = s1;
					else if( x21 && ~x26 && x7 && ~x8 && ~x6 && ~x10 && ~x22 )
						nx_state = s1;
					else if( x21 && ~x26 && ~x7 && x8 && x6 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y42 = 1'b1;	
							nx_state = s1628;
						end
					else if( x21 && ~x26 && ~x7 && x8 && ~x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( x21 && ~x26 && ~x7 && ~x8 && x6 && x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( x21 && ~x26 && ~x7 && ~x8 && x6 && ~x11 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x21 && ~x26 && ~x7 && ~x8 && x6 && ~x11 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x21 && ~x26 && ~x7 && ~x8 && x6 && ~x11 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x21 && ~x26 && ~x7 && ~x8 && x6 && ~x11 && x22 && ~x23 )
						nx_state = s1;
					else if( x21 && ~x26 && ~x7 && ~x8 && x6 && ~x11 && ~x22 )
						nx_state = s1;
					else if( x21 && ~x26 && ~x7 && ~x8 && ~x6 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else if( ~x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y28 = 1'b1;	y29 = 1'b1;	
							nx_state = s1629;
						end
					else nx_state = s1611;
				s1612 : if( x19 && x18 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( x19 && ~x18 )
						begin
							y23 = 1'b1;	y27 = 1'b1;	y48 = 1'b1;	
							nx_state = s1725;
						end
					else if( ~x19 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else nx_state = s1612;
				s1613 : if( 1'b1 )
						begin
							y2 = 1'b1;	
							nx_state = s1726;
						end
					else nx_state = s1613;
				s1614 : if( 1'b1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y5 = 1'b1;	
							y22 = 1'b1;	y23 = 1'b1;	
							nx_state = s1541;
						end
					else nx_state = s1614;
				s1615 : if( x18 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1727;
						end
					else if( ~x18 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s1615;
						end
					else nx_state = s1615;
				s1616 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y19 = 1'b1;	
							nx_state = s1728;
						end
					else nx_state = s1616;
				s1617 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s1729;
						end
					else nx_state = s1617;
				s1618 : if( 1'b1 )
						begin
							y3 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	y32 = 1'b1;	
							nx_state = s1575;
						end
					else nx_state = s1618;
				s1619 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y19 = 1'b1;	
							nx_state = s1730;
						end
					else nx_state = s1619;
				s1620 : if( x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s1616;
						end
					else if( ~x4 && x5 && x6 && x7 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s1617;
						end
					else if( ~x4 && x5 && x6 && ~x7 )
						begin
							y3 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	y30 = 1'b1;	
							nx_state = s1618;
						end
					else if( ~x4 && x5 && ~x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1571;
						end
					else if( ~x4 && ~x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s1619;
						end
					else nx_state = s1620;
				s1621 : if( 1'b1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							nx_state = s1103;
						end
					else nx_state = s1621;
				s1622 : if( x19 && x23 && x4 && x5 && x3 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x19 && x23 && x4 && x5 && x3 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x19 && x23 && x4 && x5 && x3 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( x19 && x23 && x4 && x5 && x3 && ~x21 )
						nx_state = s1;
					else if( x19 && x23 && x4 && x5 && ~x3 && x12 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y23 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s535;
						end
					else if( x19 && x23 && x4 && x5 && ~x3 && ~x12 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x19 && x23 && x4 && x5 && ~x3 && ~x12 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x19 && x23 && x4 && x5 && ~x3 && ~x12 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( x19 && x23 && x4 && x5 && ~x3 && ~x12 && ~x21 )
						nx_state = s1;
					else if( x19 && x23 && x4 && ~x5 && x3 )
						begin
							y6 = 1'b1;	
							nx_state = s1506;
						end
					else if( x19 && x23 && x4 && ~x5 && ~x3 && x11 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y23 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s535;
						end
					else if( x19 && x23 && x4 && ~x5 && ~x3 && ~x11 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x19 && x23 && x4 && ~x5 && ~x3 && ~x11 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x19 && x23 && x4 && ~x5 && ~x3 && ~x11 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( x19 && x23 && x4 && ~x5 && ~x3 && ~x11 && ~x21 )
						nx_state = s1;
					else if( x19 && x23 && ~x4 && x3 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s1155;
						end
					else if( x19 && x23 && ~x4 && x3 && ~x5 && x13 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y23 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s535;
						end
					else if( x19 && x23 && ~x4 && x3 && ~x5 && ~x13 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x19 && x23 && ~x4 && x3 && ~x5 && ~x13 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x19 && x23 && ~x4 && x3 && ~x5 && ~x13 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( x19 && x23 && ~x4 && x3 && ~x5 && ~x13 && ~x21 )
						nx_state = s1;
					else if( x19 && x23 && ~x4 && ~x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y23 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s535;
						end
					else if( x19 && ~x23 && x22 && x4 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y9 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s1684;
						end
					else if( x19 && ~x23 && x22 && x4 && ~x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( x19 && ~x23 && x22 && ~x4 )
						begin
							y6 = 1'b1;	
							nx_state = s368;
						end
					else if( x19 && ~x23 && ~x22 )
						begin
							y6 = 1'b1;	
							nx_state = s1506;
						end
					else if( ~x19 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y23 = 1'b1;	
							y27 = 1'b1;	y28 = 1'b1;	
							nx_state = s1685;
						end
					else nx_state = s1622;
				s1623 : if( x14 && x21 && x9 )
						begin
							y44 = 1'b1;	
							nx_state = s755;
						end
					else if( x14 && x21 && ~x9 )
						begin
							y44 = 1'b1;	
							nx_state = s1138;
						end
					else if( x14 && ~x21 && x5 && x8 && x7 )
						begin
							y44 = 1'b1;	
							nx_state = s755;
						end
					else if( x14 && ~x21 && x5 && x8 && ~x7 && x9 && x18 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1263;
						end
					else if( x14 && ~x21 && x5 && x8 && ~x7 && x9 && ~x18 && x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x14 && ~x21 && x5 && x8 && ~x7 && x9 && ~x18 && x10 && ~x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x14 && ~x21 && x5 && x8 && ~x7 && x9 && ~x18 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x14 && ~x21 && x5 && x8 && ~x7 && x9 && ~x18 && ~x10 )
						nx_state = s1;
					else if( x14 && ~x21 && x5 && x8 && ~x7 && ~x9 && x19 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1263;
						end
					else if( x14 && ~x21 && x5 && x8 && ~x7 && ~x9 && ~x19 && x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x14 && ~x21 && x5 && x8 && ~x7 && ~x9 && ~x19 && x10 && ~x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x14 && ~x21 && x5 && x8 && ~x7 && ~x9 && ~x19 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x14 && ~x21 && x5 && x8 && ~x7 && ~x9 && ~x19 && ~x10 )
						nx_state = s1;
					else if( x14 && ~x21 && x5 && ~x8 && x7 && x9 )
						begin
							y2 = 1'b1;	
							nx_state = s437;
						end
					else if( x14 && ~x21 && x5 && ~x8 && x7 && ~x9 && x20 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1263;
						end
					else if( x14 && ~x21 && x5 && ~x8 && x7 && ~x9 && ~x20 && x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x14 && ~x21 && x5 && ~x8 && x7 && ~x9 && ~x20 && x10 && ~x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x14 && ~x21 && x5 && ~x8 && x7 && ~x9 && ~x20 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( x14 && ~x21 && x5 && ~x8 && x7 && ~x9 && ~x20 && ~x10 )
						nx_state = s1;
					else if( x14 && ~x21 && x5 && ~x8 && ~x7 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s1263;
						end
					else if( x14 && ~x21 && ~x5 )
						begin
							y44 = 1'b1;	
							nx_state = s755;
						end
					else if( ~x14 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y21 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s1264;
						end
					else nx_state = s1623;
				s1624 : if( 1'b1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y8 = 1'b1;	y10 = 1'b1;	y26 = 1'b1;	
							nx_state = s1444;
						end
					else nx_state = s1624;
				s1625 : if( x64 && x20 )
						begin
							y7 = 1'b1;	y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s467;
						end
					else if( x64 && ~x20 )
						begin
							y14 = 1'b1;	
							nx_state = s366;
						end
					else if( ~x64 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	
							nx_state = s328;
						end
					else nx_state = s1625;
				s1626 : if( 1'b1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s371;
						end
					else nx_state = s1626;
				s1627 : if( x63 )
						begin
							y9 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x63 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else nx_state = s1627;
				s1628 : if( 1'b1 )
						begin
							y11 = 1'b1;	
							nx_state = s271;
						end
					else nx_state = s1628;
				s1629 : if( x26 && x27 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x26 && x27 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( x26 && x27 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( x26 && x27 && x22 && ~x23 )
						nx_state = s1;
					else if( x26 && x27 && ~x22 )
						nx_state = s1;
					else if( x26 && ~x27 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1627;
						end
					else if( ~x26 && x7 && x8 && x6 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x26 && x7 && x8 && x6 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x26 && x7 && x8 && x6 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x26 && x7 && x8 && x6 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x26 && x7 && x8 && x6 && ~x22 )
						nx_state = s1;
					else if( ~x26 && x7 && x8 && ~x6 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( ~x26 && x7 && x8 && ~x6 && ~x9 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x26 && x7 && x8 && ~x6 && ~x9 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x26 && x7 && x8 && ~x6 && ~x9 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x26 && x7 && x8 && ~x6 && ~x9 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x26 && x7 && x8 && ~x6 && ~x9 && ~x22 )
						nx_state = s1;
					else if( ~x26 && x7 && ~x8 && x6 )
						begin
							y11 = 1'b1;	
							nx_state = s241;
						end
					else if( ~x26 && x7 && ~x8 && ~x6 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( ~x26 && x7 && ~x8 && ~x6 && ~x10 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x26 && x7 && ~x8 && ~x6 && ~x10 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x26 && x7 && ~x8 && ~x6 && ~x10 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x26 && x7 && ~x8 && ~x6 && ~x10 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x26 && x7 && ~x8 && ~x6 && ~x10 && ~x22 )
						nx_state = s1;
					else if( ~x26 && ~x7 && x8 && x6 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	y42 = 1'b1;	
							nx_state = s1628;
						end
					else if( ~x26 && ~x7 && x8 && ~x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( ~x26 && ~x7 && ~x8 && x6 && x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( ~x26 && ~x7 && ~x8 && x6 && ~x11 && x22 && x23 && x24 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x26 && ~x7 && ~x8 && x6 && ~x11 && x22 && x23 && ~x24 && x25 )
						begin
							y59 = 1'b1;	
							nx_state = s417;
						end
					else if( ~x26 && ~x7 && ~x8 && x6 && ~x11 && x22 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x26 && ~x7 && ~x8 && x6 && ~x11 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x26 && ~x7 && ~x8 && x6 && ~x11 && ~x22 )
						nx_state = s1;
					else if( ~x26 && ~x7 && ~x8 && ~x6 )
						begin
							y49 = 1'b1;	
							nx_state = s528;
						end
					else nx_state = s1629;
				s1630 : if( 1'b1 )
						begin
							y25 = 1'b1;	
							nx_state = s1731;
						end
					else nx_state = s1630;
				s1631 : if( 1'b1 )
						begin
							y25 = 1'b1;	
							nx_state = s53;
						end
					else nx_state = s1631;
				s1632 : if( 1'b1 )
						begin
							y10 = 1'b1;	y25 = 1'b1;	y26 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s1632;
				s1633 : if( 1'b1 )
						begin
							y74 = 1'b1;	
							nx_state = s1732;
						end
					else nx_state = s1633;
				s1634 : if( x14 && x7 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1635;
						end
					else if( x14 && ~x7 && x5 && x10 && x9 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1636;
						end
					else if( x14 && ~x7 && x5 && x10 && ~x9 && x11 && x16 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1455;
						end
					else if( x14 && ~x7 && x5 && x10 && ~x9 && x11 && ~x16 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x14 && ~x7 && x5 && x10 && ~x9 && x11 && ~x16 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x14 && ~x7 && x5 && x10 && ~x9 && x11 && ~x16 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x14 && ~x7 && x5 && x10 && ~x9 && x11 && ~x16 && ~x19 )
						nx_state = s1;
					else if( x14 && ~x7 && x5 && x10 && ~x9 && ~x11 && x17 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1455;
						end
					else if( x14 && ~x7 && x5 && x10 && ~x9 && ~x11 && ~x17 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x14 && ~x7 && x5 && x10 && ~x9 && ~x11 && ~x17 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x14 && ~x7 && x5 && x10 && ~x9 && ~x11 && ~x17 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x14 && ~x7 && x5 && x10 && ~x9 && ~x11 && ~x17 && ~x19 )
						nx_state = s1;
					else if( x14 && ~x7 && x5 && ~x10 && x11 && x9 )
						begin
							y6 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s80;
						end
					else if( x14 && ~x7 && x5 && ~x10 && x11 && ~x9 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1455;
						end
					else if( x14 && ~x7 && x5 && ~x10 && ~x11 && x9 && x15 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1455;
						end
					else if( x14 && ~x7 && x5 && ~x10 && ~x11 && x9 && ~x15 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x14 && ~x7 && x5 && ~x10 && ~x11 && x9 && ~x15 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x14 && ~x7 && x5 && ~x10 && ~x11 && x9 && ~x15 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x14 && ~x7 && x5 && ~x10 && ~x11 && x9 && ~x15 && ~x19 )
						nx_state = s1;
					else if( x14 && ~x7 && x5 && ~x10 && ~x11 && ~x9 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( x14 && ~x7 && ~x5 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1637;
						end
					else if( ~x14 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	y18 = 1'b1;	
							nx_state = s1638;
						end
					else nx_state = s1634;
				s1635 : if( 1'b1 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y43 = 1'b1;	
							y44 = 1'b1;	y45 = 1'b1;	
							nx_state = s1733;
						end
					else nx_state = s1635;
				s1636 : if( 1'b1 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y43 = 1'b1;	
							y44 = 1'b1;	y45 = 1'b1;	
							nx_state = s1734;
						end
					else nx_state = s1636;
				s1637 : if( 1'b1 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y43 = 1'b1;	
							y44 = 1'b1;	y45 = 1'b1;	
							nx_state = s1735;
						end
					else nx_state = s1637;
				s1638 : if( x7 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1635;
						end
					else if( ~x7 && x5 && x10 && x9 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1636;
						end
					else if( ~x7 && x5 && x10 && ~x9 && x11 && x16 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1455;
						end
					else if( ~x7 && x5 && x10 && ~x9 && x11 && ~x16 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x7 && x5 && x10 && ~x9 && x11 && ~x16 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x7 && x5 && x10 && ~x9 && x11 && ~x16 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x7 && x5 && x10 && ~x9 && x11 && ~x16 && ~x19 )
						nx_state = s1;
					else if( ~x7 && x5 && x10 && ~x9 && ~x11 && x17 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1455;
						end
					else if( ~x7 && x5 && x10 && ~x9 && ~x11 && ~x17 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x7 && x5 && x10 && ~x9 && ~x11 && ~x17 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x7 && x5 && x10 && ~x9 && ~x11 && ~x17 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x7 && x5 && x10 && ~x9 && ~x11 && ~x17 && ~x19 )
						nx_state = s1;
					else if( ~x7 && x5 && ~x10 && x11 && x9 )
						begin
							y6 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s80;
						end
					else if( ~x7 && x5 && ~x10 && x11 && ~x9 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1455;
						end
					else if( ~x7 && x5 && ~x10 && ~x11 && x9 && x15 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y15 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1455;
						end
					else if( ~x7 && x5 && ~x10 && ~x11 && x9 && ~x15 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x7 && x5 && ~x10 && ~x11 && x9 && ~x15 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x7 && x5 && ~x10 && ~x11 && x9 && ~x15 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x7 && x5 && ~x10 && ~x11 && x9 && ~x15 && ~x19 )
						nx_state = s1;
					else if( ~x7 && x5 && ~x10 && ~x11 && ~x9 )
						begin
							y24 = 1'b1;	
							nx_state = s257;
						end
					else if( ~x7 && ~x5 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1637;
						end
					else nx_state = s1638;
				s1639 : if( 1'b1 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y46 = 1'b1;	
							y47 = 1'b1;	
							nx_state = s1736;
						end
					else nx_state = s1639;
				s1640 : if( 1'b1 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y52 = 1'b1;	
							y53 = 1'b1;	
							nx_state = s1737;
						end
					else nx_state = s1640;
				s1641 : if( x62 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x62 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x62 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x62 && ~x19 )
						nx_state = s1;
					else if( ~x62 && x14 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x62 && x14 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x62 && x14 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x62 && x14 && ~x23 )
						nx_state = s1;
					else if( ~x62 && ~x14 )
						begin
							y47 = 1'b1;	y57 = 1'b1;	y61 = 1'b1;	
							y71 = 1'b1;	
							nx_state = s1271;
						end
					else nx_state = s1641;
				s1642 : if( 1'b1 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y48 = 1'b1;	
							nx_state = s1455;
						end
					else nx_state = s1642;
				s1643 : if( 1'b1 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y54 = 1'b1;	
							nx_state = s1455;
						end
					else nx_state = s1643;
				s1644 : if( 1'b1 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1738;
						end
					else nx_state = s1644;
				s1645 : if( 1'b1 )
						begin
							y7 = 1'b1;	y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s467;
						end
					else nx_state = s1645;
				s1646 : if( 1'b1 )
						begin
							y1 = 1'b1;	y37 = 1'b1;	y39 = 1'b1;	
							nx_state = s584;
						end
					else nx_state = s1646;
				s1647 : if( 1'b1 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else nx_state = s1647;
				s1648 : if( x17 )
						begin
							y24 = 1'b1;	
							nx_state = s590;
						end
					else if( ~x17 )
						begin
							y5 = 1'b1;	y13 = 1'b1;	y17 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1648;
						end
					else nx_state = s1648;
				s1649 : if( 1'b1 )
						begin
							y25 = 1'b1;	
							nx_state = s1641;
						end
					else nx_state = s1649;
				s1650 : if( 1'b1 )
						begin
							y6 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s1739;
						end
					else nx_state = s1650;
				s1651 : if( x5 && x21 && x7 && x9 )
						begin
							y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x5 && x21 && x7 && ~x9 )
						begin
							y50 = 1'b1;	
							nx_state = s658;
						end
					else if( x5 && x21 && ~x7 && x8 && x9 && x12 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x5 && x21 && ~x7 && x8 && x9 && ~x12 && x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x5 && x21 && ~x7 && x8 && x9 && ~x12 && x10 && ~x11 )
						nx_state = s1;
					else if( x5 && x21 && ~x7 && x8 && x9 && ~x12 && ~x10 )
						nx_state = s1;
					else if( x5 && x21 && ~x7 && x8 && ~x9 && x11 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x5 && x21 && ~x7 && x8 && ~x9 && ~x11 && x10 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( x5 && x21 && ~x7 && x8 && ~x9 && ~x11 && x10 && ~x12 )
						nx_state = s1;
					else if( x5 && x21 && ~x7 && x8 && ~x9 && ~x11 && ~x10 )
						nx_state = s1;
					else if( x5 && x21 && ~x7 && ~x8 && x9 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							y39 = 1'b1;	y40 = 1'b1;	
							nx_state = s1263;
						end
					else if( x5 && x21 && ~x7 && ~x8 && ~x9 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y16 = 1'b1;	
							y42 = 1'b1;	y51 = 1'b1;	
							nx_state = s1263;
						end
					else if( x5 && ~x21 && x16 )
						begin
							y34 = 1'b1;	
							nx_state = s103;
						end
					else if( x5 && ~x21 && ~x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1264;
						end
					else if( ~x5 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1264;
						end
					else if( ~x5 && ~x6 && x8 && x9 && x21 && x7 )
						begin
							y36 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x5 && ~x6 && x8 && x9 && x21 && ~x7 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1740;
						end
					else if( ~x5 && ~x6 && x8 && x9 && ~x21 && x7 )
						begin
							y6 = 1'b1;	y30 = 1'b1;	y31 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s1263;
						end
					else if( ~x5 && ~x6 && x8 && x9 && ~x21 && ~x7 )
						begin
							y6 = 1'b1;	y29 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	y32 = 1'b1;	
							nx_state = s1263;
						end
					else if( ~x5 && ~x6 && x8 && ~x9 && x21 && x7 )
						begin
							y37 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x5 && ~x6 && x8 && ~x9 && x21 && ~x7 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y31 = 1'b1;	
							y47 = 1'b1;	
							nx_state = s1263;
						end
					else if( ~x5 && ~x6 && x8 && ~x9 && ~x21 && x7 )
						begin
							y6 = 1'b1;	y30 = 1'b1;	y31 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s1263;
						end
					else if( ~x5 && ~x6 && x8 && ~x9 && ~x21 && ~x7 )
						begin
							y6 = 1'b1;	y29 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	y32 = 1'b1;	
							nx_state = s1263;
						end
					else if( ~x5 && ~x6 && ~x8 && x21 && x9 && x7 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x5 && ~x6 && ~x8 && x21 && x9 && ~x7 )
						begin
							y6 = 1'b1;	y30 = 1'b1;	y31 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s1263;
						end
					else if( ~x5 && ~x6 && ~x8 && x21 && ~x9 && x7 )
						begin
							y6 = 1'b1;	y30 = 1'b1;	y31 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s1263;
						end
					else if( ~x5 && ~x6 && ~x8 && x21 && ~x9 && ~x7 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y32 = 1'b1;	
							nx_state = s1263;
						end
					else if( ~x5 && ~x6 && ~x8 && ~x21 && x7 && x9 )
						begin
							y6 = 1'b1;	y30 = 1'b1;	y31 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s1263;
						end
					else if( ~x5 && ~x6 && ~x8 && ~x21 && x7 && ~x9 )
						begin
							y6 = 1'b1;	y30 = 1'b1;	y31 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s1263;
						end
					else if( ~x5 && ~x6 && ~x8 && ~x21 && ~x7 )
						begin
							y6 = 1'b1;	y29 = 1'b1;	y30 = 1'b1;	
							y31 = 1'b1;	y32 = 1'b1;	
							nx_state = s1263;
						end
					else nx_state = s1651;
				s1652 : if( 1'b1 )
						begin
							y11 = 1'b1;	y41 = 1'b1;	y45 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s1741;
						end
					else nx_state = s1652;
				s1653 : if( x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s654;
						end
					else if( ~x5 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x5 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x5 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( ~x5 && ~x22 )
						nx_state = s1;
					else nx_state = s1653;
				s1654 : if( 1'b1 )
						begin
							y11 = 1'b1;	y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s1654;
				s1655 : if( 1'b1 )
						begin
							y28 = 1'b1;	
							nx_state = s1326;
						end
					else nx_state = s1655;
				s1656 : if( x20 )
						begin
							y6 = 1'b1;	y9 = 1'b1;	y25 = 1'b1;	
							y56 = 1'b1;	
							nx_state = s1512;
						end
					else if( ~x20 && x13 && x21 && x14 && x15 )
						begin
							y13 = 1'b1;	
							nx_state = s484;
						end
					else if( ~x20 && x13 && x21 && x14 && ~x15 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( ~x20 && x13 && x21 && x14 && ~x15 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( ~x20 && x13 && x21 && ~x14 && x15 && x17 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( ~x20 && x13 && x21 && ~x14 && x15 && x17 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( ~x20 && x13 && x21 && ~x14 && x15 && ~x17 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && x13 && x21 && ~x14 && x15 && ~x17 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && x13 && x21 && ~x14 && x15 && ~x17 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x20 && x13 && x21 && ~x14 && x15 && ~x17 && ~x10 )
						nx_state = s1;
					else if( ~x20 && x13 && x21 && ~x14 && ~x15 && x9 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( ~x20 && x13 && x21 && ~x14 && ~x15 && x9 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( ~x20 && x13 && x21 && ~x14 && ~x15 && ~x9 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && x13 && x21 && ~x14 && ~x15 && ~x9 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && x13 && x21 && ~x14 && ~x15 && ~x9 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x20 && x13 && x21 && ~x14 && ~x15 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x20 && x13 && ~x21 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							nx_state = s1213;
						end
					else if( ~x20 && ~x13 && x14 && x21 && x15 && x18 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( ~x20 && ~x13 && x14 && x21 && x15 && x18 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( ~x20 && ~x13 && x14 && x21 && x15 && ~x18 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && ~x13 && x14 && x21 && x15 && ~x18 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && ~x13 && x14 && x21 && x15 && ~x18 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x20 && ~x13 && x14 && x21 && x15 && ~x18 && ~x10 )
						nx_state = s1;
					else if( ~x20 && ~x13 && x14 && x21 && ~x15 && x19 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else if( ~x20 && ~x13 && x14 && x21 && ~x15 && x19 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1206;
						end
					else if( ~x20 && ~x13 && x14 && x21 && ~x15 && ~x19 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && ~x13 && x14 && x21 && ~x15 && ~x19 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && ~x13 && x14 && x21 && ~x15 && ~x19 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x20 && ~x13 && x14 && x21 && ~x15 && ~x19 && ~x10 )
						nx_state = s1;
					else if( ~x20 && ~x13 && x14 && ~x21 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y22 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s722;
						end
					else if( ~x20 && ~x13 && ~x14 && x21 && x15 && x5 )
						begin
							y14 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x20 && ~x13 && ~x14 && x21 && x15 && ~x5 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1207;
						end
					else if( ~x20 && ~x13 && ~x14 && x21 && ~x15 && x7 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1208;
						end
					else if( ~x20 && ~x13 && ~x14 && x21 && ~x15 && ~x7 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1209;
						end
					else if( ~x20 && ~x13 && ~x14 && ~x21 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && ~x13 && ~x14 && ~x21 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && ~x13 && ~x14 && ~x21 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x20 && ~x13 && ~x14 && ~x21 && ~x10 )
						nx_state = s1;
					else nx_state = s1656;
				s1657 : if( x20 && x14 && x15 )
						begin
							y6 = 1'b1;	y11 = 1'b1;	y26 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1307;
						end
					else if( x20 && x14 && ~x15 )
						begin
							y6 = 1'b1;	y11 = 1'b1;	y42 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1068;
						end
					else if( x20 && ~x14 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y44 = 1'b1;	
							y45 = 1'b1;	y49 = 1'b1;	
							nx_state = s1482;
						end
					else if( ~x20 && x21 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1259;
						end
					else if( ~x20 && ~x21 && x13 )
						begin
							y6 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							nx_state = s1213;
						end
					else if( ~x20 && ~x21 && ~x13 && x14 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y22 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s722;
						end
					else if( ~x20 && ~x21 && ~x13 && ~x14 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && ~x21 && ~x13 && ~x14 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x20 && ~x21 && ~x13 && ~x14 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x20 && ~x21 && ~x13 && ~x14 && ~x10 )
						nx_state = s1;
					else nx_state = s1657;
				s1658 : if( 1'b1 )
						begin
							y15 = 1'b1;	
							nx_state = s885;
						end
					else nx_state = s1658;
				s1659 : if( 1'b1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1527;
						end
					else nx_state = s1659;
				s1660 : if( 1'b1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s1657;
						end
					else nx_state = s1660;
				s1661 : if( x65 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1742;
						end
					else if( ~x65 )
						begin
							y6 = 1'b1;	y41 = 1'b1;	y43 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s1028;
						end
					else nx_state = s1661;
				s1662 : if( x16 )
						begin
							y6 = 1'b1;	y40 = 1'b1;	y41 = 1'b1;	
							y42 = 1'b1;	y50 = 1'b1;	
							nx_state = s1028;
						end
					else if( ~x16 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x16 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x16 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x16 && ~x10 )
						nx_state = s1;
					else nx_state = s1662;
				s1663 : if( 1'b1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y74 = 1'b1;	
							nx_state = s1743;
						end
					else nx_state = s1663;
				s1664 : if( x62 && x33 && x32 )
						nx_state = s1;
					else if( x62 && x33 && ~x32 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s470;
						end
					else if( x62 && ~x33 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s470;
						end
					else if( ~x62 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y30 = 1'b1;	
							nx_state = s1744;
						end
					else nx_state = s1664;
				s1665 : if( 1'b1 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y63 = 1'b1;	
							nx_state = s1046;
						end
					else nx_state = s1665;
				s1666 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s1745;
						end
					else nx_state = s1666;
				s1667 : if( 1'b1 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	y21 = 1'b1;	
							nx_state = s820;
						end
					else nx_state = s1667;
				s1668 : if( 1'b1 )
						begin
							y10 = 1'b1;	y41 = 1'b1;	y42 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s1668;
				s1669 : if( 1'b1 )
						begin
							y25 = 1'b1;	
							nx_state = s1360;
						end
					else nx_state = s1669;
				s1670 : if( 1'b1 )
						begin
							y25 = 1'b1;	
							nx_state = s1746;
						end
					else nx_state = s1670;
				s1671 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y45 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s1747;
						end
					else nx_state = s1671;
				s1672 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y8 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s654;
						end
					else nx_state = s1672;
				s1673 : if( x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y8 = 1'b1;	
							nx_state = s1748;
						end
					else if( ~x6 && x10 && x2 && x3 && x4 && x9 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x6 && x10 && x2 && x3 && x4 && x9 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x6 && x10 && x2 && x3 && x4 && x9 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x6 && x10 && x2 && x3 && x4 && x9 && ~x1 )
						nx_state = s1;
					else if( ~x6 && x10 && x2 && x3 && x4 && ~x9 && x8 )
						begin
							y45 = 1'b1;	
							nx_state = s286;
						end
					else if( ~x6 && x10 && x2 && x3 && x4 && ~x9 && ~x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x6 && x10 && x2 && x3 && ~x4 && x9 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x6 && x10 && x2 && x3 && ~x4 && ~x9 && x8 )
						begin
							y44 = 1'b1;	
							nx_state = s1138;
						end
					else if( ~x6 && x10 && x2 && x3 && ~x4 && ~x9 && ~x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x6 && x10 && x2 && ~x3 && x4 && x9 )
						begin
							y3 = 1'b1;	y18 = 1'b1;	y21 = 1'b1;	
							nx_state = s1382;
						end
					else if( ~x6 && x10 && x2 && ~x3 && x4 && ~x9 && x8 )
						begin
							y46 = 1'b1;	
							nx_state = s531;
						end
					else if( ~x6 && x10 && x2 && ~x3 && x4 && ~x9 && ~x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x6 && x10 && x2 && ~x3 && ~x4 && x9 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( ~x6 && x10 && x2 && ~x3 && ~x4 && x9 && ~x13 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x6 && x10 && x2 && ~x3 && ~x4 && x9 && ~x13 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x6 && x10 && x2 && ~x3 && ~x4 && x9 && ~x13 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x6 && x10 && x2 && ~x3 && ~x4 && x9 && ~x13 && ~x1 )
						nx_state = s1;
					else if( ~x6 && x10 && x2 && ~x3 && ~x4 && ~x9 && x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x6 && x10 && x2 && ~x3 && ~x4 && ~x9 && ~x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x6 && x10 && ~x2 && x4 && x3 && x9 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( ~x6 && x10 && ~x2 && x4 && x3 && x9 && ~x14 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x6 && x10 && ~x2 && x4 && x3 && x9 && ~x14 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x6 && x10 && ~x2 && x4 && x3 && x9 && ~x14 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x6 && x10 && ~x2 && x4 && x3 && x9 && ~x14 && ~x1 )
						nx_state = s1;
					else if( ~x6 && x10 && ~x2 && x4 && x3 && ~x9 && x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y37 = 1'b1;	
							nx_state = s1540;
						end
					else if( ~x6 && x10 && ~x2 && x4 && x3 && ~x9 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x6 && x10 && ~x2 && x4 && ~x3 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( ~x6 && x10 && ~x2 && x4 && ~x3 && ~x9 && x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x6 && x10 && ~x2 && x4 && ~x3 && ~x9 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x6 && x10 && ~x2 && ~x4 && x9 && x3 && x12 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( ~x6 && x10 && ~x2 && ~x4 && x9 && x3 && ~x12 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x6 && x10 && ~x2 && ~x4 && x9 && x3 && ~x12 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x6 && x10 && ~x2 && ~x4 && x9 && x3 && ~x12 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x6 && x10 && ~x2 && ~x4 && x9 && x3 && ~x12 && ~x1 )
						nx_state = s1;
					else if( ~x6 && x10 && ~x2 && ~x4 && x9 && ~x3 )
						begin
							y26 = 1'b1;	
							nx_state = s1197;
						end
					else if( ~x6 && x10 && ~x2 && ~x4 && ~x9 && x8 && x3 )
						begin
							y3 = 1'b1;	y18 = 1'b1;	y42 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x6 && x10 && ~x2 && ~x4 && ~x9 && x8 && ~x3 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x6 && x10 && ~x2 && ~x4 && ~x9 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x6 && ~x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y36 = 1'b1;	y40 = 1'b1;	
							nx_state = s1705;
						end
					else nx_state = s1673;
				s1674 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y13 = 1'b1;	
							y14 = 1'b1;	
							nx_state = s1749;
						end
					else nx_state = s1674;
				s1675 : if( 1'b1 )
						begin
							y42 = 1'b1;	
							nx_state = s1670;
						end
					else nx_state = s1675;
				s1676 : if( 1'b1 )
						begin
							y42 = 1'b1;	
							nx_state = s1103;
						end
					else nx_state = s1676;
				s1677 : if( x15 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s376;
						end
					else if( ~x15 )
						begin
							y58 = 1'b1;	
							nx_state = s1265;
						end
					else nx_state = s1677;
				s1678 : if( 1'b1 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s1750;
						end
					else nx_state = s1678;
				s1679 : if( 1'b1 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s1751;
						end
					else nx_state = s1679;
				s1680 : if( 1'b1 )
						begin
							y24 = 1'b1;	
							nx_state = s590;
						end
					else nx_state = s1680;
				s1681 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1752;
						end
					else nx_state = s1681;
				s1682 : if( x15 )
						begin
							y6 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1753;
						end
					else if( ~x15 )
						begin
							y6 = 1'b1;	y25 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	y45 = 1'b1;	y46 = 1'b1;	
							nx_state = s1754;
						end
					else nx_state = s1682;
				s1683 : if( x19 && x18 )
						begin
							y2 = 1'b1;	
							nx_state = s768;
						end
					else if( x19 && ~x18 )
						begin
							y23 = 1'b1;	y28 = 1'b1;	y48 = 1'b1;	
							nx_state = s1755;
						end
					else if( ~x19 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else nx_state = s1683;
				s1684 : if( 1'b1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s1186;
						end
					else nx_state = s1684;
				s1685 : if( x23 && x4 && x5 && x3 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x23 && x4 && x5 && x3 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x23 && x4 && x5 && x3 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( x23 && x4 && x5 && x3 && ~x21 )
						nx_state = s1;
					else if( x23 && x4 && x5 && ~x3 && x12 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y23 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s535;
						end
					else if( x23 && x4 && x5 && ~x3 && ~x12 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x23 && x4 && x5 && ~x3 && ~x12 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x23 && x4 && x5 && ~x3 && ~x12 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( x23 && x4 && x5 && ~x3 && ~x12 && ~x21 )
						nx_state = s1;
					else if( x23 && x4 && ~x5 && x3 )
						begin
							y6 = 1'b1;	
							nx_state = s1506;
						end
					else if( x23 && x4 && ~x5 && ~x3 && x11 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y23 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s535;
						end
					else if( x23 && x4 && ~x5 && ~x3 && ~x11 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x23 && x4 && ~x5 && ~x3 && ~x11 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x23 && x4 && ~x5 && ~x3 && ~x11 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( x23 && x4 && ~x5 && ~x3 && ~x11 && ~x21 )
						nx_state = s1;
					else if( x23 && ~x4 && x3 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s1155;
						end
					else if( x23 && ~x4 && x3 && ~x5 && x13 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y23 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s535;
						end
					else if( x23 && ~x4 && x3 && ~x5 && ~x13 && x21 && x16 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x23 && ~x4 && x3 && ~x5 && ~x13 && x21 && ~x16 && x15 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( x23 && ~x4 && x3 && ~x5 && ~x13 && x21 && ~x16 && ~x15 )
						nx_state = s1;
					else if( x23 && ~x4 && x3 && ~x5 && ~x13 && ~x21 )
						nx_state = s1;
					else if( x23 && ~x4 && ~x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y23 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s535;
						end
					else if( ~x23 && x22 && x4 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y9 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s1684;
						end
					else if( ~x23 && x22 && x4 && ~x5 )
						begin
							y6 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x23 && x22 && ~x4 )
						begin
							y6 = 1'b1;	
							nx_state = s368;
						end
					else if( ~x23 && ~x22 )
						begin
							y6 = 1'b1;	
							nx_state = s1506;
						end
					else nx_state = s1685;
				s1686 : if( 1'b1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y27 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1756;
						end
					else nx_state = s1686;
				s1687 : if( 1'b1 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s1028;
						end
					else nx_state = s1687;
				s1688 : if( x12 && x11 && x6 )
						begin
							y5 = 1'b1;	y27 = 1'b1;	y49 = 1'b1;	
							y50 = 1'b1;	
							nx_state = s1006;
						end
					else if( x12 && x11 && ~x6 && x10 )
						begin
							y47 = 1'b1;	
							nx_state = s675;
						end
					else if( x12 && x11 && ~x6 && ~x10 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y29 = 1'b1;	
							y35 = 1'b1;	y36 = 1'b1;	
							nx_state = s749;
						end
					else if( x12 && ~x11 && x6 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y27 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s749;
						end
					else if( x12 && ~x11 && ~x6 && x10 )
						begin
							y56 = 1'b1;	
							nx_state = s1007;
						end
					else if( x12 && ~x11 && ~x6 && ~x10 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y28 = 1'b1;	
							y35 = 1'b1;	y36 = 1'b1;	
							nx_state = s749;
						end
					else if( ~x12 && x11 && x6 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y14 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s1008;
						end
					else if( ~x12 && x11 && ~x6 && x10 )
						begin
							y48 = 1'b1;	
							nx_state = s1009;
						end
					else if( ~x12 && x11 && ~x6 && ~x10 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y30 = 1'b1;	
							y35 = 1'b1;	y36 = 1'b1;	
							nx_state = s749;
						end
					else if( ~x12 && ~x11 && x6 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x12 && ~x11 && x6 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x12 && ~x11 && x6 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x12 && ~x11 && x6 && ~x18 )
						nx_state = s1;
					else if( ~x12 && ~x11 && ~x6 && x10 )
						begin
							y54 = 1'b1;	
							nx_state = s525;
						end
					else if( ~x12 && ~x11 && ~x6 && ~x10 && x18 && x14 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x12 && ~x11 && ~x6 && ~x10 && x18 && ~x14 && x13 )
						begin
							y56 = 1'b1;	
							nx_state = s746;
						end
					else if( ~x12 && ~x11 && ~x6 && ~x10 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x12 && ~x11 && ~x6 && ~x10 && ~x18 )
						nx_state = s1;
					else nx_state = s1688;
				s1689 : if( 1'b1 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s296;
						end
					else nx_state = s1689;
				s1690 : if( 1'b1 )
						begin
							y3 = 1'b1;	y18 = 1'b1;	y43 = 1'b1;	
							nx_state = s1539;
						end
					else nx_state = s1690;
				s1691 : if( 1'b1 )
						begin
							y10 = 1'b1;	
							nx_state = s841;
						end
					else nx_state = s1691;
				s1692 : if( 1'b1 )
						begin
							y4 = 1'b1;	y31 = 1'b1;	y39 = 1'b1;	
							nx_state = s1757;
						end
					else nx_state = s1692;
				s1693 : if( 1'b1 )
						begin
							y4 = 1'b1;	y31 = 1'b1;	y39 = 1'b1;	
							nx_state = s1758;
						end
					else nx_state = s1693;
				s1694 : if( x8 && x9 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x8 && x9 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x8 && x9 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x8 && x9 && ~x14 )
						nx_state = s1;
					else if( x8 && ~x9 && x11 && x10 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x8 && ~x9 && x11 && x10 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x8 && ~x9 && x11 && x10 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x8 && ~x9 && x11 && x10 && ~x14 )
						nx_state = s1;
					else if( x8 && ~x9 && x11 && ~x10 )
						begin
							y2 = 1'b1;	
							nx_state = s768;
						end
					else if( x8 && ~x9 && ~x11 && x10 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y18 = 1'b1;	y20 = 1'b1;	
							nx_state = s1692;
						end
					else if( x8 && ~x9 && ~x11 && ~x10 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x8 && ~x9 && ~x11 && ~x10 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x8 && ~x9 && ~x11 && ~x10 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x8 && ~x9 && ~x11 && ~x10 && ~x14 )
						nx_state = s1;
					else if( ~x8 && x6 && x10 && x11 && x9 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x8 && x6 && x10 && x11 && x9 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x8 && x6 && x10 && x11 && x9 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( ~x8 && x6 && x10 && x11 && x9 && ~x14 )
						nx_state = s1;
					else if( ~x8 && x6 && x10 && x11 && ~x9 && x18 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s1430;
						end
					else if( ~x8 && x6 && x10 && x11 && ~x9 && ~x18 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x8 && x6 && x10 && x11 && ~x9 && ~x18 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x8 && x6 && x10 && x11 && ~x9 && ~x18 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( ~x8 && x6 && x10 && x11 && ~x9 && ~x18 && ~x14 )
						nx_state = s1;
					else if( ~x8 && x6 && x10 && ~x11 && x9 )
						begin
							y44 = 1'b1;	
							nx_state = s755;
						end
					else if( ~x8 && x6 && x10 && ~x11 && ~x9 && x17 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s1430;
						end
					else if( ~x8 && x6 && x10 && ~x11 && ~x9 && ~x17 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x8 && x6 && x10 && ~x11 && ~x9 && ~x17 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x8 && x6 && x10 && ~x11 && ~x9 && ~x17 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( ~x8 && x6 && x10 && ~x11 && ~x9 && ~x17 && ~x14 )
						nx_state = s1;
					else if( ~x8 && x6 && ~x10 && x11 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s1693;
						end
					else if( ~x8 && x6 && ~x10 && x11 && ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s1430;
						end
					else if( ~x8 && x6 && ~x10 && ~x11 && x9 && x19 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s1430;
						end
					else if( ~x8 && x6 && ~x10 && ~x11 && x9 && ~x19 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x8 && x6 && ~x10 && ~x11 && x9 && ~x19 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x8 && x6 && ~x10 && ~x11 && x9 && ~x19 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( ~x8 && x6 && ~x10 && ~x11 && x9 && ~x19 && ~x14 )
						nx_state = s1;
					else if( ~x8 && x6 && ~x10 && ~x11 && ~x9 )
						begin
							y44 = 1'b1;	
							nx_state = s1138;
						end
					else if( ~x8 && ~x6 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else nx_state = s1694;
				s1695 : if( x63 )
						begin
							y23 = 1'b1;	y29 = 1'b1;	y48 = 1'b1;	
							nx_state = s820;
						end
					else if( ~x63 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y20 = 1'b1;	
							nx_state = s1759;
						end
					else nx_state = s1695;
				s1696 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y26 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s1760;
						end
					else nx_state = s1696;
				s1697 : if( x66 && x7 && x11 && x13 && x15 && x14 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	
							nx_state = s220;
						end
					else if( x66 && x7 && x11 && x13 && x15 && ~x14 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y58 = 1'b1;	
							nx_state = s1493;
						end
					else if( x66 && x7 && x11 && x13 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y59 = 1'b1;	
							nx_state = s1494;
						end
					else if( x66 && x7 && x11 && x13 && ~x15 && ~x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y29 = 1'b1;	
							nx_state = s1495;
						end
					else if( x66 && x7 && x11 && ~x13 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && x7 && x11 && ~x13 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && x7 && x11 && ~x13 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x66 && x7 && x11 && ~x13 && ~x8 )
						nx_state = s1;
					else if( x66 && x7 && ~x11 && x12 && x15 && x13 && x14 )
						begin
							y61 = 1'b1;	
							nx_state = s1098;
						end
					else if( x66 && x7 && ~x11 && x12 && x15 && x13 && ~x14 && x16 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( x66 && x7 && ~x11 && x12 && x15 && x13 && ~x14 && ~x16 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && x7 && ~x11 && x12 && x15 && x13 && ~x14 && ~x16 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && x7 && ~x11 && x12 && x15 && x13 && ~x14 && ~x16 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x66 && x7 && ~x11 && x12 && x15 && x13 && ~x14 && ~x16 && ~x8 )
						nx_state = s1;
					else if( x66 && x7 && ~x11 && x12 && x15 && ~x13 && x14 && x18 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1078;
						end
					else if( x66 && x7 && ~x11 && x12 && x15 && ~x13 && x14 && ~x18 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && x7 && ~x11 && x12 && x15 && ~x13 && x14 && ~x18 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && x7 && ~x11 && x12 && x15 && ~x13 && x14 && ~x18 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x66 && x7 && ~x11 && x12 && x15 && ~x13 && x14 && ~x18 && ~x8 )
						nx_state = s1;
					else if( x66 && x7 && ~x11 && x12 && x15 && ~x13 && ~x14 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( x66 && x7 && ~x11 && x12 && ~x15 && x13 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( x66 && x7 && ~x11 && x12 && ~x15 && x13 && ~x14 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( x66 && x7 && ~x11 && x12 && ~x15 && x13 && ~x14 && ~x17 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && x7 && ~x11 && x12 && ~x15 && x13 && ~x14 && ~x17 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && x7 && ~x11 && x12 && ~x15 && x13 && ~x14 && ~x17 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x66 && x7 && ~x11 && x12 && ~x15 && x13 && ~x14 && ~x17 && ~x8 )
						nx_state = s1;
					else if( x66 && x7 && ~x11 && x12 && ~x15 && ~x13 && x14 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y62 = 1'b1;	
							nx_state = s1496;
						end
					else if( x66 && x7 && ~x11 && x12 && ~x15 && ~x13 && ~x14 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && x7 && ~x11 && x12 && ~x15 && ~x13 && ~x14 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x66 && x7 && ~x11 && x12 && ~x15 && ~x13 && ~x14 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x66 && x7 && ~x11 && x12 && ~x15 && ~x13 && ~x14 && ~x8 )
						nx_state = s1;
					else if( x66 && x7 && ~x11 && ~x12 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y29 = 1'b1;	
							nx_state = s1497;
						end
					else if( x66 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y28 = 1'b1;	y29 = 1'b1;	
							nx_state = s1761;
						end
					else if( ~x66 && x26 && x25 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x66 && x26 && ~x25 && x24 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x66 && x26 && ~x25 && ~x24 )
						nx_state = s1;
					else if( ~x66 && ~x26 )
						nx_state = s1;
					else nx_state = s1697;
				s1698 : if( 1'b1 )
						begin
							y44 = 1'b1;	
							nx_state = s755;
						end
					else nx_state = s1698;
				s1699 : if( x11 && x6 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( x11 && x6 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( x11 && ~x6 && x7 && x10 )
						begin
							y48 = 1'b1;	
							nx_state = s1009;
						end
					else if( x11 && ~x6 && x7 && ~x10 && x12 && x18 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y47 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s720;
						end
					else if( x11 && ~x6 && x7 && ~x10 && x12 && ~x18 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x11 && ~x6 && x7 && ~x10 && x12 && ~x18 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x11 && ~x6 && x7 && ~x10 && x12 && ~x18 && x19 && ~x14 && ~x13 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( x11 && ~x6 && x7 && ~x10 && x12 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x11 && ~x6 && x7 && ~x10 && ~x12 && x17 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y47 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s720;
						end
					else if( x11 && ~x6 && x7 && ~x10 && ~x12 && ~x17 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x11 && ~x6 && x7 && ~x10 && ~x12 && ~x17 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x11 && ~x6 && x7 && ~x10 && ~x12 && ~x17 && x19 && ~x14 && ~x13 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( x11 && ~x6 && x7 && ~x10 && ~x12 && ~x17 && ~x19 )
						nx_state = s1;
					else if( x11 && ~x6 && ~x7 && x12 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	y38 = 1'b1;	y40 = 1'b1;	
							nx_state = s720;
						end
					else if( x11 && ~x6 && ~x7 && ~x12 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	y38 = 1'b1;	y41 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x11 && x6 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x11 && ~x6 && x7 && x12 && x10 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y45 = 1'b1;	
							y49 = 1'b1;	
							nx_state = s1576;
						end
					else if( ~x11 && ~x6 && x7 && x12 && ~x10 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y47 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x11 && ~x6 && x7 && ~x12 && x10 && x16 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y47 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x11 && ~x6 && x7 && ~x12 && x10 && ~x16 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( ~x11 && ~x6 && x7 && ~x12 && x10 && ~x16 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( ~x11 && ~x6 && x7 && ~x12 && x10 && ~x16 && x19 && ~x14 && ~x13 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x11 && ~x6 && x7 && ~x12 && x10 && ~x16 && ~x19 )
						nx_state = s1;
					else if( ~x11 && ~x6 && x7 && ~x12 && ~x10 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x11 && ~x6 && ~x7 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	y38 = 1'b1;	y42 = 1'b1;	
							nx_state = s720;
						end
					else nx_state = s1699;
				s1700 : if( x65 )
						begin
							y42 = 1'b1;	
							nx_state = s1630;
						end
					else if( ~x65 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s1762;
						end
					else nx_state = s1700;
				s1701 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else nx_state = s1701;
				s1702 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y26 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1314;
						end
					else nx_state = s1702;
				s1703 : if( 1'b1 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s1763;
						end
					else nx_state = s1703;
				s1704 : if( x19 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1564;
						end
					else if( ~x19 && x11 )
						begin
							y28 = 1'b1;	
							nx_state = s1565;
						end
					else if( ~x19 && ~x11 )
						begin
							y29 = 1'b1;	
							nx_state = s1017;
						end
					else nx_state = s1704;
				s1705 : if( x2 && x3 && x4 && x9 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x2 && x3 && x4 && x9 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x2 && x3 && x4 && x9 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x2 && x3 && x4 && x9 && ~x1 )
						nx_state = s1;
					else if( x2 && x3 && x4 && ~x9 && x8 )
						begin
							y45 = 1'b1;	
							nx_state = s286;
						end
					else if( x2 && x3 && x4 && ~x9 && ~x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x2 && x3 && ~x4 && x9 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s602;
						end
					else if( x2 && x3 && ~x4 && x9 && ~x6 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( x2 && x3 && ~x4 && ~x9 && x8 )
						begin
							y44 = 1'b1;	
							nx_state = s1138;
						end
					else if( x2 && x3 && ~x4 && ~x9 && ~x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x2 && ~x3 && x4 && x9 )
						begin
							y3 = 1'b1;	y18 = 1'b1;	y21 = 1'b1;	
							nx_state = s1382;
						end
					else if( x2 && ~x3 && x4 && ~x9 && x8 )
						begin
							y46 = 1'b1;	
							nx_state = s531;
						end
					else if( x2 && ~x3 && x4 && ~x9 && ~x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x2 && ~x3 && ~x4 && x9 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( x2 && ~x3 && ~x4 && x9 && ~x13 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x2 && ~x3 && ~x4 && x9 && ~x13 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( x2 && ~x3 && ~x4 && x9 && ~x13 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( x2 && ~x3 && ~x4 && x9 && ~x13 && ~x1 )
						nx_state = s1;
					else if( x2 && ~x3 && ~x4 && ~x9 && x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( x2 && ~x3 && ~x4 && ~x9 && ~x8 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x2 && x4 && x3 && x9 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( ~x2 && x4 && x3 && x9 && ~x14 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x2 && x4 && x3 && x9 && ~x14 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x2 && x4 && x3 && x9 && ~x14 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x2 && x4 && x3 && x9 && ~x14 && ~x1 )
						nx_state = s1;
					else if( ~x2 && x4 && x3 && ~x9 && x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y37 = 1'b1;	
							nx_state = s1540;
						end
					else if( ~x2 && x4 && x3 && ~x9 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x2 && x4 && ~x3 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( ~x2 && x4 && ~x3 && ~x9 && x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x2 && x4 && ~x3 && ~x9 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x2 && ~x4 && x9 && x3 && x12 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( ~x2 && ~x4 && x9 && x3 && ~x12 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x2 && ~x4 && x9 && x3 && ~x12 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x2 && ~x4 && x9 && x3 && ~x12 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x2 && ~x4 && x9 && x3 && ~x12 && ~x1 )
						nx_state = s1;
					else if( ~x2 && ~x4 && x9 && ~x3 )
						begin
							y26 = 1'b1;	
							nx_state = s1197;
						end
					else if( ~x2 && ~x4 && ~x9 && x8 && x3 )
						begin
							y3 = 1'b1;	y18 = 1'b1;	y42 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x2 && ~x4 && ~x9 && x8 && ~x3 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x2 && ~x4 && ~x9 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	y38 = 1'b1;	
							nx_state = s1539;
						end
					else nx_state = s1705;
				s1706 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y49 = 1'b1;	
							y50 = 1'b1;	
							nx_state = s1764;
						end
					else nx_state = s1706;
				s1707 : if( x12 )
						begin
							y61 = 1'b1;	
							nx_state = s1098;
						end
					else if( ~x12 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x12 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x12 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x12 && ~x15 )
						nx_state = s1;
					else nx_state = s1707;
				s1708 : if( 1'b1 )
						begin
							y5 = 1'b1;	y19 = 1'b1;	y25 = 1'b1;	
							y27 = 1'b1;	y30 = 1'b1;	
							nx_state = s1765;
						end
					else nx_state = s1708;
				s1709 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y26 = 1'b1;	
							nx_state = s1766;
						end
					else nx_state = s1709;
				s1710 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y55 = 1'b1;	
							y63 = 1'b1;	
							nx_state = s1400;
						end
					else nx_state = s1710;
				s1711 : if( 1'b1 )
						begin
							y3 = 1'b1;	y26 = 1'b1;	y55 = 1'b1;	
							y62 = 1'b1;	
							nx_state = s1400;
						end
					else nx_state = s1711;
				s1712 : if( x63 )
						begin
							y24 = 1'b1;	
							nx_state = s1317;
						end
					else if( ~x63 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y31 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s1400;
						end
					else nx_state = s1712;
				s1713 : if( x12 )
						begin
							y9 = 1'b1;	
							nx_state = s967;
						end
					else if( ~x12 && x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x12 && x15 && ~x16 && x17 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x12 && x15 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x12 && ~x15 )
						nx_state = s1;
					else nx_state = s1713;
				s1714 : if( 1'b1 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y19 = 1'b1;	
							y25 = 1'b1;	y30 = 1'b1;	
							nx_state = s1400;
						end
					else nx_state = s1714;
				s1715 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y54 = 1'b1;	
							y55 = 1'b1;	
							nx_state = s1400;
						end
					else nx_state = s1715;
				s1716 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y53 = 1'b1;	
							y55 = 1'b1;	
							nx_state = s1400;
						end
					else nx_state = s1716;
				s1717 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y28 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s1417;
						end
					else nx_state = s1717;
				s1718 : if( x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s1583;
						end
					else if( ~x5 && x7 && x11 && x13 && x15 && x14 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	
							nx_state = s220;
						end
					else if( ~x5 && x7 && x11 && x13 && x15 && ~x14 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y58 = 1'b1;	
							nx_state = s1493;
						end
					else if( ~x5 && x7 && x11 && x13 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y59 = 1'b1;	
							nx_state = s1494;
						end
					else if( ~x5 && x7 && x11 && x13 && ~x15 && ~x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y29 = 1'b1;	
							nx_state = s1495;
						end
					else if( ~x5 && x7 && x11 && ~x13 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x5 && x7 && x11 && ~x13 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x5 && x7 && x11 && ~x13 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x5 && x7 && x11 && ~x13 && ~x8 )
						nx_state = s1;
					else if( ~x5 && x7 && ~x11 && x12 && x15 && x13 && x14 )
						begin
							y61 = 1'b1;	
							nx_state = s1098;
						end
					else if( ~x5 && x7 && ~x11 && x12 && x15 && x13 && ~x14 && x16 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x5 && x7 && ~x11 && x12 && x15 && x13 && ~x14 && ~x16 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x5 && x7 && ~x11 && x12 && x15 && x13 && ~x14 && ~x16 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x5 && x7 && ~x11 && x12 && x15 && x13 && ~x14 && ~x16 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x5 && x7 && ~x11 && x12 && x15 && x13 && ~x14 && ~x16 && ~x8 )
						nx_state = s1;
					else if( ~x5 && x7 && ~x11 && x12 && x15 && ~x13 && x14 && x18 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1078;
						end
					else if( ~x5 && x7 && ~x11 && x12 && x15 && ~x13 && x14 && ~x18 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x5 && x7 && ~x11 && x12 && x15 && ~x13 && x14 && ~x18 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x5 && x7 && ~x11 && x12 && x15 && ~x13 && x14 && ~x18 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x5 && x7 && ~x11 && x12 && x15 && ~x13 && x14 && ~x18 && ~x8 )
						nx_state = s1;
					else if( ~x5 && x7 && ~x11 && x12 && x15 && ~x13 && ~x14 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x5 && x7 && ~x11 && x12 && ~x15 && x13 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x5 && x7 && ~x11 && x12 && ~x15 && x13 && ~x14 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x5 && x7 && ~x11 && x12 && ~x15 && x13 && ~x14 && ~x17 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x5 && x7 && ~x11 && x12 && ~x15 && x13 && ~x14 && ~x17 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x5 && x7 && ~x11 && x12 && ~x15 && x13 && ~x14 && ~x17 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x5 && x7 && ~x11 && x12 && ~x15 && x13 && ~x14 && ~x17 && ~x8 )
						nx_state = s1;
					else if( ~x5 && x7 && ~x11 && x12 && ~x15 && ~x13 && x14 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y62 = 1'b1;	
							nx_state = s1496;
						end
					else if( ~x5 && x7 && ~x11 && x12 && ~x15 && ~x13 && ~x14 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x5 && x7 && ~x11 && x12 && ~x15 && ~x13 && ~x14 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x5 && x7 && ~x11 && x12 && ~x15 && ~x13 && ~x14 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x5 && x7 && ~x11 && x12 && ~x15 && ~x13 && ~x14 && ~x8 )
						nx_state = s1;
					else if( ~x5 && x7 && ~x11 && ~x12 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y29 = 1'b1;	
							nx_state = s1497;
						end
					else if( ~x5 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y28 = 1'b1;	y29 = 1'b1;	
							nx_state = s1761;
						end
					else nx_state = s1718;
				s1719 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y42 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s1767;
						end
					else nx_state = s1719;
				s1720 : if( x14 && x13 )
						begin
							y5 = 1'b1;	y29 = 1'b1;	y36 = 1'b1;	
							y38 = 1'b1;	y53 = 1'b1;	
							nx_state = s1078;
						end
					else if( x14 && ~x13 && x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y48 = 1'b1;	
							y49 = 1'b1;	
							nx_state = s1768;
						end
					else if( x14 && ~x13 && ~x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y45 = 1'b1;	
							y46 = 1'b1;	
							nx_state = s1769;
						end
					else if( ~x14 && x15 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y36 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1078;
						end
					else if( ~x14 && x15 && ~x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y24 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1770;
						end
					else if( ~x14 && ~x15 && x13 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y38 = 1'b1;	
							y53 = 1'b1;	y54 = 1'b1;	
							nx_state = s1078;
						end
					else if( ~x14 && ~x15 && ~x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y24 = 1'b1;	
							y36 = 1'b1;	
							nx_state = s1771;
						end
					else nx_state = s1720;
				s1721 : if( x4 )
						begin
							y6 = 1'b1;	
							nx_state = s1506;
						end
					else if( ~x4 && x12 && x11 && x14 && x15 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y24 = 1'b1;	
							y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s1078;
						end
					else if( ~x4 && x12 && x11 && x14 && x15 && ~x13 )
						begin
							y35 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x4 && x12 && x11 && x14 && ~x15 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	y34 = 1'b1;	
							nx_state = s1078;
						end
					else if( ~x4 && x12 && x11 && x14 && ~x15 && ~x13 )
						begin
							y18 = 1'b1;	
							nx_state = s221;
						end
					else if( ~x4 && x12 && x11 && ~x14 && x13 && x15 && x9 )
						begin
							y11 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x4 && x12 && x11 && ~x14 && x13 && x15 && ~x9 && x8 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x4 && x12 && x11 && ~x14 && x13 && x15 && ~x9 && x8 && ~x10 )
						nx_state = s1;
					else if( ~x4 && x12 && x11 && ~x14 && x13 && x15 && ~x9 && ~x8 )
						nx_state = s1;
					else if( ~x4 && x12 && x11 && ~x14 && x13 && ~x15 && x10 )
						begin
							y11 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x4 && x12 && x11 && ~x14 && x13 && ~x15 && ~x10 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x4 && x12 && x11 && ~x14 && x13 && ~x15 && ~x10 && x8 && ~x9 )
						nx_state = s1;
					else if( ~x4 && x12 && x11 && ~x14 && x13 && ~x15 && ~x10 && ~x8 )
						nx_state = s1;
					else if( ~x4 && x12 && x11 && ~x14 && ~x13 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x4 && x12 && x11 && ~x14 && ~x13 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x4 && x12 && x11 && ~x14 && ~x13 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x4 && x12 && x11 && ~x14 && ~x13 && ~x8 )
						nx_state = s1;
					else if( ~x4 && x12 && ~x11 && x13 && x14 && x15 )
						begin
							y61 = 1'b1;	
							nx_state = s1098;
						end
					else if( ~x4 && x12 && ~x11 && x13 && x14 && ~x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1226;
						end
					else if( ~x4 && x12 && ~x11 && x13 && ~x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1226;
						end
					else if( ~x4 && x12 && ~x11 && ~x13 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1226;
						end
					else if( ~x4 && ~x12 && x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s1226;
						end
					else if( ~x4 && ~x12 && ~x5 && x11 && x14 && x15 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y38 = 1'b1;	
							nx_state = s1078;
						end
					else if( ~x4 && ~x12 && ~x5 && x11 && x14 && x15 && ~x13 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y38 = 1'b1;	
							y42 = 1'b1;	
							nx_state = s1078;
						end
					else if( ~x4 && ~x12 && ~x5 && x11 && x14 && ~x15 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y23 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1438;
						end
					else if( ~x4 && ~x12 && ~x5 && x11 && x14 && ~x15 && ~x13 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x4 && ~x12 && ~x5 && x11 && ~x14 && x15 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s1078;
						end
					else if( ~x4 && ~x12 && ~x5 && x11 && ~x14 && x15 && ~x13 )
						begin
							y40 = 1'b1;	
							nx_state = s751;
						end
					else if( ~x4 && ~x12 && ~x5 && x11 && ~x14 && ~x15 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y23 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s1772;
						end
					else if( ~x4 && ~x12 && ~x5 && x11 && ~x14 && ~x15 && ~x13 )
						begin
							y39 = 1'b1;	
							nx_state = s277;
						end
					else if( ~x4 && ~x12 && ~x5 && ~x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y23 = 1'b1;	
							y24 = 1'b1;	
							nx_state = s1720;
						end
					else nx_state = s1721;
				s1722 : if( 1'b1 )
						begin
							y2 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1773;
						end
					else nx_state = s1722;
				s1723 : if( 1'b1 )
						begin
							y3 = 1'b1;	y18 = 1'b1;	y48 = 1'b1;	
							nx_state = s1774;
						end
					else nx_state = s1723;
				s1724 : if( 1'b1 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y57 = 1'b1;	
							nx_state = s1775;
						end
					else nx_state = s1724;
				s1725 : if( 1'b1 )
						begin
							y2 = 1'b1;	
							nx_state = s1776;
						end
					else nx_state = s1725;
				s1726 : if( 1'b1 )
						begin
							y23 = 1'b1;	y28 = 1'b1;	y48 = 1'b1;	
							nx_state = s1777;
						end
					else nx_state = s1726;
				s1727 : if( 1'b1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s1778;
						end
					else nx_state = s1727;
				s1728 : if( x18 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s1728;
						end
					else if( ~x18 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y15 = 1'b1;	
							nx_state = s1779;
						end
					else nx_state = s1728;
				s1729 : if( x18 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s1689;
						end
					else if( ~x18 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s1729;
						end
					else nx_state = s1729;
				s1730 : if( x18 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s1780;
						end
					else if( ~x18 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s1730;
						end
					else nx_state = s1730;
				s1731 : if( x64 )
						begin
							y26 = 1'b1;	
							nx_state = s413;
						end
					else if( ~x64 && x14 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x64 && x14 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x64 && x14 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x64 && x14 && ~x23 )
						nx_state = s1;
					else if( ~x64 && ~x14 )
						begin
							y47 = 1'b1;	y53 = 1'b1;	y61 = 1'b1;	
							y71 = 1'b1;	
							nx_state = s1554;
						end
					else nx_state = s1731;
				s1732 : if( x15 )
						begin
							y46 = 1'b1;	y47 = 1'b1;	
							nx_state = s516;
						end
					else if( ~x15 && x6 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x15 && x6 && ~x7 && x8 )
						begin
							y15 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x15 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x15 && ~x6 )
						nx_state = s1;
					else nx_state = s1732;
				s1733 : if( 1'b1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y18 = 1'b1;	y20 = 1'b1;	
							nx_state = s1781;
						end
					else nx_state = s1733;
				s1734 : if( 1'b1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y18 = 1'b1;	
							y20 = 1'b1;	y42 = 1'b1;	
							nx_state = s1782;
						end
					else nx_state = s1734;
				s1735 : if( 1'b1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y6 = 1'b1;	
							y18 = 1'b1;	y20 = 1'b1;	
							nx_state = s1783;
						end
					else nx_state = s1735;
				s1736 : if( 1'b1 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y48 = 1'b1;	
							y49 = 1'b1;	
							nx_state = s1455;
						end
					else nx_state = s1736;
				s1737 : if( 1'b1 )
						begin
							y9 = 1'b1;	y18 = 1'b1;	y48 = 1'b1;	
							y54 = 1'b1;	
							nx_state = s1455;
						end
					else nx_state = s1737;
				s1738 : if( 1'b1 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s1455;
						end
					else nx_state = s1738;
				s1739 : if( x21 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y27 = 1'b1;	
							y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s1263;
						end
					else if( ~x21 && x8 && x9 )
						begin
							y6 = 1'b1;	y30 = 1'b1;	y31 = 1'b1;	
							y32 = 1'b1;	y38 = 1'b1;	
							nx_state = s1263;
						end
					else if( ~x21 && x8 && ~x9 )
						begin
							y6 = 1'b1;	y30 = 1'b1;	y31 = 1'b1;	
							y32 = 1'b1;	y38 = 1'b1;	
							nx_state = s1263;
						end
					else if( ~x21 && ~x8 )
						begin
							y6 = 1'b1;	y30 = 1'b1;	y31 = 1'b1;	
							y32 = 1'b1;	y38 = 1'b1;	
							nx_state = s1263;
						end
					else nx_state = s1739;
				s1740 : if( 1'b1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y31 = 1'b1;	
							y47 = 1'b1;	
							nx_state = s1784;
						end
					else nx_state = s1740;
				s1741 : if( x16 )
						begin
							y6 = 1'b1;	y40 = 1'b1;	y41 = 1'b1;	
							y42 = 1'b1;	y50 = 1'b1;	
							nx_state = s1028;
						end
					else if( ~x16 && x10 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x16 && x10 && ~x11 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x16 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x16 && ~x10 )
						nx_state = s1;
					else nx_state = s1741;
				s1742 : if( x11 && x10 && x2 )
						nx_state = s1;
					else if( x11 && x10 && ~x2 && x3 && x4 && x5 && x1 )
						begin
							y31 = 1'b1;	
							nx_state = s292;
						end
					else if( x11 && x10 && ~x2 && x3 && x4 && x5 && ~x1 )
						begin
							y41 = 1'b1;	y45 = 1'b1;	y46 = 1'b1;	
							nx_state = s654;
						end
					else if( x11 && x10 && ~x2 && x3 && x4 && ~x5 && x1 )
						begin
							y13 = 1'b1;	
							nx_state = s210;
						end
					else if( x11 && x10 && ~x2 && x3 && x4 && ~x5 && ~x1 )
						begin
							y39 = 1'b1;	y43 = 1'b1;	y44 = 1'b1;	
							nx_state = s654;
						end
					else if( x11 && x10 && ~x2 && x3 && ~x4 && x5 && x1 )
						begin
							y51 = 1'b1;	
							nx_state = s655;
						end
					else if( x11 && x10 && ~x2 && x3 && ~x4 && x5 && ~x1 )
						begin
							y41 = 1'b1;	y42 = 1'b1;	
							nx_state = s654;
						end
					else if( x11 && x10 && ~x2 && x3 && ~x4 && ~x5 && x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y48 = 1'b1;	
							y50 = 1'b1;	
							nx_state = s654;
						end
					else if( x11 && x10 && ~x2 && x3 && ~x4 && ~x5 && ~x1 )
						begin
							y39 = 1'b1;	y40 = 1'b1;	
							nx_state = s654;
						end
					else if( x11 && x10 && ~x2 && ~x3 && x4 && x5 && x1 && x6 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s651;
						end
					else if( x11 && x10 && ~x2 && ~x3 && x4 && x5 && x1 && ~x6 && x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s651;
						end
					else if( x11 && x10 && ~x2 && ~x3 && x4 && x5 && x1 && ~x6 && ~x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s652;
						end
					else if( x11 && x10 && ~x2 && ~x3 && x4 && x5 && ~x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y47 = 1'b1;	y48 = 1'b1;	
							nx_state = s654;
						end
					else if( x11 && x10 && ~x2 && ~x3 && x4 && ~x5 && x1 && x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s653;
						end
					else if( x11 && x10 && ~x2 && ~x3 && x4 && ~x5 && x1 && ~x6 && x7 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y19 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s653;
						end
					else if( x11 && x10 && ~x2 && ~x3 && x4 && ~x5 && x1 && ~x6 && ~x7 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s654;
						end
					else if( x11 && x10 && ~x2 && ~x3 && x4 && ~x5 && ~x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y48 = 1'b1;	y49 = 1'b1;	
							nx_state = s654;
						end
					else if( x11 && x10 && ~x2 && ~x3 && ~x4 && x1 && x5 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s654;
						end
					else if( x11 && x10 && ~x2 && ~x3 && ~x4 && x1 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y4 = 1'b1;	
							y48 = 1'b1;	
							nx_state = s654;
						end
					else if( x11 && x10 && ~x2 && ~x3 && ~x4 && ~x1 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y20 = 1'b1;	
							y32 = 1'b1;	y48 = 1'b1;	
							nx_state = s654;
						end
					else if( x11 && ~x10 )
						begin
							y28 = 1'b1;	
							nx_state = s1326;
						end
					else if( ~x11 )
						begin
							y29 = 1'b1;	
							nx_state = s1661;
						end
					else nx_state = s1742;
				s1743 : if( x14 && x6 && x8 && x7 )
						begin
							y63 = 1'b1;	
							nx_state = s483;
						end
					else if( x14 && x6 && x8 && ~x7 && x9 && x18 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y45 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s672;
						end
					else if( x14 && x6 && x8 && ~x7 && x9 && ~x18 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x14 && x6 && x8 && ~x7 && x9 && ~x18 && x20 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x14 && x6 && x8 && ~x7 && x9 && ~x18 && x20 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x14 && x6 && x8 && ~x7 && x9 && ~x18 && ~x20 )
						nx_state = s1;
					else if( x14 && x6 && x8 && ~x7 && ~x9 && x19 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y45 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s672;
						end
					else if( x14 && x6 && x8 && ~x7 && ~x9 && ~x19 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x14 && x6 && x8 && ~x7 && ~x9 && ~x19 && x20 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x14 && x6 && x8 && ~x7 && ~x9 && ~x19 && x20 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x14 && x6 && x8 && ~x7 && ~x9 && ~x19 && ~x20 )
						nx_state = s1;
					else if( x14 && x6 && ~x8 && x9 && x7 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y5 = 1'b1;	
							y74 = 1'b1;	
							nx_state = s1217;
						end
					else if( x14 && x6 && ~x8 && x9 && ~x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y45 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s672;
						end
					else if( x14 && x6 && ~x8 && ~x9 && x7 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y45 = 1'b1;	
							y64 = 1'b1;	
							nx_state = s672;
						end
					else if( x14 && x6 && ~x8 && ~x9 && x7 && ~x17 && x20 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x14 && x6 && ~x8 && ~x9 && x7 && ~x17 && x20 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s88;
						end
					else if( x14 && x6 && ~x8 && ~x9 && x7 && ~x17 && x20 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x14 && x6 && ~x8 && ~x9 && x7 && ~x17 && ~x20 )
						nx_state = s1;
					else if( x14 && x6 && ~x8 && ~x9 && ~x7 )
						begin
							y65 = 1'b1;	
							nx_state = s393;
						end
					else if( x14 && ~x6 )
						begin
							y57 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x14 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y40 = 1'b1;	y45 = 1'b1;	
							nx_state = s1218;
						end
					else nx_state = s1743;
				s1744 : if( 1'b1 )
						begin
							y9 = 1'b1;	
							nx_state = s709;
						end
					else nx_state = s1744;
				s1745 : if( 1'b1 )
						begin
							y9 = 1'b1;	
							nx_state = s1785;
						end
					else nx_state = s1745;
				s1746 : if( x64 )
						begin
							y26 = 1'b1;	
							nx_state = s1468;
						end
					else if( ~x64 && x14 && x23 && x24 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x64 && x14 && x23 && ~x24 && x25 )
						begin
							y10 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x64 && x14 && x23 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x64 && x14 && ~x23 )
						nx_state = s1;
					else if( ~x64 && ~x14 )
						begin
							y47 = 1'b1;	y55 = 1'b1;	y61 = 1'b1;	
							y71 = 1'b1;	
							nx_state = s1513;
						end
					else nx_state = s1746;
				s1747 : if( 1'b1 )
						begin
							y23 = 1'b1;	y72 = 1'b1;	y73 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s1747;
				s1748 : if( 1'b1 )
						begin
							y35 = 1'b1;	
							nx_state = s1025;
						end
					else nx_state = s1748;
				s1749 : if( x5 )
						begin
							y15 = 1'b1;	
							nx_state = s1625;
						end
					else if( ~x5 && x8 && x9 && x3 && x2 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x5 && x8 && x9 && x3 && x2 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x5 && x8 && x9 && x3 && x2 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x5 && x8 && x9 && x3 && x2 && ~x1 )
						nx_state = s1;
					else if( ~x5 && x8 && x9 && x3 && ~x2 && x4 && x17 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x5 && x8 && x9 && x3 && ~x2 && x4 && ~x17 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x5 && x8 && x9 && x3 && ~x2 && x4 && ~x17 && x1 && ~x16 )
						nx_state = s1;
					else if( ~x5 && x8 && x9 && x3 && ~x2 && x4 && ~x17 && ~x1 )
						nx_state = s1;
					else if( ~x5 && x8 && x9 && x3 && ~x2 && ~x4 && x16 )
						begin
							y17 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x5 && x8 && x9 && x3 && ~x2 && ~x4 && ~x16 && x1 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x5 && x8 && x9 && x3 && ~x2 && ~x4 && ~x16 && x1 && ~x17 )
						nx_state = s1;
					else if( ~x5 && x8 && x9 && x3 && ~x2 && ~x4 && ~x16 && ~x1 )
						nx_state = s1;
					else if( ~x5 && x8 && x9 && ~x3 && x4 && x2 )
						begin
							y32 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x5 && x8 && x9 && ~x3 && x4 && ~x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	y29 = 1'b1;	
							nx_state = s673;
						end
					else if( ~x5 && x8 && x9 && ~x3 && ~x4 && x2 )
						begin
							y33 = 1'b1;	
							nx_state = s589;
						end
					else if( ~x5 && x8 && x9 && ~x3 && ~x4 && ~x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y29 = 1'b1;	
							y30 = 1'b1;	y31 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x5 && x8 && ~x9 && x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y22 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s1712;
						end
					else if( ~x5 && x8 && ~x9 && ~x6 && x3 && x4 && x2 )
						begin
							y45 = 1'b1;	
							nx_state = s286;
						end
					else if( ~x5 && x8 && ~x9 && ~x6 && x3 && x4 && ~x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y37 = 1'b1;	
							nx_state = s1786;
						end
					else if( ~x5 && x8 && ~x9 && ~x6 && x3 && ~x4 && x2 )
						begin
							y44 = 1'b1;	
							nx_state = s1138;
						end
					else if( ~x5 && x8 && ~x9 && ~x6 && x3 && ~x4 && ~x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y37 = 1'b1;	
							y39 = 1'b1;	
							nx_state = s1595;
						end
					else if( ~x5 && x8 && ~x9 && ~x6 && ~x3 && x4 && x2 )
						begin
							y46 = 1'b1;	
							nx_state = s531;
						end
					else if( ~x5 && x8 && ~x9 && ~x6 && ~x3 && x4 && ~x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y22 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x5 && x8 && ~x9 && ~x6 && ~x3 && ~x4 && x2 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x5 && x8 && ~x9 && ~x6 && ~x3 && ~x4 && ~x2 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x5 && ~x8 && x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y22 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s1712;
						end
					else if( ~x5 && ~x8 && ~x6 && x2 && x3 && x4 && x9 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x5 && ~x8 && ~x6 && x2 && x3 && x4 && x9 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x5 && ~x8 && ~x6 && x2 && x3 && x4 && x9 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x5 && ~x8 && ~x6 && x2 && x3 && x4 && x9 && ~x1 )
						nx_state = s1;
					else if( ~x5 && ~x8 && ~x6 && x2 && x3 && x4 && ~x9 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x5 && ~x8 && ~x6 && x2 && x3 && ~x4 && x9 )
						begin
							y16 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x5 && ~x8 && ~x6 && x2 && x3 && ~x4 && ~x9 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x5 && ~x8 && ~x6 && x2 && ~x3 && x4 && x9 )
						begin
							y3 = 1'b1;	y18 = 1'b1;	y21 = 1'b1;	
							nx_state = s1382;
						end
					else if( ~x5 && ~x8 && ~x6 && x2 && ~x3 && x4 && ~x9 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x5 && ~x8 && ~x6 && x2 && ~x3 && ~x4 && x9 && x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( ~x5 && ~x8 && ~x6 && x2 && ~x3 && ~x4 && x9 && ~x13 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x5 && ~x8 && ~x6 && x2 && ~x3 && ~x4 && x9 && ~x13 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x5 && ~x8 && ~x6 && x2 && ~x3 && ~x4 && x9 && ~x13 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x5 && ~x8 && ~x6 && x2 && ~x3 && ~x4 && x9 && ~x13 && ~x1 )
						nx_state = s1;
					else if( ~x5 && ~x8 && ~x6 && x2 && ~x3 && ~x4 && ~x9 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x5 && ~x8 && ~x6 && ~x2 && x4 && x3 && x9 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( ~x5 && ~x8 && ~x6 && ~x2 && x4 && x3 && x9 && ~x14 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x5 && ~x8 && ~x6 && ~x2 && x4 && x3 && x9 && ~x14 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x5 && ~x8 && ~x6 && ~x2 && x4 && x3 && x9 && ~x14 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x5 && ~x8 && ~x6 && ~x2 && x4 && x3 && x9 && ~x14 && ~x1 )
						nx_state = s1;
					else if( ~x5 && ~x8 && ~x6 && ~x2 && x4 && x3 && ~x9 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	y40 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x5 && ~x8 && ~x6 && ~x2 && x4 && ~x3 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( ~x5 && ~x8 && ~x6 && ~x2 && x4 && ~x3 && ~x9 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	y40 = 1'b1;	
							nx_state = s1539;
						end
					else if( ~x5 && ~x8 && ~x6 && ~x2 && ~x4 && x9 && x3 && x12 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( ~x5 && ~x8 && ~x6 && ~x2 && ~x4 && x9 && x3 && ~x12 && x1 && x16 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x5 && ~x8 && ~x6 && ~x2 && ~x4 && x9 && x3 && ~x12 && x1 && ~x16 && x17 )
						begin
							y33 = 1'b1;	
							nx_state = s289;
						end
					else if( ~x5 && ~x8 && ~x6 && ~x2 && ~x4 && x9 && x3 && ~x12 && x1 && ~x16 && ~x17 )
						nx_state = s1;
					else if( ~x5 && ~x8 && ~x6 && ~x2 && ~x4 && x9 && x3 && ~x12 && ~x1 )
						nx_state = s1;
					else if( ~x5 && ~x8 && ~x6 && ~x2 && ~x4 && x9 && ~x3 )
						begin
							y26 = 1'b1;	
							nx_state = s1197;
						end
					else if( ~x5 && ~x8 && ~x6 && ~x2 && ~x4 && ~x9 )
						begin
							y5 = 1'b1;	y36 = 1'b1;	y37 = 1'b1;	
							y38 = 1'b1;	y40 = 1'b1;	
							nx_state = s1539;
						end
					else nx_state = s1749;
				s1750 : if( 1'b1 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s1787;
						end
					else nx_state = s1750;
				s1751 : if( 1'b1 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s1788;
						end
					else nx_state = s1751;
				s1752 : if( x15 && x11 && x6 && x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( x15 && x11 && x6 && ~x12 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( x15 && x11 && ~x6 && x7 && x10 )
						begin
							y48 = 1'b1;	
							nx_state = s1009;
						end
					else if( x15 && x11 && ~x6 && x7 && ~x10 && x12 && x18 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y47 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s720;
						end
					else if( x15 && x11 && ~x6 && x7 && ~x10 && x12 && ~x18 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x15 && x11 && ~x6 && x7 && ~x10 && x12 && ~x18 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x15 && x11 && ~x6 && x7 && ~x10 && x12 && ~x18 && x19 && ~x14 && ~x13 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y21 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s719;
						end
					else if( x15 && x11 && ~x6 && x7 && ~x10 && x12 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x15 && x11 && ~x6 && x7 && ~x10 && ~x12 && x17 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y47 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s720;
						end
					else if( x15 && x11 && ~x6 && x7 && ~x10 && ~x12 && ~x17 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x15 && x11 && ~x6 && x7 && ~x10 && ~x12 && ~x17 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x15 && x11 && ~x6 && x7 && ~x10 && ~x12 && ~x17 && x19 && ~x14 && ~x13 )
						begin
							y2 = 1'b1;	y31 = 1'b1;	y37 = 1'b1;	
							nx_state = s720;
						end
					else if( x15 && x11 && ~x6 && x7 && ~x10 && ~x12 && ~x17 && ~x19 )
						nx_state = s1;
					else if( x15 && x11 && ~x6 && ~x7 && x12 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	y38 = 1'b1;	y40 = 1'b1;	
							nx_state = s720;
						end
					else if( x15 && x11 && ~x6 && ~x7 && ~x12 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	y38 = 1'b1;	y41 = 1'b1;	
							nx_state = s720;
						end
					else if( x15 && ~x11 && x6 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( x15 && ~x11 && ~x6 && x7 && x12 && x10 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y45 = 1'b1;	
							y49 = 1'b1;	
							nx_state = s1576;
						end
					else if( x15 && ~x11 && ~x6 && x7 && x12 && ~x10 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y47 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s720;
						end
					else if( x15 && ~x11 && ~x6 && x7 && ~x12 && x10 && x16 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y47 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s720;
						end
					else if( x15 && ~x11 && ~x6 && x7 && ~x12 && x10 && ~x16 && x19 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x15 && ~x11 && ~x6 && x7 && ~x12 && x10 && ~x16 && x19 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s616;
						end
					else if( x15 && ~x11 && ~x6 && x7 && ~x12 && x10 && ~x16 && x19 && ~x14 && ~x13 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s720;
						end
					else if( x15 && ~x11 && ~x6 && x7 && ~x12 && x10 && ~x16 && ~x19 )
						nx_state = s1;
					else if( x15 && ~x11 && ~x6 && x7 && ~x12 && ~x10 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( x15 && ~x11 && ~x6 && ~x7 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y34 = 1'b1;	y38 = 1'b1;	y42 = 1'b1;	
							nx_state = s720;
						end
					else if( ~x15 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y33 = 1'b1;	
							y40 = 1'b1;	y47 = 1'b1;	
							nx_state = s1699;
						end
					else nx_state = s1752;
				s1753 : if( x17 )
						begin
							y43 = 1'b1;	
							nx_state = s410;
						end
					else if( ~x17 && x10 && x11 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x17 && x10 && ~x11 && x12 )
						begin
							y41 = 1'b1;	
							nx_state = s753;
						end
					else if( ~x17 && x10 && ~x11 && ~x12 )
						nx_state = s1;
					else if( ~x17 && ~x10 )
						nx_state = s1;
					else nx_state = s1753;
				s1754 : if( 1'b1 )
						begin
							y44 = 1'b1;	y48 = 1'b1;	y49 = 1'b1;	
							nx_state = s1525;
						end
					else nx_state = s1754;
				s1755 : if( 1'b1 )
						begin
							y2 = 1'b1;	
							nx_state = s1789;
						end
					else nx_state = s1755;
				s1756 : if( 1'b1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y20 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s535;
						end
					else nx_state = s1756;
				s1757 : if( x3 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x3 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x3 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x3 && ~x14 )
						nx_state = s1;
					else if( ~x3 )
						begin
							y14 = 1'b1;	y37 = 1'b1;	y43 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s1692;
						end
					else nx_state = s1757;
				s1758 : if( x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y10 = 1'b1;	
							y39 = 1'b1;	y41 = 1'b1;	
							nx_state = s1430;
						end
					else if( ~x3 )
						begin
							y14 = 1'b1;	y37 = 1'b1;	y43 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s1693;
						end
					else nx_state = s1758;
				s1759 : if( x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y7 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1790;
						end
					else if( ~x3 )
						begin
							y14 = 1'b1;	y37 = 1'b1;	y43 = 1'b1;	
							y44 = 1'b1;	
							nx_state = s1791;
						end
					else nx_state = s1759;
				s1760 : if( 1'b1 )
						begin
							y3 = 1'b1;	y13 = 1'b1;	y29 = 1'b1;	
							nx_state = s1417;
						end
					else nx_state = s1760;
				s1761 : if( x11 && x13 && x15 && x14 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	
							nx_state = s220;
						end
					else if( x11 && x13 && x15 && ~x14 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y58 = 1'b1;	
							nx_state = s1493;
						end
					else if( x11 && x13 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y59 = 1'b1;	
							nx_state = s1494;
						end
					else if( x11 && x13 && ~x15 && ~x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y29 = 1'b1;	
							nx_state = s1495;
						end
					else if( x11 && ~x13 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x11 && ~x13 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( x11 && ~x13 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x11 && ~x13 && ~x8 )
						nx_state = s1;
					else if( ~x11 && x12 && x15 && x13 && x14 )
						begin
							y61 = 1'b1;	
							nx_state = s1098;
						end
					else if( ~x11 && x12 && x15 && x13 && ~x14 && x16 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x11 && x12 && x15 && x13 && ~x14 && ~x16 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x11 && x12 && x15 && x13 && ~x14 && ~x16 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x11 && x12 && x15 && x13 && ~x14 && ~x16 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x11 && x12 && x15 && x13 && ~x14 && ~x16 && ~x8 )
						nx_state = s1;
					else if( ~x11 && x12 && x15 && ~x13 && x14 && x18 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1078;
						end
					else if( ~x11 && x12 && x15 && ~x13 && x14 && ~x18 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x11 && x12 && x15 && ~x13 && x14 && ~x18 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x11 && x12 && x15 && ~x13 && x14 && ~x18 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x11 && x12 && x15 && ~x13 && x14 && ~x18 && ~x8 )
						nx_state = s1;
					else if( ~x11 && x12 && x15 && ~x13 && ~x14 )
						begin
							y9 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x11 && x12 && ~x15 && x13 && x14 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x11 && x12 && ~x15 && x13 && ~x14 && x17 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s1346;
						end
					else if( ~x11 && x12 && ~x15 && x13 && ~x14 && ~x17 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x11 && x12 && ~x15 && x13 && ~x14 && ~x17 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x11 && x12 && ~x15 && x13 && ~x14 && ~x17 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x11 && x12 && ~x15 && x13 && ~x14 && ~x17 && ~x8 )
						nx_state = s1;
					else if( ~x11 && x12 && ~x15 && ~x13 && x14 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y62 = 1'b1;	
							nx_state = s1496;
						end
					else if( ~x11 && x12 && ~x15 && ~x13 && ~x14 && x8 && x9 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x11 && x12 && ~x15 && ~x13 && ~x14 && x8 && ~x9 && x10 )
						begin
							y64 = 1'b1;	
							nx_state = s485;
						end
					else if( ~x11 && x12 && ~x15 && ~x13 && ~x14 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x11 && x12 && ~x15 && ~x13 && ~x14 && ~x8 )
						nx_state = s1;
					else if( ~x11 && ~x12 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	y29 = 1'b1;	
							nx_state = s1497;
						end
					else nx_state = s1761;
				s1762 : if( 1'b1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s1792;
						end
					else nx_state = s1762;
				s1763 : if( 1'b1 )
						begin
							y2 = 1'b1;	y15 = 1'b1;	y31 = 1'b1;	
							nx_state = s1793;
						end
					else nx_state = s1763;
				s1764 : if( 1'b1 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y47 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s720;
						end
					else nx_state = s1764;
				s1765 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y27 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s1400;
						end
					else nx_state = s1765;
				s1766 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y13 = 1'b1;	
							y27 = 1'b1;	
							nx_state = s1697;
						end
					else nx_state = s1766;
				s1767 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y32 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1078;
						end
					else nx_state = s1767;
				s1768 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y50 = 1'b1;	
							nx_state = s1078;
						end
					else nx_state = s1768;
				s1769 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y47 = 1'b1;	
							nx_state = s1078;
						end
					else nx_state = s1769;
				s1770 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y45 = 1'b1;	
							y46 = 1'b1;	
							nx_state = s1794;
						end
					else nx_state = s1770;
				s1771 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y48 = 1'b1;	
							y49 = 1'b1;	
							nx_state = s1795;
						end
					else nx_state = s1771;
				s1772 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y36 = 1'b1;	
							y37 = 1'b1;	
							nx_state = s1796;
						end
					else nx_state = s1772;
				s1773 : if( 1'b1 )
						begin
							y2 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s1797;
						end
					else nx_state = s1773;
				s1774 : if( 1'b1 )
						begin
							y8 = 1'b1;	y54 = 1'b1;	
							nx_state = s1798;
						end
					else nx_state = s1774;
				s1775 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y32 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1078;
						end
					else nx_state = s1775;
				s1776 : if( 1'b1 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s1683;
						end
					else nx_state = s1776;
				s1777 : if( 1'b1 )
						begin
							y2 = 1'b1;	
							nx_state = s1695;
						end
					else nx_state = s1777;
				s1778 : if( x19 && x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s1616;
						end
					else if( x19 && ~x4 && x5 && x6 && x7 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s1617;
						end
					else if( x19 && ~x4 && x5 && x6 && ~x7 )
						begin
							y3 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							y27 = 1'b1;	y30 = 1'b1;	
							nx_state = s1618;
						end
					else if( x19 && ~x4 && x5 && ~x6 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1571;
						end
					else if( x19 && ~x4 && ~x5 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y15 = 1'b1;	y18 = 1'b1;	
							nx_state = s1619;
						end
					else if( ~x19 )
						begin
							y4 = 1'b1;	y20 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s1620;
						end
					else nx_state = s1778;
				s1779 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y23 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s1571;
						end
					else nx_state = s1779;
				s1780 : if( x5 )
						begin
							y5 = 1'b1;	y23 = 1'b1;	y34 = 1'b1;	
							y35 = 1'b1;	
							nx_state = s1571;
						end
					else if( ~x5 )
						begin
							y5 = 1'b1;	y23 = 1'b1;	y32 = 1'b1;	
							y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s1571;
						end
					else nx_state = s1780;
				s1781 : if( x9 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x9 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x9 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x9 && ~x19 )
						nx_state = s1;
					else if( ~x9 && x11 && x10 )
						begin
							y9 = 1'b1;	y21 = 1'b1;	y30 = 1'b1;	
							nx_state = s1799;
						end
					else if( ~x9 && x11 && ~x10 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1455;
						end
					else if( ~x9 && ~x11 && x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s1800;
						end
					else if( ~x9 && ~x11 && ~x10 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x9 && ~x11 && ~x10 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x9 && ~x11 && ~x10 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x9 && ~x11 && ~x10 && ~x19 )
						nx_state = s1;
					else nx_state = s1781;
				s1782 : if( 1'b1 )
						begin
							y9 = 1'b1;	y21 = 1'b1;	y44 = 1'b1;	
							nx_state = s1186;
						end
					else nx_state = s1782;
				s1783 : if( x10 && x9 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x10 && x9 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x10 && x9 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x10 && x9 && ~x19 )
						nx_state = s1;
					else if( x10 && ~x9 && x11 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x10 && ~x9 && x11 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( x10 && ~x9 && x11 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x10 && ~x9 && x11 && ~x19 )
						nx_state = s1;
					else if( x10 && ~x9 && ~x11 )
						begin
							y5 = 1'b1;	y18 = 1'b1;	y31 = 1'b1;	
							y36 = 1'b1;	y37 = 1'b1;	
							nx_state = s1455;
						end
					else if( ~x10 && x9 && x11 && x19 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x10 && x9 && x11 && x19 && ~x13 && x12 )
						begin
							y25 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x10 && x9 && x11 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x10 && x9 && x11 && ~x19 )
						nx_state = s1;
					else if( ~x10 && x9 && ~x11 )
						begin
							y5 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							y34 = 1'b1;	y35 = 1'b1;	
							nx_state = s1455;
						end
					else if( ~x10 && ~x9 )
						begin
							y5 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	y34 = 1'b1;	
							nx_state = s1455;
						end
					else nx_state = s1783;
				s1784 : if( 1'b1 )
						begin
							y4 = 1'b1;	y6 = 1'b1;	y27 = 1'b1;	
							y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s1263;
						end
					else nx_state = s1784;
				s1785 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y31 = 1'b1;	
							nx_state = s1720;
						end
					else nx_state = s1785;
				s1786 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y22 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1801;
						end
					else nx_state = s1786;
				s1787 : if( 1'b1 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s1802;
						end
					else nx_state = s1787;
				s1788 : if( 1'b1 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s1803;
						end
					else nx_state = s1788;
				s1789 : if( 1'b1 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	y17 = 1'b1;	
							y26 = 1'b1;	y49 = 1'b1;	
							nx_state = s873;
						end
					else nx_state = s1789;
				s1790 : if( x13 && x8 && x9 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x13 && x8 && x9 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x13 && x8 && x9 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x13 && x8 && x9 && ~x14 )
						nx_state = s1;
					else if( x13 && x8 && ~x9 && x11 && x10 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x13 && x8 && ~x9 && x11 && x10 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x13 && x8 && ~x9 && x11 && x10 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x13 && x8 && ~x9 && x11 && x10 && ~x14 )
						nx_state = s1;
					else if( x13 && x8 && ~x9 && x11 && ~x10 )
						begin
							y2 = 1'b1;	
							nx_state = s768;
						end
					else if( x13 && x8 && ~x9 && ~x11 && x10 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y18 = 1'b1;	y20 = 1'b1;	
							nx_state = s1692;
						end
					else if( x13 && x8 && ~x9 && ~x11 && ~x10 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x13 && x8 && ~x9 && ~x11 && ~x10 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x13 && x8 && ~x9 && ~x11 && ~x10 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x13 && x8 && ~x9 && ~x11 && ~x10 && ~x14 )
						nx_state = s1;
					else if( x13 && ~x8 && x6 && x10 && x11 && x9 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x13 && ~x8 && x6 && x10 && x11 && x9 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x13 && ~x8 && x6 && x10 && x11 && x9 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x13 && ~x8 && x6 && x10 && x11 && x9 && ~x14 )
						nx_state = s1;
					else if( x13 && ~x8 && x6 && x10 && x11 && ~x9 && x18 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s1430;
						end
					else if( x13 && ~x8 && x6 && x10 && x11 && ~x9 && ~x18 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x13 && ~x8 && x6 && x10 && x11 && ~x9 && ~x18 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x13 && ~x8 && x6 && x10 && x11 && ~x9 && ~x18 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x13 && ~x8 && x6 && x10 && x11 && ~x9 && ~x18 && ~x14 )
						nx_state = s1;
					else if( x13 && ~x8 && x6 && x10 && ~x11 && x9 )
						begin
							y44 = 1'b1;	
							nx_state = s755;
						end
					else if( x13 && ~x8 && x6 && x10 && ~x11 && ~x9 && x17 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s1430;
						end
					else if( x13 && ~x8 && x6 && x10 && ~x11 && ~x9 && ~x17 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x13 && ~x8 && x6 && x10 && ~x11 && ~x9 && ~x17 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x13 && ~x8 && x6 && x10 && ~x11 && ~x9 && ~x17 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x13 && ~x8 && x6 && x10 && ~x11 && ~x9 && ~x17 && ~x14 )
						nx_state = s1;
					else if( x13 && ~x8 && x6 && ~x10 && x11 && x9 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s1693;
						end
					else if( x13 && ~x8 && x6 && ~x10 && x11 && ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s1430;
						end
					else if( x13 && ~x8 && x6 && ~x10 && ~x11 && x9 && x19 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y39 = 1'b1;	
							y40 = 1'b1;	
							nx_state = s1430;
						end
					else if( x13 && ~x8 && x6 && ~x10 && ~x11 && x9 && ~x19 && x14 && x15 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x13 && ~x8 && x6 && ~x10 && ~x11 && x9 && ~x19 && x14 && ~x15 && x16 )
						begin
							y46 = 1'b1;	
							nx_state = s283;
						end
					else if( x13 && ~x8 && x6 && ~x10 && ~x11 && x9 && ~x19 && x14 && ~x15 && ~x16 )
						nx_state = s1;
					else if( x13 && ~x8 && x6 && ~x10 && ~x11 && x9 && ~x19 && ~x14 )
						nx_state = s1;
					else if( x13 && ~x8 && x6 && ~x10 && ~x11 && ~x9 )
						begin
							y44 = 1'b1;	
							nx_state = s1138;
						end
					else if( x13 && ~x8 && ~x6 )
						begin
							y2 = 1'b1;	
							nx_state = s422;
						end
					else if( ~x13 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y17 = 1'b1;	
							y27 = 1'b1;	y45 = 1'b1;	
							nx_state = s1694;
						end
					else nx_state = s1790;
				s1791 : if( 1'b1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y20 = 1'b1;	
							nx_state = s1759;
						end
					else nx_state = s1791;
				s1792 : if( x14 && x6 && x5 )
						nx_state = s1;
					else if( x14 && x6 && ~x5 && x7 && x8 )
						begin
							y46 = 1'b1;	
							nx_state = s1428;
						end
					else if( x14 && x6 && ~x5 && x7 && ~x8 && x9 )
						begin
							y3 = 1'b1;	y19 = 1'b1;	y42 = 1'b1;	
							y43 = 1'b1;	
							nx_state = s1555;
						end
					else if( x14 && x6 && ~x5 && x7 && ~x8 && ~x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( x14 && x6 && ~x5 && ~x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s1137;
						end
					else if( x14 && ~x6 )
						begin
							y46 = 1'b1;	
							nx_state = s1428;
						end
					else if( ~x14 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y40 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s1556;
						end
					else nx_state = s1792;
				s1793 : if( 1'b1 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s1804;
						end
					else nx_state = s1793;
				s1794 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y50 = 1'b1;	
							y52 = 1'b1;	
							nx_state = s1078;
						end
					else nx_state = s1794;
				s1795 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y47 = 1'b1;	
							y51 = 1'b1;	
							nx_state = s1078;
						end
					else nx_state = s1795;
				s1796 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y32 = 1'b1;	
							y38 = 1'b1;	
							nx_state = s1078;
						end
					else nx_state = s1796;
				s1797 : if( x14 )
						begin
							y22 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x14 && x22 && x21 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x14 && x22 && ~x21 && x18 )
						begin
							y52 = 1'b1;	
							nx_state = s714;
						end
					else if( ~x14 && x22 && ~x21 && ~x18 )
						nx_state = s1;
					else if( ~x14 && ~x22 )
						nx_state = s1;
					else nx_state = s1797;
				s1798 : if( 1'b1 )
						begin
							y13 = 1'b1;	y55 = 1'b1;	y56 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s1798;
				s1799 : if( 1'b1 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y21 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1805;
						end
					else nx_state = s1799;
				s1800 : if( 1'b1 )
						begin
							y9 = 1'b1;	y21 = 1'b1;	y41 = 1'b1;	
							y45 = 1'b1;	
							nx_state = s1806;
						end
					else nx_state = s1800;
				s1801 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y39 = 1'b1;	
							y41 = 1'b1;	
							nx_state = s1539;
						end
					else nx_state = s1801;
				s1802 : if( 1'b1 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s1536;
						end
					else nx_state = s1802;
				s1803 : if( 1'b1 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s1325;
						end
					else nx_state = s1803;
				s1804 : if( 1'b1 )
						begin
							y2 = 1'b1;	y15 = 1'b1;	y31 = 1'b1;	
							nx_state = s1276;
						end
					else nx_state = s1804;
				s1805 : if( 1'b1 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s1455;
						end
					else nx_state = s1805;
				s1806 : if( 1'b1 )
						begin
							y9 = 1'b1;	y21 = 1'b1;	y44 = 1'b1;	
							nx_state = s1455;
						end
					else nx_state = s1806;

			default : nx_state = 0;
		endcase
	end
endmodule
