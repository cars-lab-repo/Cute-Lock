library ieee;
use ieee.std_logic_1164.all;

entity group15m is
   port ( clk,rst,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,
	x16,x17,x18,x19,x20,x21,x22,x23,x24,x25,x26,x42,x45,x51,x59,
	x60,x61,x62,x63,x64,x65,x66,x67,x68 : in std_logic;
        y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,
	y16,y17,y18,y19,y20,y21,y22,y23,y24,y25,y26,y27,y28,y29,y30,
	y31,y32,y33,y34,y35,y36,y37,y38,y112 : out std_logic );
end group15m;

architecture ARC of group15m is

   type states_group15m is ( s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,
	s16,s17,s18,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29,s30,
	s31,s32,s33,s34,s35,s36,s37,s38,s39,s40,s41,s42,s43,s44,s45,
	s46,s47,s48,s49,s50,s51,s52,s53,s54,s55,s56,s57,s58,s59,s60,
	s61,s62,s63,s64,s65,s66,s67,s68,s69,s70,s71,s72,s73,s74,s75,
	s76,s77,s78,s79,s80,s81,s82,s83,s84,s85,s86,s87,s88,s89,s90,
	s91,s92,s93,s94,s95,s96,s97,s98,s99,s100,s101,s102,s103,s104,s105,
	s106,s107,s108,s109,s110,s111,s112,s113,s114,s115,s116,s117,s118,s119,s120,
	s121,s122,s123,s124,s125,s126,s127,s128,s129,s130,s131,s132,s133,s134,s135,
	s136,s137,s138,s139,s140,s141,s142,s143,s144,s145,s146,s147,s148,s149,s150,
	s151,s152,s153,s154,s155,s156,s157,s158,s159,s160,s161,s162,s163,s164,s165,
	s166,s167,s168,s169,s170,s171,s172,s173,s174,s175,s176,s177,s178,s179,s180,
	s181,s182,s183,s184,s185,s186,s187,s188,s189,s190,s191,s192,s193,s194,s195,
	s196,s197,s198,s199,s200,s201,s202,s203,s204,s205,s206,s207,s208,s209,s210,
	s211,s212,s213,s214,s215,s216,s217,s218,s219,s220,s221,s222,s223,s224,s225,
	s226,s227,s228,s229,s230,s231,s232,s233,s234,s235,s236,s237,s238,s239,s240,
	s241,s242,s243,s244,s245,s246,s247,s248,s249,s250,s251,s252,s253,s254,s255,
	s256,s257,s258,s259,s260,s261,s262,s263,s264,s265,s266,s267,s268,s269,s270,
	s271,s272,s273,s274,s275,s276,s277,s278,s279,s280,s281,s282,s283,s284,s285,
	s286,s287,s288,s289,s290,s291,s292,s293,s294,s295,s296,s297,s298,s299,s300,
	s301,s302,s303,s304,s305,s306,s307,s308,s309,s310,s311,s312,s313,s314,s315,
	s316,s317,s318,s319,s320,s321,s322,s323,s324,s325,s326,s327,s328,s329,s330,
	s331,s332,s333,s334,s335,s336,s337,s338,s339,s340,s341,s342,s343,s344,s345,
	s346,s347,s348,s349,s350,s351,s352,s353,s354,s355,s356,s357,s358,s359,s360,
	s361,s362,s363,s364,s365,s366,s367,s368,s369,s370,s371,s372,s373,s374,s375,
	s376,s377,s378,s379,s380,s381,s382,s383,s384,s385,s386,s387,s388,s389,s390,
	s391,s392,s393,s394,s395,s396,s397,s398,s399,s400,s401,s402,s403,s404,s405,
	s406,s407,s408,s409,s410,s411,s412,s413,s414,s415,s416,s417,s418,s419,s420,
	s421,s422 );
   signal current_group15m : states_group15m;

begin
   process (clk , rst)
   procedure proc_group15m is
   begin

	y1   <= '0' ;	y2   <= '0' ;	y3   <= '0' ;	y4   <= '0' ;
	y5   <= '0' ;	y6   <= '0' ;	y7   <= '0' ;	y8   <= '0' ;
	y9   <= '0' ;	y10  <= '0' ;	y11  <= '0' ;	y12  <= '0' ;
	y13  <= '0' ;	y14  <= '0' ;	y15  <= '0' ;	y16  <= '0' ;
	y17  <= '0' ;	y18  <= '0' ;	y19  <= '0' ;	y20  <= '0' ;
	y21  <= '0' ;	y22  <= '0' ;	y23  <= '0' ;	y24  <= '0' ;
	y25  <= '0' ;	y26  <= '0' ;	y27  <= '0' ;	y28  <= '0' ;
	y29  <= '0' ;	y30  <= '0' ;	y31  <= '0' ;	y32  <= '0' ;
	y33  <= '0' ;	y34  <= '0' ;	y35  <= '0' ;	y36  <= '0' ;
	y37  <= '0' ;	y38  <= '0' ;	y112 <= '0' ;

   case current_group15m is
   when s1 =>
      if ( x67 and x66 and x65 and x22 and x5 and x21 and x1 ) = '1' then
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s2;

      elsif ( x67 and x66 and x65 and x22 and x5 and x21 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and x65 and x22 and x5 and not x21 and x1 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x67 and x66 and x65 and x22 and x5 and not x21 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and x65 and x22 and not x5 and x6 and x1 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x67 and x66 and x65 and x22 and not x5 and x6 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and x65 and x22 and not x5 and not x6 and x1 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s5;

      elsif ( x67 and x66 and x65 and x22 and not x5 and not x6 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and x65 and not x22 and x4 and x17 and x23 and x1 ) = '1' then
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s1;

      elsif ( x67 and x66 and x65 and not x22 and x4 and x17 and x23 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and x65 and not x22 and x4 and x17 and not x23 and x1 ) = '1' then
         y3 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s6;

      elsif ( x67 and x66 and x65 and not x22 and x4 and x17 and not x23 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and x65 and not x22 and x4 and not x17 and x23 and x1 ) = '1' then
         y3 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s6;

      elsif ( x67 and x66 and x65 and not x22 and x4 and not x17 and x23 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and x65 and not x22 and x4 and not x17 and not x23 and x1 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x67 and x66 and x65 and not x22 and x4 and not x17 and not x23 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and x65 and not x22 and not x4 and x5 and x23 and x1 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s8;

      elsif ( x67 and x66 and x65 and not x22 and not x4 and x5 and x23 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and x65 and not x22 and not x4 and x5 and not x23 and x1 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y10 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s9;

      elsif ( x67 and x66 and x65 and not x22 and not x4 and x5 and not x23 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and x65 and not x22 and not x4 and not x5 and x23 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x67 and x66 and x65 and not x22 and not x4 and not x5 and x23 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and x65 and not x22 and not x4 and not x5 and not x23 and x1 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s5;

      elsif ( x67 and x66 and x65 and not x22 and not x4 and not x5 and not x23 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and not x65 and x68 and x1 and x21 and x6 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( x67 and x66 and not x65 and x68 and x1 and x21 and not x6 and x5 and x18 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x67 and x66 and not x65 and x68 and x1 and x21 and not x6 and x5 and not x18 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x67 and x66 and not x65 and x68 and x1 and x21 and not x6 and not x5 and x4 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s14;

      elsif ( x67 and x66 and not x65 and x68 and x1 and x21 and not x6 and not x5 and not x4 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s15;

      elsif ( x67 and x66 and not x65 and x68 and x1 and not x21 and x4 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( x67 and x66 and not x65 and x68 and x1 and not x21 and not x4 and x5 and x18 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x67 and x66 and not x65 and x68 and x1 and not x21 and not x4 and x5 and not x18 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x67 and x66 and not x65 and x68 and x1 and not x21 and not x4 and not x5 and x6 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x67 and x66 and not x65 and x68 and x1 and not x21 and not x4 and not x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s15;

      elsif ( x67 and x66 and not x65 and x68 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and not x65 and not x68 and x62 and x5 and x51 and x1 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s17;

      elsif ( x67 and x66 and not x65 and not x68 and x62 and x5 and x51 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and not x65 and not x68 and x62 and x5 and not x51 and x1 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s1;

      elsif ( x67 and x66 and not x65 and not x68 and x62 and x5 and not x51 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and not x65 and not x68 and x62 and not x5 and x2 and x1 ) = '1' then
         y14 <= '1' ;
         y28 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_group15m <= s18;

      elsif ( x67 and x66 and not x65 and not x68 and x62 and not x5 and x2 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and not x65 and not x68 and x62 and not x5 and not x2 and x1 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s19;

      elsif ( x67 and x66 and not x65 and not x68 and x62 and not x5 and not x2 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and x63 and x64 and x4 and x5 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s20;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and x63 and x64 and x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and x63 and x64 and not x4 and x5 and x3 ) = '1' then
         y34 <= '1' ;
         current_group15m <= s21;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and x63 and x64 and not x4 and x5 and not x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s22;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and x63 and x64 and not x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and x63 and not x64 and x2 and x1 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and x63 and not x64 and x2 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and x63 and not x64 and not x2 and x4 and x1 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and x63 and not x64 and not x2 and x4 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and x63 and not x64 and not x2 and not x4 and x1 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s22;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and x63 and not x64 and not x2 and not x4 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and not x63 and x64 and x5 and x17 and x1 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s22;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and not x63 and x64 and x5 and x17 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and not x63 and x64 and x5 and not x17 and x1 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and not x63 and x64 and x5 and not x17 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and not x63 and x64 and not x5 and x2 and x1 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and not x63 and x64 and not x5 and x2 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and not x63 and x64 and not x5 and not x2 and x1 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and not x63 and x64 and not x5 and not x2 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and not x63 and not x64 and x5 and x18 and x1 ) = '1' then
         y35 <= '1' ;
         current_group15m <= s26;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and not x63 and not x64 and x5 and x18 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and not x63 and not x64 and x5 and not x18 and x1 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and not x63 and not x64 and x5 and not x18 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and not x63 and not x64 and not x5 and x2 and x1 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and not x63 and not x64 and not x5 and x2 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and not x63 and not x64 and not x5 and not x2 and x1 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s22;

      elsif ( x67 and x66 and not x65 and not x68 and not x62 and not x63 and not x64 and not x5 and not x2 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and x65 and x68 and x21 and x7 and x1 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x67 and not x66 and x65 and x68 and x21 and x7 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and x65 and x68 and x21 and not x7 and x11 and x2 and x1 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s28;

      elsif ( x67 and not x66 and x65 and x68 and x21 and not x7 and x11 and x2 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and x65 and x68 and x21 and not x7 and x11 and not x2 and x1 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x67 and not x66 and x65 and x68 and x21 and not x7 and x11 and not x2 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and x65 and x68 and x21 and not x7 and not x11 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x67 and not x66 and x65 and x68 and x21 and not x7 and not x11 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and x22 and x23 and x9 and x1 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and x22 and x23 and x9 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and x22 and x23 and not x9 and x2 and x3 and x1 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s31;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and x22 and x23 and not x9 and x2 and x3 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and x22 and x23 and not x9 and x2 and not x3 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and x22 and x23 and not x9 and x2 and not x3 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and x22 and x23 and not x9 and not x2 and x1 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s32;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and x22 and x23 and not x9 and not x2 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and x22 and not x23 and x4 and x7 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and x22 and not x23 and x4 and not x7 and x2 and x1 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s33;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and x22 and not x23 and x4 and not x7 and x2 and not x1 ) = '1' then
         y3 <= '1' ;
         y12 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s34;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and x22 and not x23 and x4 and not x7 and not x2 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s35;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and x22 and not x23 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and not x22 and x23 and x7 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and not x22 and x23 and x7 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and not x22 and x23 and not x7 and x2 and x8 and x1 ) = '1' then
         y15 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s36;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and not x22 and x23 and not x7 and x2 and x8 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and not x22 and x23 and not x7 and x2 and not x8 and x1 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s33;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and not x22 and x23 and not x7 and x2 and not x8 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and not x22 and x23 and not x7 and not x2 and x1 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and not x22 and x23 and not x7 and not x2 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and not x22 and not x23 and x9 and x1 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and not x22 and not x23 and x9 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and not x22 and not x23 and not x9 and x2 and x3 and x1 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s31;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and not x22 and not x23 and not x9 and x2 and x3 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and not x22 and not x23 and not x9 and x2 and not x3 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and not x22 and not x23 and not x9 and x2 and not x3 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and not x22 and not x23 and not x9 and not x2 and x1 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s32;

      elsif ( x67 and not x66 and x65 and x68 and not x21 and not x22 and not x23 and not x9 and not x2 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and x65 and not x68 and x9 and x1 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s37;

      elsif ( x67 and not x66 and x65 and not x68 and x9 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and x65 and not x68 and not x9 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s38;

      elsif ( x67 and not x66 and x65 and not x68 and not x9 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and x68 and x20 and x4 and x19 and x2 ) = '1' then
         current_group15m <= s39;

      elsif ( x67 and not x66 and not x65 and x68 and x20 and x4 and x19 and not x2 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and x68 and x20 and x4 and not x19 and x2 ) = '1' then
         current_group15m <= s40;

      elsif ( x67 and not x66 and not x65 and x68 and x20 and x4 and not x19 and not x2 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and x68 and x20 and not x4 and x3 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s41;

      elsif ( x67 and not x66 and not x65 and x68 and x20 and not x4 and x3 and not x2 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and x68 and x20 and not x4 and not x3 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x67 and not x66 and not x65 and x68 and x20 and not x4 and not x3 and not x2 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and x68 and not x20 and x21 and x4 and x19 and x1 ) = '1' then
         y3 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s42;

      elsif ( x67 and not x66 and not x65 and x68 and not x20 and x21 and x4 and x19 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and x68 and not x20 and x21 and x4 and not x19 and x1 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( x67 and not x66 and not x65 and x68 and not x20 and x21 and x4 and not x19 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and x68 and not x20 and x21 and not x4 and x5 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s44;

      elsif ( x67 and not x66 and not x65 and x68 and not x20 and x21 and not x4 and x5 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and x68 and not x20 and x21 and not x4 and not x5 and x1 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( x67 and not x66 and not x65 and x68 and not x20 and x21 and not x4 and not x5 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and x68 and not x20 and not x21 and x5 and x1 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( x67 and not x66 and not x65 and x68 and not x20 and not x21 and x5 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and x68 and not x20 and not x21 and not x5 and x4 and x1 ) = '1' then
         y4 <= '1' ;
         y16 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s45;

      elsif ( x67 and not x66 and not x65 and x68 and not x20 and not x21 and not x5 and x4 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and x68 and not x20 and not x21 and not x5 and not x4 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s44;

      elsif ( x67 and not x66 and not x65 and x68 and not x20 and not x21 and not x5 and not x4 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and not x68 and x24 and x26 and x6 and x1 ) = '1' then
         y15 <= '1' ;
         y112 <= '1' ;
         current_group15m <= s46;

      elsif ( x67 and not x66 and not x65 and not x68 and x24 and x26 and x6 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and not x68 and x24 and x26 and not x6 and x5 and x1 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( x67 and not x66 and not x65 and not x68 and x24 and x26 and not x6 and x5 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and not x68 and x24 and x26 and not x6 and not x5 and x1 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( x67 and not x66 and not x65 and not x68 and x24 and x26 and not x6 and not x5 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and not x68 and x24 and not x26 and x5 and x18 and x1 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s48;

      elsif ( x67 and not x66 and not x65 and not x68 and x24 and not x26 and x5 and x18 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and not x68 and x24 and not x26 and x5 and not x18 and x1 ) = '1' then
         y12 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s49;

      elsif ( x67 and not x66 and not x65 and not x68 and x24 and not x26 and x5 and not x18 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and not x68 and x24 and not x26 and not x5 and x2 and x1 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s50;

      elsif ( x67 and not x66 and not x65 and not x68 and x24 and not x26 and not x5 and x2 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and not x68 and x24 and not x26 and not x5 and not x2 and x1 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( x67 and not x66 and not x65 and not x68 and x24 and not x26 and not x5 and not x2 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and x25 and x26 and x6 and x2 and x17 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s50;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and x25 and x26 and x6 and x2 and not x17 ) = '1' then
         y15 <= '1' ;
         y112 <= '1' ;
         current_group15m <= s46;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and x25 and x26 and x6 and not x2 and x5 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s51;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and x25 and x26 and x6 and not x2 and not x5 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s19;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and x25 and x26 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and x25 and not x26 and x3 and x17 and x1 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and x25 and not x26 and x3 and x17 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and x25 and not x26 and x3 and not x17 and x1 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s48;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and x25 and not x26 and x3 and not x17 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and x25 and not x26 and not x3 and x4 and x1 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and x25 and not x26 and not x3 and x4 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and x25 and not x26 and not x3 and not x4 and x1 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and x25 and not x26 and not x3 and not x4 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and not x25 and x26 and x6 and x1 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and not x25 and x26 and x6 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and not x25 and x26 and not x6 and x5 and x1 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and not x25 and x26 and not x6 and x5 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and not x25 and x26 and not x6 and not x5 and x1 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and not x25 and x26 and not x6 and not x5 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and not x25 and not x26 and x6 and x19 and x1 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and not x25 and not x26 and x6 and x19 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and not x25 and not x26 and x6 and not x19 and x1 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and not x25 and not x26 and x6 and not x19 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and not x25 and not x26 and not x6 and x2 and x1 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and not x25 and not x26 and not x6 and x2 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and not x25 and not x26 and not x6 and not x2 and x1 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( x67 and not x66 and not x65 and not x68 and not x24 and not x25 and not x26 and not x6 and not x2 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and x68 and x1 and x21 and x20 and x3 and x19 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x67 and x66 and x65 and x68 and x1 and x21 and x20 and x3 and not x19 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s57;

      elsif ( not x67 and x66 and x65 and x68 and x1 and x21 and x20 and not x3 and x4 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s58;

      elsif ( not x67 and x66 and x65 and x68 and x1 and x21 and x20 and not x3 and not x4 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s44;

      elsif ( not x67 and x66 and x65 and x68 and x1 and x21 and not x20 and x6 and x17 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s58;

      elsif ( not x67 and x66 and x65 and x68 and x1 and x21 and not x20 and x6 and not x17 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s59;

      elsif ( not x67 and x66 and x65 and x68 and x1 and x21 and not x20 and not x6 and x4 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s60;

      elsif ( not x67 and x66 and x65 and x68 and x1 and x21 and not x20 and not x6 and not x4 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s44;

      elsif ( not x67 and x66 and x65 and x68 and x1 and not x21 and x6 and x20 and x17 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x67 and x66 and x65 and x68 and x1 and not x21 and x6 and x20 and not x17 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s61;

      elsif ( not x67 and x66 and x65 and x68 and x1 and not x21 and x6 and not x20 and x17 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s61;

      elsif ( not x67 and x66 and x65 and x68 and x1 and not x21 and x6 and not x20 and not x17 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x67 and x66 and x65 and x68 and x1 and not x21 and not x6 and x5 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s58;

      elsif ( not x67 and x66 and x65 and x68 and x1 and not x21 and not x6 and not x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s44;

      elsif ( not x67 and x66 and x65 and x68 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and x60 and x5 and x4 and x17 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and x60 and x5 and x4 and not x17 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s63;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and x60 and x5 and not x4 and x6 ) = '1' then
         y4 <= '1' ;
         y13 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s64;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and x60 and x5 and not x4 and not x6 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s65;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and x60 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and not x60 and x62 and x59 and x19 and x1 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and not x60 and x62 and x59 and x19 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and not x60 and x62 and x59 and not x19 and x1 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s67;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and not x60 and x62 and x59 and not x19 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and not x60 and x62 and not x59 and x6 and x1 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s68;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and not x60 and x62 and not x59 and x6 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and not x60 and x62 and not x59 and not x6 and x1 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s69;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and not x60 and x62 and not x59 and not x6 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and not x60 and not x62 and x3 and x17 and x1 ) = '1' then
         current_group15m <= s70;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and not x60 and not x62 and x3 and x17 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and not x60 and not x62 and x3 and not x17 and x1 ) = '1' then
         current_group15m <= s71;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and not x60 and not x62 and x3 and not x17 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and not x60 and not x62 and not x3 and x6 and x1 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and not x60 and not x62 and not x3 and x6 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and not x60 and not x62 and not x3 and not x6 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( not x67 and x66 and x65 and not x68 and x61 and not x60 and not x62 and not x3 and not x6 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and x60 and x3 and x17 and x1 ) = '1' then
         current_group15m <= s70;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and x60 and x3 and x17 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and x60 and x3 and not x17 and x1 ) = '1' then
         current_group15m <= s71;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and x60 and x3 and not x17 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and x60 and not x3 and x6 and x1 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and x60 and not x3 and x6 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and x60 and not x3 and not x6 and x1 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and x60 and not x3 and not x6 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and not x60 and x62 and x3 and x1 ) = '1' then
         current_group15m <= s71;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and not x60 and x62 and x3 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and not x60 and x62 and not x3 and x5 and x1 ) = '1' then
         current_group15m <= s73;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and not x60 and x62 and not x3 and x5 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and not x60 and x62 and not x3 and not x5 and x15 and x16 and x1 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s74;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and not x60 and x62 and not x3 and not x5 and x15 and x16 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and not x60 and x62 and not x3 and not x5 and x15 and not x16 and x1 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s75;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and not x60 and x62 and not x3 and not x5 and x15 and not x16 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and not x60 and x62 and not x3 and not x5 and not x15 and x1 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s75;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and not x60 and x62 and not x3 and not x5 and not x15 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and not x60 and not x62 and x6 and x1 ) = '1' then
         current_group15m <= s71;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and not x60 and not x62 and x6 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and not x60 and not x62 and not x6 and x2 and x1 ) = '1' then
         current_group15m <= s73;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and not x60 and not x62 and not x6 and x2 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and not x60 and not x62 and not x6 and not x2 and x1 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( not x67 and x66 and x65 and not x68 and not x61 and not x60 and not x62 and not x6 and not x2 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and x1 and x21 and x68 and x3 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x67 and x66 and not x65 and x1 and x21 and x68 and not x3 and x18 and x19 ) = '1' then
         y25 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and x1 and x21 and x68 and not x3 and x18 and not x19 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( not x67 and x66 and not x65 and x1 and x21 and x68 and not x3 and not x18 ) = '1' then
         y2 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s79;

      elsif ( not x67 and x66 and not x65 and x1 and x21 and not x68 and x6 and x17 ) = '1' then
         current_group15m <= s40;

      elsif ( not x67 and x66 and not x65 and x1 and x21 and not x68 and x6 and not x17 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s80;

      elsif ( not x67 and x66 and not x65 and x1 and x21 and not x68 and not x6 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s81;

      elsif ( not x67 and x66 and not x65 and x1 and x21 and not x68 and not x6 and not x2 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x67 and x66 and not x65 and x1 and not x21 and x22 and x68 and x3 ) = '1' then
         y8 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s82;

      elsif ( not x67 and x66 and not x65 and x1 and not x21 and x22 and x68 and not x3 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and x1 and not x21 and x22 and not x68 and x23 and x5 and x19 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x67 and x66 and not x65 and x1 and not x21 and x22 and not x68 and x23 and x5 and not x19 ) = '1' then
         y2 <= '1' ;
         y8 <= '1' ;
         y13 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and x1 and not x21 and x22 and not x68 and x23 and not x5 and x6 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s84;

      elsif ( not x67 and x66 and not x65 and x1 and not x21 and x22 and not x68 and x23 and not x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s5;

      elsif ( not x67 and x66 and not x65 and x1 and not x21 and x22 and not x68 and not x23 and x4 and x17 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x67 and x66 and not x65 and x1 and not x21 and x22 and not x68 and not x23 and x4 and not x17 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s22;

      elsif ( not x67 and x66 and not x65 and x1 and not x21 and x22 and not x68 and not x23 and not x4 and x5 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s5;

      elsif ( not x67 and x66 and not x65 and x1 and not x21 and x22 and not x68 and not x23 and not x4 and not x5 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s85;

      elsif ( not x67 and x66 and not x65 and x1 and not x21 and not x22 and x68 and x9 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s28;

      elsif ( not x67 and x66 and not x65 and x1 and not x21 and not x22 and x68 and not x9 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( not x67 and x66 and not x65 and x1 and not x21 and not x22 and not x68 and x5 and x17 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s22;

      elsif ( not x67 and x66 and not x65 and x1 and not x21 and not x22 and not x68 and x5 and not x17 and x23 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x67 and x66 and not x65 and x1 and not x21 and not x22 and not x68 and x5 and not x17 and not x23 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x67 and x66 and not x65 and x1 and not x21 and not x22 and not x68 and not x5 and x6 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x67 and x66 and not x65 and x1 and not x21 and not x22 and not x68 and not x5 and not x6 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s5;

      elsif ( not x67 and x66 and not x65 and not x1 and x22 and x19 and x20 and x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and x22 and x19 and x20 and not x21 and x68 and x3 ) = '1' then
         y25 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and x22 and x19 and x20 and not x21 and x68 and not x3 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and x22 and x19 and x20 and not x21 and not x68 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and x22 and x19 and not x20 and x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and x22 and x19 and not x20 and not x21 and x68 and x3 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x67 and x66 and not x65 and not x1 and x22 and x19 and not x20 and not x21 and x68 and not x3 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and x22 and x19 and not x20 and not x21 and not x68 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and x22 and not x19 and x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and x22 and not x19 and not x21 and x68 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( not x67 and x66 and not x65 and not x1 and x22 and not x19 and not x21 and x68 and not x3 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and x22 and not x19 and not x21 and not x68 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and x17 and x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and x17 and not x10 and x68 and x16 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and x17 and not x10 and x68 and not x16 and x15 and x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and x17 and not x10 and x68 and not x16 and x15 and not x14 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and x17 and not x10 and x68 and not x16 and x15 and not x14 and not x3 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and x17 and not x10 and x68 and not x16 and not x15 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and x17 and not x10 and x68 and not x16 and not x15 and not x3 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and x17 and not x10 and not x68 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and not x17 and x14 and x68 and x16 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and not x17 and x14 and x68 and x16 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and not x17 and x14 and x68 and x16 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and not x17 and x14 and x68 and not x16 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and not x17 and x14 and not x68 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and not x17 and not x14 and x15 and x16 and x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and not x17 and not x14 and x15 and x16 and not x10 and x68 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and not x17 and not x14 and x15 and x16 and not x10 and x68 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and not x17 and not x14 and x15 and x16 and not x10 and x68 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and not x17 and not x14 and x15 and x16 and not x10 and x68 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and not x17 and not x14 and x15 and x16 and not x10 and not x68 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and not x17 and not x14 and x15 and not x16 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and not x17 and not x14 and not x15 and x68 and x16 and x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and not x17 and not x14 and not x15 and x68 and x16 and not x10 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and not x17 and not x14 and not x15 and x68 and x16 and not x10 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and not x17 and not x14 and not x15 and x68 and x16 and not x10 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and not x17 and not x14 and not x15 and x68 and not x16 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x66 and not x65 and not x1 and not x22 and not x21 and not x17 and not x14 and not x15 and not x68 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and x68 and x10 and x1 ) = '1' then
         y28 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s90;

      elsif ( not x67 and not x66 and x65 and x68 and x10 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and x68 and not x10 and x1 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s65;

      elsif ( not x67 and not x66 and x65 and x68 and not x10 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and x21 and x4 and x20 and x1 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x67 and not x66 and x65 and not x68 and x21 and x4 and x20 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and x21 and x4 and not x20 and x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and x21 and x4 and not x20 and not x18 and x1 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( not x67 and not x66 and x65 and not x68 and x21 and x4 and not x20 and not x18 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and x21 and not x4 and x3 and x1 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x67 and not x66 and x65 and not x68 and x21 and not x4 and x3 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and x21 and not x4 and not x3 and x1 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x67 and not x66 and x65 and not x68 and x21 and not x4 and not x3 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and x22 and x2 and x20 and x23 and x1 ) = '1' then
         y1 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s93;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and x22 and x2 and x20 and x23 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and x22 and x2 and x20 and not x23 ) = '1' then
         y28 <= '1' ;
         current_group15m <= s94;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and x22 and x2 and not x20 and x23 and x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and x22 and x2 and not x20 and x23 and not x19 and x1 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and x22 and x2 and not x20 and x23 and not x19 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and x22 and x2 and not x20 and not x23 and x4 and x19 ) = '1' then
         y1 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s93;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and x22 and x2 and not x20 and not x23 and x4 and not x19 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and x22 and x2 and not x20 and not x23 and not x4 and x3 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and x22 and x2 and not x20 and not x23 and not x4 and not x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and x22 and not x2 and x3 and x23 and x1 ) = '1' then
         y31 <= '1' ;
         current_group15m <= s96;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and x22 and not x2 and x3 and x23 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and x22 and not x2 and x3 and not x23 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and x22 and not x2 and not x3 and x23 and x1 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and x22 and not x2 and not x3 and x23 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and x22 and not x2 and not x3 and not x23 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and not x22 and x19 and x23 and x1 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and not x22 and x19 and x23 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and not x22 and x19 and not x23 and x1 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s97;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and not x22 and x19 and not x23 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and not x22 and not x19 and x4 and x23 and x18 and x1 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and not x22 and not x19 and x4 and x23 and x18 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and not x22 and not x19 and x4 and x23 and not x18 and x1 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s97;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and not x22 and not x19 and x4 and x23 and not x18 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and not x22 and not x19 and x4 and not x23 and x20 and x1 ) = '1' then
         y2 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s98;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and not x22 and not x19 and x4 and not x23 and x20 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and not x22 and not x19 and x4 and not x23 and not x20 and x1 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and not x22 and not x19 and x4 and not x23 and not x20 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and not x22 and not x19 and not x4 and x3 and x23 and x1 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and not x22 and not x19 and not x4 and x3 and x23 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and not x22 and not x19 and not x4 and x3 and not x23 and x1 ) = '1' then
         y1 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s93;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and not x22 and not x19 and not x4 and x3 and not x23 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and not x22 and not x19 and not x4 and not x3 and x1 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x67 and not x66 and x65 and not x68 and not x21 and not x22 and not x19 and not x4 and not x3 and not x1 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and not x65 and x1 and x21 and x68 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x67 and not x66 and not x65 and x1 and x21 and x68 and not x6 and x10 and x11 ) = '1' then
         y6 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s102;

      elsif ( not x67 and not x66 and not x65 and x1 and x21 and x68 and not x6 and x10 and not x11 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x67 and not x66 and not x65 and x1 and x21 and x68 and not x6 and not x10 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( not x67 and not x66 and not x65 and x1 and x21 and not x68 and x10 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s103;

      elsif ( not x67 and not x66 and not x65 and x1 and x21 and not x68 and not x10 and x12 and x11 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( not x67 and not x66 and not x65 and x1 and x21 and not x68 and not x10 and x12 and not x11 ) = '1' then
         y10 <= '1' ;
         y17 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s104;

      elsif ( not x67 and not x66 and not x65 and x1 and x21 and not x68 and not x10 and not x12 and x2 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( not x67 and not x66 and not x65 and x1 and x21 and not x68 and not x10 and not x12 and not x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and x22 and x68 and x9 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s105;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and x22 and x68 and not x9 and x10 and x18 and x19 and x11 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and x22 and x68 and not x9 and x10 and x18 and x19 and not x11 ) = '1' then
         y6 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s102;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and x22 and x68 and not x9 and x10 and x18 and not x19 and x12 and x16 and x11 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and x22 and x68 and not x9 and x10 and x18 and not x19 and x12 and x16 and not x11 ) = '1' then
         y6 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s102;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and x22 and x68 and not x9 and x10 and x18 and not x19 and x12 and not x16 and x11 ) = '1' then
         y6 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s102;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and x22 and x68 and not x9 and x10 and x18 and not x19 and x12 and not x16 and not x11 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and x22 and x68 and not x9 and x10 and x18 and not x19 and not x12 and x11 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and x22 and x68 and not x9 and x10 and x18 and not x19 and not x12 and not x11 ) = '1' then
         y6 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s102;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and x22 and x68 and not x9 and x10 and not x18 and x11 ) = '1' then
         y6 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s102;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and x22 and x68 and not x9 and x10 and not x18 and not x11 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and x22 and x68 and not x9 and not x10 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and x22 and not x68 and x3 ) = '1' then
         y8 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s106;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and x22 and not x68 and not x3 and x11 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s107;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and x22 and not x68 and not x3 and x11 and not x2 ) = '1' then
         current_group15m <= s40;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and x22 and not x68 and not x3 and not x11 and x9 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and x22 and not x68 and not x3 and not x11 and not x9 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and x68 and x11 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and x68 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and not x68 and x19 and x20 and x13 and x9 and x11 ) = '1' then
         current_group15m <= s40;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and not x68 and x19 and x20 and x13 and x9 and not x11 and x2 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and not x68 and x19 and x20 and x13 and x9 and not x11 and not x2 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and not x68 and x19 and x20 and x13 and not x9 and x8 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s108;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and not x68 and x19 and x20 and x13 and not x9 and not x8 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and not x68 and x19 and x20 and not x13 and x2 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and not x68 and x19 and x20 and not x13 and not x2 and x9 and x11 ) = '1' then
         current_group15m <= s40;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and not x68 and x19 and x20 and not x13 and not x2 and x9 and not x11 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and not x68 and x19 and x20 and not x13 and not x2 and not x9 and x8 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s108;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and not x68 and x19 and x20 and not x13 and not x2 and not x9 and not x8 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and not x68 and x19 and not x20 and x2 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and not x68 and x19 and not x20 and not x2 and x9 and x11 ) = '1' then
         current_group15m <= s40;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and not x68 and x19 and not x20 and not x2 and x9 and not x11 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and not x68 and x19 and not x20 and not x2 and not x9 and x8 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s108;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and not x68 and x19 and not x20 and not x2 and not x9 and not x8 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and not x68 and not x19 and x2 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and not x68 and not x19 and not x2 and x9 and x11 ) = '1' then
         current_group15m <= s40;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and not x68 and not x19 and not x2 and x9 and not x11 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and not x68 and not x19 and not x2 and not x9 and x8 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s108;

      elsif ( not x67 and not x66 and not x65 and x1 and not x21 and not x22 and not x68 and not x19 and not x2 and not x9 and not x8 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( not x67 and not x66 and not x65 and not x1 and x68 and x22 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and not x65 and not x1 and x68 and not x22 and x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x66 and not x65 and not x1 and x68 and not x22 and not x21 and x11 and x3 and x6 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s109;

      elsif ( not x67 and not x66 and not x65 and not x1 and x68 and not x22 and not x21 and x11 and x3 and not x6 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x67 and not x66 and not x65 and not x1 and x68 and not x22 and not x21 and x11 and not x3 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x67 and not x66 and not x65 and not x1 and x68 and not x22 and not x21 and not x11 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s2 =>
      if ( x22 ) = '1' then
         current_group15m <= s1;

      elsif ( not x22 and x15 and x8 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s8;

      elsif ( not x22 and x15 and not x8 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s111;

      elsif ( not x22 and not x15 and x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s50;

      else
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      end if;

   when s3 =>
      if ( x65 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and x16 and x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s113;

      elsif ( not x65 and x21 and x16 and not x10 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and x21 and not x16 ) = '1' then
         y5 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s115;

      else
         current_group15m <= s1;

      end if;

   when s4 =>
      if ( x65 and x67 and x66 and x22 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y10 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s9;

      elsif ( x65 and x67 and x66 and not x22 and x23 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y10 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s9;

      elsif ( x65 and x67 and x66 and not x22 and not x23 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x66 and x21 and x18 ) = '1' then
         y14 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s116;

      elsif ( x65 and x67 and not x66 and x21 and not x18 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s117;

      elsif ( x65 and x67 and not x66 and not x21 and x22 and x8 and x23 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x66 and not x21 and x22 and x8 and x23 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x66 and not x21 and x22 and x8 and x23 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x66 and not x21 and x22 and x8 and not x23 and x9 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x66 and not x21 and x22 and x8 and not x23 and not x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x66 and not x21 and x22 and x8 and not x23 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x66 and not x21 and x22 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x66 and not x21 and not x22 and x23 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x66 and not x21 and not x22 and x23 and x9 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x66 and not x21 and not x22 and x23 and x9 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x66 and not x21 and not x22 and x23 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x66 and not x21 and not x22 and not x23 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x66 and not x21 and not x22 and not x23 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x66 and not x21 and not x22 and not x23 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x66 and not x21 and not x22 and not x23 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and x68 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and not x68 and x61 and x60 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x67 and x66 and not x68 and x61 and x60 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x67 and x66 and not x68 and x61 and x60 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and not x68 and x61 and x60 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and not x68 and x61 and not x60 and x62 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x67 and x66 and not x68 and x61 and not x60 and not x62 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s118;

      elsif ( x65 and not x67 and x66 and not x68 and not x61 and x60 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s118;

      elsif ( x65 and not x67 and x66 and not x68 and not x61 and not x60 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and not x67 and not x66 and x21 and x18 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x65 and not x67 and not x66 and x21 and not x18 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x67 and not x66 and x21 and not x18 and x19 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x67 and not x66 and x21 and not x18 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x66 and x21 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x66 and not x21 and x23 and x22 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( x65 and not x67 and not x66 and not x21 and x23 and x22 and not x19 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x67 and not x66 and not x21 and x23 and x22 and not x19 and x17 and not x14 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x67 and not x66 and not x21 and x23 and x22 and not x19 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x66 and not x21 and x23 and x22 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x66 and not x21 and x23 and not x22 and x20 and x14 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x67 and not x66 and not x21 and x23 and not x22 and x20 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x67 and not x66 and not x21 and x23 and not x22 and x20 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x66 and not x21 and x23 and not x22 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x66 and not x21 and not x23 and x18 and x14 and x22 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x67 and not x66 and not x21 and not x23 and x18 and x14 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x67 and not x66 and not x21 and not x23 and x18 and not x14 and x13 and x22 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x67 and not x66 and not x21 and not x23 and x18 and not x14 and x13 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x67 and not x66 and not x21 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x66 and not x21 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x68 and x21 and x19 and x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and x68 and x21 and x19 and not x15 and x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and x68 and x21 and x19 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x68 and x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x68 and not x21 and x20 and x15 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( not x65 and x68 and not x21 and x20 and not x15 and x14 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( not x65 and x68 and not x21 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x68 and not x21 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x68 and x62 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x68 and not x62 and x63 and x17 and x13 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and not x68 and not x62 and x63 and x17 and x13 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x68 and not x62 and x63 and x17 and not x13 and x12 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and not x68 and not x62 and x63 and x17 and not x13 and x12 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x68 and not x62 and x63 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x68 and not x62 and x63 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x68 and not x62 and not x63 and x19 and x13 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x68 and not x62 and not x63 and x19 and x13 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and not x68 and not x62 and not x63 and x19 and not x13 and x12 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x68 and not x62 and not x63 and x19 and not x13 and x12 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and not x68 and not x62 and not x63 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s5 =>
      if ( x65 and x22 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x65 and not x22 ) = '1' then
         y2 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s121;

      elsif ( not x65 and x21 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and not x21 and x23 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( not x65 and not x21 and not x23 and x22 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      else
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      end if;

   when s6 =>
      if ( x22 ) = '1' then
         y9 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s111;

      else
         current_group15m <= s1;

      end if;

   when s7 =>
      if ( x65 and x67 and x66 and x22 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and x66 and not x22 and x23 and x19 and x15 and x8 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x65 and x67 and x66 and not x22 and x23 and x19 and x15 and not x8 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x65 and x67 and x66 and not x22 and x23 and x19 and not x15 and x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s50;

      elsif ( x65 and x67 and x66 and not x22 and x23 and x19 and not x15 and not x16 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s122;

      elsif ( x65 and x67 and x66 and not x22 and x23 and not x19 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x67 and x66 and not x22 and not x23 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x66 and x21 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x65 and x67 and not x66 and not x21 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and x68 and x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and x68 and not x20 and x21 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and not x67 and x66 and x68 and not x20 and x21 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and not x67 and x66 and x68 and not x20 and x21 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and x68 and not x20 and x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and x68 and not x20 and not x21 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and not x68 and x60 and x61 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x67 and x66 and not x68 and x60 and x61 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x67 and x66 and not x68 and x60 and x61 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and not x68 and x60 and x61 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and not x68 and x60 and not x61 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and not x67 and x66 and not x68 and not x60 and x61 and x62 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and not x67 and x66 and not x68 and not x60 and x61 and x62 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and not x67 and x66 and not x68 and not x60 and x61 and x62 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and not x68 and not x60 and x61 and x62 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and not x68 and not x60 and x61 and not x62 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and not x67 and x66 and not x68 and not x60 and not x61 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and not x67 and not x66 and x21 and x18 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x65 and not x67 and not x66 and x21 and not x18 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x67 and not x66 and x21 and not x18 and x19 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x67 and not x66 and x21 and not x18 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x66 and x21 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x66 and not x21 and x23 and x22 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( x65 and not x67 and not x66 and not x21 and x23 and x22 and not x19 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x67 and not x66 and not x21 and x23 and x22 and not x19 and x17 and not x14 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x67 and not x66 and not x21 and x23 and x22 and not x19 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x66 and not x21 and x23 and x22 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x66 and not x21 and x23 and not x22 and x20 and x14 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x67 and not x66 and not x21 and x23 and not x22 and x20 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x67 and not x66 and not x21 and x23 and not x22 and x20 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x66 and not x21 and x23 and not x22 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x66 and not x21 and not x23 and x18 and x14 and x22 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x67 and not x66 and not x21 and not x23 and x18 and x14 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x67 and not x66 and not x21 and not x23 and x18 and not x14 and x13 and x22 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x67 and not x66 and not x21 and not x23 and x18 and not x14 and x13 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x67 and not x66 and not x21 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x66 and not x21 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x68 and x21 and x19 and x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and x66 and x68 and x21 and x19 and not x15 and x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and x66 and x68 and x21 and x19 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x68 and x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x68 and not x21 and x20 and x15 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( not x65 and x66 and x68 and not x21 and x20 and not x15 and x14 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( not x65 and x66 and x68 and not x21 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x68 and not x21 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x68 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x21 and x22 ) = '1' then
         y10 <= '1' ;
         y17 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s104;

      else
         y2 <= '1' ;
         y6 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      end if;

   when s8 =>
      if ( x65 and x23 ) = '1' then
         y2 <= '1' ;
         y16 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s124;

      elsif ( x65 and not x23 and x18 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and not x23 and x18 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and not x23 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s9 =>
      if ( x22 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s125;

      elsif ( not x22 and x23 and x15 and x8 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( not x22 and x23 and x15 and not x8 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x22 and x23 and not x15 and x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s50;

      elsif ( not x22 and x23 and not x15 and not x16 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s122;

      else
         y2 <= '1' ;
         y16 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s124;

      end if;

   when s10 =>
      if ( x65 and x66 and x67 and x22 and x16 and x15 and x8 and x14 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x65 and x66 and x67 and x22 and x16 and x15 and x8 and not x14 and x7 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s126;

      elsif ( x65 and x66 and x67 and x22 and x16 and x15 and x8 and not x14 and not x7 and x12 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s85;

      elsif ( x65 and x66 and x67 and x22 and x16 and x15 and x8 and not x14 and not x7 and not x12 and x17 and x18 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and x67 and x22 and x16 and x15 and x8 and not x14 and not x7 and not x12 and x17 and not x18 and x19 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and x67 and x22 and x16 and x15 and x8 and not x14 and not x7 and not x12 and x17 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x67 and x22 and x16 and x15 and x8 and not x14 and not x7 and not x12 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x67 and x22 and x16 and x15 and not x8 and x14 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( x65 and x66 and x67 and x22 and x16 and x15 and not x8 and not x14 and x7 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         y12 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s127;

      elsif ( x65 and x66 and x67 and x22 and x16 and x15 and not x8 and not x14 and not x7 and x13 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s85;

      elsif ( x65 and x66 and x67 and x22 and x16 and x15 and not x8 and not x14 and not x7 and not x13 and x17 and x18 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and x67 and x22 and x16 and x15 and not x8 and not x14 and not x7 and not x13 and x17 and not x18 and x19 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and x67 and x22 and x16 and x15 and not x8 and not x14 and not x7 and not x13 and x17 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x67 and x22 and x16 and x15 and not x8 and not x14 and not x7 and not x13 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and x8 and x9 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and x8 and x9 and not x2 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and x8 and x9 and not x2 and not x4 ) = '1' then
         y4 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s111;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and x8 and not x9 and x7 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and x8 and not x9 and x7 and not x2 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and x8 and not x9 and x7 and not x2 and not x4 ) = '1' then
         y4 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s111;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and x8 and not x9 and not x7 and x17 and x18 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and x8 and not x9 and not x7 and x17 and not x18 and x19 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and x8 and not x9 and not x7 and x17 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and x8 and not x9 and not x7 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and not x8 and x7 and x11 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and not x8 and x7 and x11 and not x2 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and not x8 and x7 and x11 and not x2 and not x4 ) = '1' then
         y4 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s111;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and not x8 and x7 and not x11 and x17 and x18 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and not x8 and x7 and not x11 and x17 and not x18 and x19 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and not x8 and x7 and not x11 and x17 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and not x8 and x7 and not x11 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and not x8 and not x7 and x10 and x17 and x18 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and not x8 and not x7 and x10 and x17 and not x18 and x19 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and not x8 and not x7 and x10 and x17 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and not x8 and not x7 and x10 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and not x8 and not x7 and not x10 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and not x8 and not x7 and not x10 and not x2 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x65 and x66 and x67 and x22 and x16 and not x15 and not x8 and not x7 and not x10 and not x2 and not x4 ) = '1' then
         y4 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s111;

      elsif ( x65 and x66 and x67 and x22 and not x16 and x15 and x7 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x65 and x66 and x67 and x22 and not x16 and x15 and not x7 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( x65 and x66 and x67 and x22 and not x16 and x15 and not x7 and not x2 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x65 and x66 and x67 and x22 and not x16 and x15 and not x7 and not x2 and not x4 and x8 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s129;

      elsif ( x65 and x66 and x67 and x22 and not x16 and x15 and not x7 and not x2 and not x4 and not x8 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s111;

      elsif ( x65 and x66 and x67 and x22 and not x16 and not x15 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( x65 and x66 and x67 and x22 and not x16 and not x15 and not x2 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x65 and x66 and x67 and x22 and not x16 and not x15 and not x2 and not x4 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( x65 and x66 and x67 and not x22 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( x65 and x66 and not x67 and x21 and x20 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s131;

      elsif ( x65 and x66 and not x67 and x21 and not x20 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s132;

      elsif ( x65 and x66 and not x67 and not x21 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s132;

      elsif ( x65 and not x66 and x21 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s32;

      elsif ( x65 and not x66 and not x21 and x23 and x22 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x23 and not x22 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s31;

      elsif ( x65 and not x66 and not x21 and not x23 and x22 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s32;

      elsif ( x65 and not x66 and not x21 and not x23 and not x22 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x20 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      else
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      end if;

   when s11 =>
      if ( x65 and x66 and x60 and x61 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x66 and x60 and x61 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x66 and x60 and x61 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x66 and x60 and x61 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x66 and x60 and not x61 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and x60 and not x61 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and x60 and not x61 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x66 and x60 and not x61 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x66 and not x60 and x61 and x62 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x66 and not x60 and x61 and x62 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x66 and not x60 and x61 and x62 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x60 and x61 and x62 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x60 and x61 and not x62 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and not x60 and x61 and not x62 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and not x60 and x61 and not x62 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x66 and not x60 and x61 and not x62 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x66 and not x60 and not x61 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and not x66 and x21 and x18 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x65 and not x66 and x21 and not x18 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x21 and not x18 and x19 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x21 and not x18 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x21 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x23 and x22 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( x65 and not x66 and not x21 and x23 and x22 and not x19 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x66 and not x21 and x23 and x22 and not x19 and x17 and not x14 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x66 and not x21 and x23 and x22 and not x19 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x23 and x22 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x23 and not x22 and x20 and x14 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x66 and not x21 and x23 and not x22 and x20 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x66 and not x21 and x23 and not x22 and x20 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x23 and not x22 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x23 and x18 and x14 and x22 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x21 and not x23 and x18 and x14 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x66 and not x21 and not x23 and x18 and not x14 and x13 and x22 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x21 and not x23 and x18 and not x14 and x13 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x66 and not x21 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x68 and x5 and x18 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x65 and x68 and x5 and not x18 and x21 and x6 ) = '1' then
         current_group15m <= s11;

      elsif ( not x65 and x68 and x5 and not x18 and x21 and not x6 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x65 and x68 and x5 and not x18 and not x21 and x4 ) = '1' then
         current_group15m <= s11;

      elsif ( not x65 and x68 and x5 and not x18 and not x21 and not x4 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x65 and x68 and not x5 and x21 and x4 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s14;

      elsif ( not x65 and x68 and not x5 and x21 and not x4 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s15;

      elsif ( not x65 and x68 and not x5 and not x21 and x6 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x65 and x68 and not x5 and not x21 and not x6 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s15;

      elsif ( not x65 and not x68 and x62 and x61 and x13 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and not x68 and x62 and x61 and not x13 and x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and not x68 and x62 and x61 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x68 and x62 and not x61 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x68 and not x62 and x63 and x17 and x13 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and not x68 and not x62 and x63 and x17 and x13 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x68 and not x62 and x63 and x17 and not x13 and x12 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and not x68 and not x62 and x63 and x17 and not x13 and x12 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x68 and not x62 and x63 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x68 and not x62 and x63 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x68 and not x62 and not x63 and x19 and x13 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x68 and not x62 and not x63 and x19 and x13 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and not x68 and not x62 and not x63 and x19 and not x13 and x12 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x68 and not x62 and not x63 and x19 and not x13 and x12 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and not x68 and not x62 and not x63 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s12 =>
      if ( x65 and x67 and x66 and x22 and x17 and x18 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and x66 and x22 and x17 and not x18 and x19 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and x66 and x22 and x17 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and x66 and x22 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and x66 and not x22 and x3 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and x66 and not x22 and not x3 and x19 and x15 and x8 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x65 and x67 and x66 and not x22 and not x3 and x19 and x15 and not x8 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x65 and x67 and x66 and not x22 and not x3 and x19 and not x15 and x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s50;

      elsif ( x65 and x67 and x66 and not x22 and not x3 and x19 and not x15 and not x16 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s122;

      elsif ( x65 and x67 and x66 and not x22 and not x3 and not x19 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x67 and not x66 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and x68 and x20 and x19 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x67 and x66 and x68 and x20 and x19 and not x14 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x67 and x66 and x68 and x20 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and x68 and x20 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and x68 and not x20 and x21 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x65 and not x67 and x66 and x68 and not x20 and not x21 and x19 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x67 and x66 and x68 and not x20 and not x21 and x19 and not x14 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x67 and x66 and x68 and not x20 and not x21 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and x68 and not x20 and not x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and not x68 and x60 and x61 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x67 and x66 and not x68 and x60 and x61 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x67 and x66 and not x68 and x60 and x61 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and not x68 and x60 and x61 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and not x68 and x60 and not x61 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x67 and x66 and not x68 and x60 and not x61 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x67 and x66 and not x68 and x60 and not x61 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and not x67 and x66 and not x68 and x60 and not x61 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and not x67 and x66 and not x68 and not x60 and x61 and x62 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and not x67 and x66 and not x68 and not x60 and x61 and x62 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and not x67 and x66 and not x68 and not x60 and x61 and x62 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and not x68 and not x60 and x61 and x62 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x66 and not x68 and not x60 and x61 and not x62 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x67 and x66 and not x68 and not x60 and x61 and not x62 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x67 and x66 and not x68 and not x60 and x61 and not x62 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and not x67 and x66 and not x68 and not x60 and x61 and not x62 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and not x67 and x66 and not x68 and not x60 and not x61 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and not x67 and not x66 and x21 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x66 and not x21 and x19 and x18 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x67 and not x66 and not x21 and x19 and not x18 ) = '1' then
         current_group15m <= s12;

      elsif ( x65 and not x67 and not x66 and not x21 and not x19 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s97;

      elsif ( not x65 and x68 and x21 and x6 and x18 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x65 and x68 and x21 and x6 and not x18 ) = '1' then
         current_group15m <= s12;

      elsif ( not x65 and x68 and x21 and not x6 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x65 and x68 and not x21 and x4 and x18 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x65 and x68 and not x21 and x4 and not x18 ) = '1' then
         current_group15m <= s12;

      elsif ( not x65 and x68 and not x21 and not x4 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x65 and not x68 and x62 and x61 and x13 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and not x68 and x62 and x61 and not x13 and x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and not x68 and x62 and x61 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x68 and x62 and not x61 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x68 and not x62 and x63 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x68 and not x62 and not x63 and x64 and x16 and x8 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and not x68 and not x62 and not x63 and x64 and x16 and not x8 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x65 and not x68 and not x62 and not x63 and x64 and not x16 and x4 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x65 and not x68 and not x62 and not x63 and x64 and not x16 and not x4 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s135;

      else
         y36 <= '1' ;
         current_group15m <= s55;

      end if;

   when s13 =>
      if ( x65 and x67 and x21 and x68 and x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x65 and x67 and x21 and x68 and x8 and not x9 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x65 and x67 and x21 and x68 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and x21 and x68 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and x21 and not x68 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x67 and x21 and not x68 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x67 and x21 and not x68 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and x21 and not x68 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x21 and x68 and x23 and x22 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x21 and x68 and x23 and x22 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x21 and x68 and x23 and x22 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x21 and x68 and x23 and x22 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x21 and x68 and x23 and not x22 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x21 and x68 and x23 and not x22 and x9 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x21 and x68 and x23 and not x22 and x9 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x21 and x68 and x23 and not x22 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x21 and x68 and not x23 and x8 and x22 and x9 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x21 and x68 and not x23 and x8 and x22 and not x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x21 and x68 and not x23 and x8 and x22 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x21 and x68 and not x23 and x8 and not x22 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x21 and x68 and not x23 and x8 and not x22 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x21 and x68 and not x23 and x8 and not x22 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x21 and x68 and not x23 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x21 and not x68 and x22 and x19 and x18 and x11 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x65 and x67 and not x21 and not x68 and x22 and x19 and x18 and not x11 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x67 and not x21 and not x68 and x22 and x19 and x18 and not x11 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x67 and not x21 and not x68 and x22 and x19 and x18 and not x11 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x21 and not x68 and x22 and x19 and x18 and not x11 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x21 and not x68 and x22 and x19 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x21 and not x68 and x22 and not x19 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x67 and not x21 and not x68 and x22 and not x19 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x67 and not x21 and not x68 and x22 and not x19 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x21 and not x68 and x22 and not x19 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x21 and not x68 and not x22 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x67 and not x21 and not x68 and not x22 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x67 and not x21 and not x68 and not x22 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x21 and not x68 and not x22 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x21 and x18 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x65 and not x67 and x21 and not x18 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x67 and x21 and not x18 and x19 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x67 and x21 and not x18 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x21 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x21 and x23 and x22 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( x65 and not x67 and not x21 and x23 and x22 and not x19 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x67 and not x21 and x23 and x22 and not x19 and x17 and not x14 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x67 and not x21 and x23 and x22 and not x19 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x21 and x23 and x22 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x21 and x23 and not x22 and x20 and x14 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x67 and not x21 and x23 and not x22 and x20 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x67 and not x21 and x23 and not x22 and x20 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x21 and x23 and not x22 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x21 and not x23 and x18 and x14 and x22 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x67 and not x21 and not x23 and x18 and x14 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x67 and not x21 and not x23 and x18 and not x14 and x13 and x22 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x67 and not x21 and not x23 and x18 and not x14 and x13 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x67 and not x21 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x21 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and x68 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x68 and x62 and x61 and x13 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and x66 and x67 and not x68 and x62 and x61 and not x13 and x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and x66 and x67 and not x68 and x62 and x61 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x68 and x62 and not x61 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and x63 and x17 and x13 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and x63 and x17 and x13 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and x63 and x17 and not x13 and x12 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and x63 and x17 and not x13 and x12 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and x63 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and x63 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and not x63 and x19 and x13 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and not x63 and x19 and x13 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and not x63 and x19 and not x13 and x12 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and not x63 and x19 and not x13 and x12 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and not x63 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and not x63 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and x21 and x17 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x66 and not x67 and x21 and x17 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x66 and not x67 and x21 and x17 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and x21 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and x8 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and not x8 and x9 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and not x8 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and not x21 and not x22 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x66 and not x67 and not x21 and not x22 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x66 and not x67 and not x21 and not x22 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and not x21 and not x22 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x22 and x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x22 and not x21 and x16 and x12 and x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x22 and not x21 and x16 and x12 and not x19 and x18 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x65 and not x66 and x22 and not x21 and x16 and x12 and not x19 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x22 and not x21 and x16 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x22 and not x21 and not x16 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s14 =>
      if ( x21 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s139;

      elsif ( not x21 and x19 and x16 and x10 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s67;

      elsif ( not x21 and x19 and x16 and not x10 ) = '1' then
         y5 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s113;

      elsif ( not x21 and x19 and not x16 and x17 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x21 and x19 and not x16 and not x17 ) = '1' then
         y5 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s115;

      else
         y13 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s141;

      end if;

   when s15 =>
      if ( x65 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      else
         y1 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s142;

      end if;

   when s16 =>
      if ( x66 and x67 and x65 and x22 and x17 and x18 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and x67 and x65 and x22 and x17 and not x18 and x19 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and x67 and x65 and x22 and x17 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x67 and x65 and x22 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x67 and x65 and not x22 and x18 and x13 and x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x66 and x67 and x65 and not x22 and x18 and x13 and not x23 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x67 and x65 and not x22 and x18 and not x13 and x12 and x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x66 and x67 and x65 and not x22 and x18 and not x13 and x12 and not x23 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x67 and x65 and not x22 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x67 and x65 and not x22 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x67 and not x65 and x68 and x21 and x19 and x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and x67 and not x65 and x68 and x21 and x19 and not x15 and x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and x67 and not x65 and x68 and x21 and x19 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x67 and not x65 and x68 and x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x67 and not x65 and x68 and not x21 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s139;

      elsif ( x66 and x67 and not x65 and not x68 and x62 and x61 and x13 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x66 and x67 and not x65 and not x68 and x62 and x61 and not x13 and x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x66 and x67 and not x65 and not x68 and x62 and x61 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x67 and not x65 and not x68 and x62 and not x61 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x67 and not x65 and not x68 and not x62 and x63 and x17 and x13 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and x67 and not x65 and not x68 and not x62 and x63 and x17 and x13 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( x66 and x67 and not x65 and not x68 and not x62 and x63 and x17 and not x13 and x12 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and x67 and not x65 and not x68 and not x62 and x63 and x17 and not x13 and x12 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( x66 and x67 and not x65 and not x68 and not x62 and x63 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x67 and not x65 and not x68 and not x62 and x63 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x67 and not x65 and not x68 and not x62 and not x63 and x19 and x13 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x66 and x67 and not x65 and not x68 and not x62 and not x63 and x19 and x13 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x66 and x67 and not x65 and not x68 and not x62 and not x63 and x19 and not x13 and x12 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x66 and x67 and not x65 and not x68 and not x62 and not x63 and x19 and not x13 and x12 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x66 and x67 and not x65 and not x68 and not x62 and not x63 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x67 and not x65 and not x68 and not x62 and not x63 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and x65 and x21 and x20 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and not x67 and x65 and x21 and x20 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and not x67 and x65 and x21 and x20 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and x65 and x21 and x20 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and x65 and x21 and not x20 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and not x67 and x65 and x21 and not x20 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and not x67 and x65 and x21 and not x20 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and x65 and x21 and not x20 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and x65 and not x21 and x19 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and not x67 and x65 and not x21 and x19 and not x14 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and not x67 and x65 and not x21 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and x65 and not x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and x21 and x68 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x66 and not x67 and not x65 and x21 and x68 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x66 and not x67 and not x65 and x21 and x68 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and x21 and x68 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and x21 and not x68 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s143;

      elsif ( x66 and not x67 and not x65 and not x21 and x68 and x22 and x9 and x7 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( x66 and not x67 and not x65 and not x21 and x68 and x22 and x9 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and x68 and x22 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and x68 and not x22 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x67 and not x65 and not x21 and x68 and not x22 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x67 and not x65 and not x21 and x68 and not x22 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and x68 and not x22 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and not x68 and x23 and x22 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x66 and not x67 and not x65 and not x21 and not x68 and x23 and not x22 and x19 and x14 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( x66 and not x67 and not x65 and not x21 and not x68 and x23 and not x22 and x19 and not x14 and x13 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( x66 and not x67 and not x65 and not x21 and not x68 and x23 and not x22 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and not x68 and x23 and not x22 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and not x68 and not x23 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x66 and x65 and x21 and x67 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and x21 and x67 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and x21 and x67 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and x21 and x67 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and x21 and not x67 and x18 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x66 and x65 and x21 and not x67 and not x18 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and x21 and not x67 and not x18 and x19 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and x21 and not x67 and not x18 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and x21 and not x67 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and x67 and x22 and x18 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and not x21 and x67 and x22 and x18 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and not x21 and x67 and x22 and x18 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and x67 and x22 and x18 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and x67 and x22 and not x18 and x10 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s146;

      elsif ( not x66 and x65 and not x21 and x67 and x22 and not x18 and not x10 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and not x21 and x67 and x22 and not x18 and not x10 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and not x21 and x67 and x22 and not x18 and not x10 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and x67 and x22 and not x18 and not x10 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and x67 and not x22 and x19 and x10 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s146;

      elsif ( not x66 and x65 and not x21 and x67 and not x22 and x19 and not x10 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and not x21 and x67 and not x22 and x19 and not x10 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and not x21 and x67 and not x22 and x19 and not x10 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and x67 and not x22 and x19 and not x10 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and x67 and not x22 and not x19 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and not x21 and x67 and not x22 and not x19 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and not x21 and x67 and not x22 and not x19 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and x67 and not x22 and not x19 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x67 and x23 and x22 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( not x66 and x65 and not x21 and not x67 and x23 and x22 and not x19 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( not x66 and x65 and not x21 and not x67 and x23 and x22 and not x19 and x17 and not x14 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( not x66 and x65 and not x21 and not x67 and x23 and x22 and not x19 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x67 and x23 and x22 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x67 and x23 and not x22 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s147;

      elsif ( not x66 and x65 and not x21 and not x67 and not x23 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s147;

      elsif ( not x66 and not x65 and x20 and x18 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x66 and not x65 and x20 and x18 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x66 and not x65 and x20 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x20 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x20 and x21 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x66 and not x65 and not x20 and x21 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x66 and not x65 and not x20 and x21 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x20 and x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x20 and not x21 and x17 and x13 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x66 and not x65 and not x20 and not x21 and x17 and not x13 and x12 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x66 and not x65 and not x20 and not x21 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s17 =>
      if ( x66 and x67 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x67 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x67 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x24 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      else
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s150;

      end if;

   when s18 =>
      if ( x63 and x62 ) = '1' then
         y34 <= '1' ;
         current_group15m <= s21;

      elsif ( x63 and not x62 and x15 and x8 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x63 and not x62 and x15 and not x8 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x63 and not x62 and not x15 and x16 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( x63 and not x62 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s135;

      else
         y34 <= '1' ;
         current_group15m <= s21;

      end if;

   when s19 =>
      if ( x66 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( not x66 and x26 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      else
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      end if;

   when s20 =>
      if ( x64 ) = '1' then
         current_group15m <= s1;

      elsif ( not x64 and x63 and x18 and x15 and x8 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x64 and x63 and x18 and x15 and not x8 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x64 and x63 and x18 and not x15 and x16 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( not x64 and x63 and x18 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s135;

      elsif ( not x64 and x63 and not x18 ) = '1' then
         y31 <= '1' ;
         current_group15m <= s96;

      else
         y15 <= '1' ;
         current_group15m <= s149;

      end if;

   when s21 =>
      if ( x63 ) = '1' then
         y35 <= '1' ;
         current_group15m <= s26;

      elsif ( not x63 and x62 ) = '1' then
         y35 <= '1' ;
         current_group15m <= s26;

      elsif ( not x63 and not x62 and x64 and x16 and x8 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x63 and not x62 and x64 and x16 and not x8 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x63 and not x62 and x64 and not x16 and x4 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( not x63 and not x62 and x64 and not x16 and not x4 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s135;

      elsif ( not x63 and not x62 and not x64 and x15 and x8 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x63 and not x62 and not x64 and x15 and not x8 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x63 and not x62 and not x64 and not x15 and x16 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s151;

      elsif ( not x63 and not x62 and not x64 and not x15 and not x16 and x14 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s135;

      else
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s152;

      end if;

   when s22 =>
      if ( x65 and x21 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( x65 and not x21 and x22 and x23 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x21 and x22 and not x23 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and not x21 and not x22 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x67 and x64 and x63 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and x67 and x64 and not x63 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and not x64 and x63 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x67 and not x64 and not x63 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( not x65 and not x67 and x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and x23 and x22 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and not x67 and not x21 and x23 and x22 and x17 and not x14 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and not x67 and not x21 and x23 and x22 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and x23 and x22 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and x23 and not x22 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s23 =>
      if ( x65 and x16 and x11 and x12 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s153;

      elsif ( x65 and x16 and x11 and not x12 and x13 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s153;

      elsif ( x65 and x16 and x11 and not x12 and not x13 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s154;

      elsif ( x65 and x16 and not x11 and x13 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s63;

      elsif ( x65 and x16 and not x11 and not x13 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( x65 and not x16 and x17 and x11 and x13 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x65 and not x16 and x17 and x11 and not x13 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( x65 and not x16 and x17 and not x11 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x65 and not x16 and not x17 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( not x65 and x66 and x62 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and x66 and not x62 and x63 and x64 and x17 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and x66 and not x62 and x63 and x64 and x17 and not x13 and x12 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and x66 and not x62 and x63 and x64 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x62 and x63 and x64 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x62 and x63 and not x64 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s156;

      elsif ( not x65 and x66 and not x62 and not x63 and x64 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s152;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and x15 and x14 and x8 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and x15 and x14 and not x8 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and x15 and not x14 and x7 and x8 ) = '1' then
         y24 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s157;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and x15 and not x14 and x7 and not x8 ) = '1' then
         y26 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s158;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and x15 and not x14 and not x7 and x8 and x12 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s65;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and x15 and not x14 and not x7 and x8 and not x12 and x19 and x13 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and x15 and not x14 and not x7 and x8 and not x12 and x19 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and x15 and not x14 and not x7 and x8 and not x12 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and x15 and not x14 and not x7 and not x8 and x13 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s65;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and x15 and not x14 and not x7 and not x8 and not x13 and x19 and x12 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and x15 and not x14 and not x7 and not x8 and not x13 and x19 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and x15 and not x14 and not x7 and not x8 and not x13 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and x8 and x7 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and x8 and x7 and not x3 and x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and x8 and x7 and not x3 and not x4 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and x8 and not x7 and x9 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and x8 and not x7 and x9 and not x3 and x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and x8 and not x7 and x9 and not x3 and not x4 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and x8 and not x7 and not x9 and x3 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and x8 and not x7 and not x9 and not x3 and x19 and x13 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and x8 and not x7 and not x9 and not x3 and x19 and not x13 and x12 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and x8 and not x7 and not x9 and not x3 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and x8 and not x7 and not x9 and not x3 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and not x8 and x7 and x11 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and not x8 and x7 and x11 and not x3 and x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and not x8 and x7 and x11 and not x3 and not x4 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and not x8 and x7 and not x11 and x3 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and not x8 and x7 and not x11 and not x3 and x19 and x13 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and not x8 and x7 and not x11 and not x3 and x19 and not x13 and x12 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and not x8 and x7 and not x11 and not x3 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and not x8 and x7 and not x11 and not x3 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and not x8 and not x7 and x10 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and not x8 and not x7 and x10 and not x3 and x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and not x8 and not x7 and x10 and not x3 and not x4 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and not x8 and not x7 and not x10 and x3 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and not x8 and not x7 and not x10 and not x3 and x19 and x13 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and not x8 and not x7 and not x10 and not x3 and x19 and not x13 and x12 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and not x8 and not x7 and not x10 and not x3 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and x16 and not x15 and not x8 and not x7 and not x10 and not x3 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and not x16 and x15 and x7 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s159;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and not x16 and x15 and not x7 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and not x16 and x15 and not x7 and not x3 and x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and not x16 and x15 and not x7 and not x3 and not x4 and x8 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and not x16 and x15 and not x7 and not x3 and not x4 and not x8 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and not x16 and not x15 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and not x16 and not x15 and not x3 and x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and not x16 and not x15 and not x3 and not x4 and x14 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s135;

      elsif ( not x65 and x66 and not x62 and not x63 and not x64 and not x16 and not x15 and not x3 and not x4 and not x14 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s156;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and x26 and x17 and x11 and x13 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s160;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and x26 and x17 and x11 and not x13 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and x26 and x17 and not x11 and x12 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and x26 and x17 and not x11 and x12 and not x13 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s48;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and x26 and x17 and not x11 and not x12 and x13 and x14 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s161;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and x26 and x17 and not x11 and not x12 and x13 and not x14 and x18 and x15 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and x26 and x17 and not x11 and not x12 and x13 and not x14 and x18 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and x26 and x17 and not x11 and not x12 and x13 and not x14 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and x26 and x17 and not x11 and not x12 and not x13 and x15 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s161;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and x26 and x17 and not x11 and not x12 and not x13 and not x15 and x18 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and x26 and x17 and not x11 and not x12 and not x13 and not x15 and x18 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and x26 and x17 and not x11 and not x12 and not x13 and not x15 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and x26 and not x17 and x13 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and x26 and not x17 and not x13 and x12 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and x26 and not x17 and not x13 and not x12 and x2 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and x26 and not x17 and not x13 and not x12 and not x2 and x11 and x4 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s50;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and x26 and not x17 and not x13 and not x12 and not x2 and x11 and not x4 ) = '1' then
         y8 <= '1' ;
         y17 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s164;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and x26 and not x17 and not x13 and not x12 and not x2 and not x11 and x4 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and x26 and not x17 and not x13 and not x12 and not x2 and not x11 and not x4 ) = '1' then
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s165;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and x17 and x11 and x13 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and x17 and x11 and not x13 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and x17 and not x11 and x12 and x13 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and x17 and not x11 and x12 and not x13 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and x17 and not x11 and not x12 and x13 and x14 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s167;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and x17 and not x11 and not x12 and x13 and not x14 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and x17 and not x11 and not x12 and x13 and not x14 and x20 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and x17 and not x11 and not x12 and x13 and not x14 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and x17 and not x11 and not x12 and not x13 and x15 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s167;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and x17 and not x11 and not x12 and not x13 and not x15 and x20 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and x17 and not x11 and not x12 and not x13 and not x15 and x20 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and x17 and not x11 and not x12 and not x13 and not x15 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and not x17 and x11 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and not x17 and x11 and not x3 and x12 and x4 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and not x17 and x11 and not x3 and x12 and not x4 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s169;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and not x17 and x11 and not x3 and not x12 and x13 and x4 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and not x17 and x11 and not x3 and not x12 and x13 and not x4 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s170;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and not x17 and x11 and not x3 and not x12 and not x13 and x4 ) = '1' then
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s165;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and not x17 and x11 and not x3 and not x12 and not x13 and not x4 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and not x17 and not x11 and x13 and x12 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s51;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and not x17 and not x11 and x13 and not x12 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s170;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and not x17 and not x11 and not x13 and x12 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and not x17 and not x11 and not x13 and not x12 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and not x17 and not x11 and not x13 and not x12 and not x3 and x4 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x66 and x67 and x24 and x16 and not x26 and not x17 and not x11 and not x13 and not x12 and not x3 and not x4 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s171;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and x13 and x11 and x9 and x18 and x15 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and x13 and x11 and x9 and x18 and not x15 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and x13 and x11 and x9 and x18 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and x13 and x11 and x9 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and x13 and x11 and not x9 and x2 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and x13 and x11 and not x9 and not x2 and x4 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and x13 and x11 and not x9 and not x2 and not x4 ) = '1' then
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s165;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and x13 and not x11 and x12 and x2 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and x13 and not x11 and x12 and not x2 and x4 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and x13 and not x11 and x12 and not x2 and not x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and x13 and not x11 and not x12 and x8 and x2 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and x13 and not x11 and not x12 and x8 and not x2 and x4 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and x13 and not x11 and not x12 and x8 and not x2 and not x4 ) = '1' then
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s165;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and x13 and not x11 and not x12 and not x8 and x18 and x15 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and x13 and not x11 and not x12 and not x8 and x18 and not x15 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and x13 and not x11 and not x12 and not x8 and x18 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and x13 and not x11 and not x12 and not x8 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and not x13 and x11 and x2 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and not x13 and x11 and not x2 and x4 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s172;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and not x13 and x11 and not x2 and not x4 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and not x13 and not x11 and x12 and x10 and x2 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and not x13 and not x11 and x12 and x10 and not x2 and x4 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and not x13 and not x11 and x12 and x10 and not x2 and not x4 ) = '1' then
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s165;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and not x13 and not x11 and x12 and not x10 and x18 and x15 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and not x13 and not x11 and x12 and not x10 and x18 and not x15 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and not x13 and not x11 and x12 and not x10 and x18 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and not x13 and not x11 and x12 and not x10 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and not x13 and not x11 and not x12 and x9 and x2 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and not x13 and not x11 and not x12 and x9 and not x2 and x4 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and not x13 and not x11 and not x12 and x9 and not x2 and not x4 ) = '1' then
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s165;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and not x13 and not x11 and not x12 and not x9 and x18 and x15 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and not x13 and not x11 and not x12 and not x9 and x18 and not x15 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and not x13 and not x11 and not x12 and not x9 and x18 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and x17 and not x13 and not x11 and not x12 and not x9 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and not x17 and x2 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and not x17 and not x2 and x4 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and x26 and not x17 and not x2 and not x4 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and x13 and x11 and x9 and x4 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and x13 and x11 and x9 and not x4 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and x13 and x11 and not x9 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and x13 and x11 and not x9 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and x13 and x11 and not x9 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and x13 and x11 and not x9 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and x13 and not x11 and x12 and x4 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and x13 and not x11 and x12 and not x4 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and x13 and not x11 and not x12 and x7 and x4 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and x13 and not x11 and not x12 and x7 and not x4 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and x13 and not x11 and not x12 and not x7 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and x13 and not x11 and not x12 and not x7 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and x13 and not x11 and not x12 and not x7 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and x13 and not x11 and not x12 and not x7 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and not x13 and x11 and x4 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s173;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and not x13 and x11 and not x4 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and not x13 and not x11 and x12 and x10 and x4 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and not x13 and not x11 and x12 and x10 and not x4 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and not x13 and not x11 and x12 and not x10 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and not x13 and not x11 and x12 and not x10 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and not x13 and not x11 and x12 and not x10 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and not x13 and not x11 and x12 and not x10 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and not x13 and not x11 and not x12 and x8 and x4 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and not x13 and not x11 and not x12 and x8 and not x4 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and not x13 and not x11 and not x12 and not x8 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and not x13 and not x11 and not x12 and not x8 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and not x13 and not x11 and not x12 and not x8 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and x17 and not x13 and not x11 and not x12 and not x8 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and not x17 and x4 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x66 and x67 and x24 and not x16 and not x26 and not x3 and not x17 and not x4 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s174;

      elsif ( not x65 and not x66 and x67 and not x24 and x25 and x26 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x66 and x67 and not x24 and x25 and not x26 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and x67 and not x24 and x25 and not x26 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and x67 and not x24 and x25 and not x26 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and not x24 and x25 and not x26 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and not x24 and not x25 and x26 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x65 and not x66 and x67 and not x24 and not x25 and x26 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x65 and not x66 and x67 and not x24 and not x25 and x26 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and not x24 and not x25 and not x26 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and x68 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x66 and not x67 and not x68 and x21 and x10 and x11 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( not x65 and not x66 and not x67 and not x68 and x21 and x10 and not x11 ) = '1' then
         current_group15m <= s23;

      elsif ( not x65 and not x66 and not x67 and not x68 and x21 and not x10 ) = '1' then
         y10 <= '1' ;
         y17 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s104;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and x8 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s176;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and not x8 and x10 and x19 and x15 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s177;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and not x8 and x10 and x19 and not x15 ) = '1' then
         y2 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and not x8 and x10 and not x19 and x20 and x15 and x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s178;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and not x8 and x10 and not x19 and x20 and x15 and not x14 and x16 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s178;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and not x8 and x10 and not x19 and x20 and x15 and not x14 and not x16 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and not x8 and x10 and not x19 and x20 and x15 and not x14 and not x16 and x5 and not x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and not x8 and x10 and not x19 and x20 and x15 and not x14 and not x16 and x5 and not x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and not x8 and x10 and not x19 and x20 and x15 and not x14 and not x16 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and not x8 and x10 and not x19 and x20 and not x15 and x14 and x18 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s178;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and not x8 and x10 and not x19 and x20 and not x15 and x14 and not x18 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and not x8 and x10 and not x19 and x20 and not x15 and x14 and not x18 and x5 and not x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and not x8 and x10 and not x19 and x20 and not x15 and x14 and not x18 and x5 and not x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and not x8 and x10 and not x19 and x20 and not x15 and x14 and not x18 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and not x8 and x10 and not x19 and x20 and not x15 and not x14 and x17 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s178;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and not x8 and x10 and not x19 and x20 and not x15 and not x14 and not x17 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and not x8 and x10 and not x19 and x20 and not x15 and not x14 and not x17 and x5 and not x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and not x8 and x10 and not x19 and x20 and not x15 and not x14 and not x17 and x5 and not x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and not x8 and x10 and not x19 and x20 and not x15 and not x14 and not x17 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and not x8 and x10 and not x19 and not x20 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s151;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x22 and not x8 and not x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and not x22 and x10 and x19 and x15 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and not x22 and x10 and x19 and not x15 ) = '1' then
         y2 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and not x22 and x10 and not x19 and x20 ) = '1' then
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s179;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and not x22 and x10 and not x19 and not x20 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s151;

      else
         y10 <= '1' ;
         y17 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s104;

      end if;

   when s24 =>
      if ( x65 and x21 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x21 and x22 and x23 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( x65 and not x21 and x22 and not x23 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x65 and not x21 and not x22 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x66 and x67 and x64 and x63 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and x66 and x67 and x64 and not x63 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x64 and x63 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x66 and x67 and not x64 and not x63 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( not x65 and x66 and not x67 and x21 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s180;

      elsif ( not x65 and x66 and not x67 and not x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x24 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and x16 and x10 and x26 and x12 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and x16 and x10 and x26 and not x12 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and x16 and x10 and not x26 and x12 ) = '1' then
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s165;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and x16 and x10 and not x26 and not x12 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and x16 and not x10 and x11 and x26 and x12 ) = '1' then
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s165;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and x16 and not x10 and x11 and x26 and not x12 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and x16 and not x10 and x11 and not x26 and x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and x16 and not x10 and x11 and not x26 and not x12 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s160;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and x16 and not x10 and not x11 and x12 and x13 and x26 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and x16 and not x10 and not x11 and x12 and x13 and not x26 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s181;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and x16 and not x10 and not x11 and x12 and not x13 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and x16 and not x10 and not x11 and x12 and not x13 and x19 and not x14 and x26 ) = '1' then
         current_group15m <= s24;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and x16 and not x10 and not x11 and x12 and not x13 and x19 and not x14 and not x26 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and x16 and not x10 and not x11 and x12 and not x13 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and x16 and not x10 and not x11 and not x12 and x14 and x26 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and x16 and not x10 and not x11 and not x12 and x14 and not x26 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s181;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and x16 and not x10 and not x11 and not x12 and not x14 and x19 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and x16 and not x10 and not x11 and not x12 and not x14 and x19 and not x13 and x26 ) = '1' then
         current_group15m <= s24;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and x16 and not x10 and not x11 and not x12 and not x14 and x19 and not x13 and not x26 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and x16 and not x10 and not x11 and not x12 and not x14 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and x26 and x10 and x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and x26 and x10 and not x3 and x1 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and x26 and x10 and not x3 and not x1 and x11 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s171;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and x26 and x10 and not x3 and not x1 and not x11 and x12 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s183;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and x26 and x10 and not x3 and not x1 and not x11 and not x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and x26 and not x10 and x11 and x12 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and x26 and not x10 and x11 and not x12 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s172;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and x26 and not x10 and not x11 and x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and x26 and not x10 and not x11 and not x3 and x12 and x1 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and x26 and not x10 and not x11 and not x3 and x12 and not x1 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s184;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and x26 and not x10 and not x11 and not x3 and not x12 and x1 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s185;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and x26 and not x10 and not x11 and not x3 and not x12 and not x1 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and not x26 and x10 and x5 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s186;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and not x26 and x10 and not x5 and x2 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s174;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and not x26 and x10 and not x5 and not x2 and x11 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s187;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and not x26 and x10 and not x5 and not x2 and not x11 and x12 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s187;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and not x26 and x10 and not x5 and not x2 and not x11 and not x12 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s171;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and not x26 and not x10 and x11 and x12 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and not x26 and not x10 and x11 and not x12 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s187;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and not x26 and not x10 and not x11 and x5 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s186;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and not x26 and not x10 and not x11 and not x5 and x2 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s174;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and not x26 and not x10 and not x11 and not x5 and not x2 and x12 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s187;

      elsif ( not x65 and not x66 and not x24 and x25 and x15 and not x16 and not x26 and not x10 and not x11 and not x5 and not x2 and not x12 ) = '1' then
         y12 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s49;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and x16 and x10 and x12 and x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and x16 and x10 and x12 and not x8 and x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and x16 and x10 and x12 and not x8 and not x3 and x1 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and x16 and x10 and x12 and not x8 and not x3 and not x1 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and x16 and x10 and not x12 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and x16 and not x10 and x12 and x7 and x11 and x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and x16 and not x10 and x12 and x7 and x11 and not x3 and x1 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and x16 and not x10 and x12 and x7 and x11 and not x3 and not x1 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and x16 and not x10 and x12 and x7 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and x16 and not x10 and x12 and not x7 and x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and x16 and not x10 and x12 and not x7 and not x3 and x1 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and x16 and not x10 and x12 and not x7 and not x3 and not x1 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and x16 and not x10 and not x12 and x11 and x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and x16 and not x10 and not x12 and x11 and not x9 and x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and x16 and not x10 and not x12 and x11 and not x9 and not x3 and x1 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and x16 and not x10 and not x12 and x11 and not x9 and not x3 and not x1 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and x16 and not x10 and not x12 and not x11 and x8 and x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and x16 and not x10 and not x12 and not x11 and x8 and not x3 and x1 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and x16 and not x10 and not x12 and not x11 and x8 and not x3 and not x1 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and x16 and not x10 and not x12 and not x11 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and not x16 and x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and not x16 and not x3 and x1 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and x26 and not x16 and not x3 and not x1 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s188;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and x5 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s186;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and x12 and x10 and x8 and x2 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s174;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and x12 and x10 and x8 and not x2 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and x12 and x10 and not x8 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and x12 and x10 and not x8 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and x12 and x10 and not x8 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and x12 and x10 and not x8 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and x12 and not x10 and x11 and x2 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s174;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and x12 and not x10 and x11 and not x2 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and x12 and not x10 and not x11 and x7 and x2 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s174;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and x12 and not x10 and not x11 and x7 and not x2 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and x12 and not x10 and not x11 and not x7 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and x12 and not x10 and not x11 and not x7 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and x12 and not x10 and not x11 and not x7 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and x12 and not x10 and not x11 and not x7 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and not x12 and x10 and x2 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s51;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and not x12 and x10 and not x2 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s174;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and not x12 and not x10 and x11 and x9 and x2 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s174;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and not x12 and not x10 and x11 and x9 and not x2 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and not x12 and not x10 and x11 and not x9 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and not x12 and not x10 and x11 and not x9 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and not x12 and not x10 and x11 and not x9 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and not x12 and not x10 and x11 and not x9 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and not x12 and not x10 and not x11 and x8 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and not x12 and not x10 and not x11 and x8 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and not x12 and not x10 and not x11 and x8 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and not x12 and not x10 and not x11 and x8 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and not x12 and not x10 and not x11 and not x8 and x2 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s174;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and x16 and not x12 and not x10 and not x11 and not x8 and not x2 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and not x16 and x2 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s174;

      elsif ( not x65 and not x66 and not x24 and x25 and not x15 and not x26 and not x5 and not x16 and not x2 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s19;

      elsif ( not x65 and not x66 and not x24 and not x25 and x26 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s189;

      else
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s190;

      end if;

   when s25 =>
      if ( x66 and x65 and x15 and x16 and x12 and x10 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x66 and x65 and x15 and x16 and x12 and not x10 and x20 and x13 and x11 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s126;

      elsif ( x66 and x65 and x15 and x16 and x12 and not x10 and x20 and x13 and not x11 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s191;

      elsif ( x66 and x65 and x15 and x16 and x12 and not x10 and x20 and not x13 and x19 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and x65 and x15 and x16 and x12 and not x10 and x20 and not x13 and x19 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and x15 and x16 and x12 and not x10 and x20 and not x13 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and x15 and x16 and x12 and not x10 and not x20 and x21 and x11 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s126;

      elsif ( x66 and x65 and x15 and x16 and x12 and not x10 and not x20 and x21 and not x11 and x13 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s125;

      elsif ( x66 and x65 and x15 and x16 and x12 and not x10 and not x20 and x21 and not x11 and not x13 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and x15 and x16 and x12 and not x10 and not x20 and x21 and not x11 and not x13 and x19 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and x15 and x16 and x12 and not x10 and not x20 and x21 and not x11 and not x13 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and x15 and x16 and x12 and not x10 and not x20 and not x21 and x13 and x11 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s126;

      elsif ( x66 and x65 and x15 and x16 and x12 and not x10 and not x20 and not x21 and x13 and not x11 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s191;

      elsif ( x66 and x65 and x15 and x16 and x12 and not x10 and not x20 and not x21 and not x13 and x19 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and x65 and x15 and x16 and x12 and not x10 and not x20 and not x21 and not x13 and x19 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and x15 and x16 and x12 and not x10 and not x20 and not x21 and not x13 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and x15 and x16 and not x12 and x10 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( x66 and x65 and x15 and x16 and not x12 and not x10 and x11 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s192;

      elsif ( x66 and x65 and x15 and x16 and not x12 and not x10 and not x11 and x14 and x20 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s191;

      elsif ( x66 and x65 and x15 and x16 and not x12 and not x10 and not x11 and x14 and not x20 and x21 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s125;

      elsif ( x66 and x65 and x15 and x16 and not x12 and not x10 and not x11 and x14 and not x20 and not x21 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s191;

      elsif ( x66 and x65 and x15 and x16 and not x12 and not x10 and not x11 and not x14 and x19 and x13 and x20 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and x65 and x15 and x16 and not x12 and not x10 and not x11 and not x14 and x19 and x13 and not x20 and x21 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and x15 and x16 and not x12 and not x10 and not x11 and not x14 and x19 and x13 and not x20 and not x21 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and x65 and x15 and x16 and not x12 and not x10 and not x11 and not x14 and x19 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and x15 and x16 and not x12 and not x10 and not x11 and not x14 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and x15 and not x16 and x10 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x66 and x65 and x15 and not x16 and x10 and not x2 and x20 and x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x66 and x65 and x15 and not x16 and x10 and not x2 and x20 and not x4 and x11 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x66 and x65 and x15 and not x16 and x10 and not x2 and x20 and not x4 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s193;

      elsif ( x66 and x65 and x15 and not x16 and x10 and not x2 and x20 and not x4 and not x11 and not x12 ) = '1' then
         y1 <= '1' ;
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s194;

      elsif ( x66 and x65 and x15 and not x16 and x10 and not x2 and not x20 and x21 and x3 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( x66 and x65 and x15 and not x16 and x10 and not x2 and not x20 and x21 and not x3 and x11 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x66 and x65 and x15 and not x16 and x10 and not x2 and not x20 and x21 and not x3 and not x11 and x12 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s193;

      elsif ( x66 and x65 and x15 and not x16 and x10 and not x2 and not x20 and x21 and not x3 and not x11 and not x12 ) = '1' then
         y8 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s195;

      elsif ( x66 and x65 and x15 and not x16 and x10 and not x2 and not x20 and not x21 and x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x66 and x65 and x15 and not x16 and x10 and not x2 and not x20 and not x21 and not x4 and x11 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x66 and x65 and x15 and not x16 and x10 and not x2 and not x20 and not x21 and not x4 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s193;

      elsif ( x66 and x65 and x15 and not x16 and x10 and not x2 and not x20 and not x21 and not x4 and not x11 and not x12 ) = '1' then
         y1 <= '1' ;
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s194;

      elsif ( x66 and x65 and x15 and not x16 and not x10 and x11 and x20 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x66 and x65 and x15 and not x16 and not x10 and x11 and not x20 and x21 and x12 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and x65 and x15 and not x16 and not x10 and x11 and not x20 and x21 and not x12 ) = '1' then
         y1 <= '1' ;
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s194;

      elsif ( x66 and x65 and x15 and not x16 and not x10 and x11 and not x20 and not x21 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x66 and x65 and x15 and not x16 and not x10 and not x11 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x66 and x65 and x15 and not x16 and not x10 and not x11 and not x2 and x20 and x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x66 and x65 and x15 and not x16 and not x10 and not x11 and not x2 and x20 and not x4 and x12 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s196;

      elsif ( x66 and x65 and x15 and not x16 and not x10 and not x11 and not x2 and x20 and not x4 and not x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s192;

      elsif ( x66 and x65 and x15 and not x16 and not x10 and not x11 and not x2 and not x20 and x21 and x3 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( x66 and x65 and x15 and not x16 and not x10 and not x11 and not x2 and not x20 and x21 and not x3 and x12 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      elsif ( x66 and x65 and x15 and not x16 and not x10 and not x11 and not x2 and not x20 and x21 and not x3 and not x12 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s198;

      elsif ( x66 and x65 and x15 and not x16 and not x10 and not x11 and not x2 and not x20 and not x21 and x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x66 and x65 and x15 and not x16 and not x10 and not x11 and not x2 and not x20 and not x21 and not x4 and x12 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s196;

      elsif ( x66 and x65 and x15 and not x16 and not x10 and not x11 and not x2 and not x20 and not x21 and not x4 and not x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s192;

      elsif ( x66 and x65 and not x15 and x20 and x16 and x10 and x12 and x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x15 and x20 and x16 and x10 and x12 and not x8 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x66 and x65 and not x15 and x20 and x16 and x10 and x12 and not x8 and not x2 and x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x66 and x65 and not x15 and x20 and x16 and x10 and x12 and not x8 and not x2 and not x4 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s199;

      elsif ( x66 and x65 and not x15 and x20 and x16 and x10 and not x12 and x9 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x66 and x65 and not x15 and x20 and x16 and x10 and not x12 and x9 and not x2 and x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s200;

      elsif ( x66 and x65 and not x15 and x20 and x16 and x10 and not x12 and x9 and not x2 and not x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x66 and x65 and not x15 and x20 and x16 and x10 and not x12 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x15 and x20 and x16 and not x10 and x12 and x7 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x66 and x65 and not x15 and x20 and x16 and not x10 and x12 and x7 and not x2 and x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x66 and x65 and not x15 and x20 and x16 and not x10 and x12 and x7 and not x2 and not x4 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s199;

      elsif ( x66 and x65 and not x15 and x20 and x16 and not x10 and x12 and not x7 and x11 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x66 and x65 and not x15 and x20 and x16 and not x10 and x12 and not x7 and x11 and not x2 and x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x66 and x65 and not x15 and x20 and x16 and not x10 and x12 and not x7 and x11 and not x2 and not x4 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s199;

      elsif ( x66 and x65 and not x15 and x20 and x16 and not x10 and x12 and not x7 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x15 and x20 and x16 and not x10 and not x12 and x11 and x9 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x66 and x65 and not x15 and x20 and x16 and not x10 and not x12 and x11 and x9 and not x2 and x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x66 and x65 and not x15 and x20 and x16 and not x10 and not x12 and x11 and x9 and not x2 and not x4 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s199;

      elsif ( x66 and x65 and not x15 and x20 and x16 and not x10 and not x12 and x11 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x15 and x20 and x16 and not x10 and not x12 and not x11 and x8 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x66 and x65 and not x15 and x20 and x16 and not x10 and not x12 and not x11 and x8 and not x2 and x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x66 and x65 and not x15 and x20 and x16 and not x10 and not x12 and not x11 and x8 and not x2 and not x4 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s199;

      elsif ( x66 and x65 and not x15 and x20 and x16 and not x10 and not x12 and not x11 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x15 and x20 and not x16 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x66 and x65 and not x15 and x20 and not x16 and not x2 and x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x66 and x65 and not x15 and x20 and not x16 and not x2 and not x4 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s201;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and x10 and x8 and x3 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s202;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and x10 and x8 and not x3 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and x10 and not x8 and x12 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and x10 and not x8 and x12 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and x10 and not x8 and x12 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and x10 and not x8 and x12 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and x10 and not x8 and not x12 and x3 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s202;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and x10 and not x8 and not x12 and not x3 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and not x10 and x12 and x11 and x3 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and not x10 and x12 and x11 and not x3 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s192;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and not x10 and x12 and not x11 and x7 and x3 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s202;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and not x10 and x12 and not x11 and x7 and not x3 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and not x10 and x12 and not x11 and not x7 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and not x10 and x12 and not x11 and not x7 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and not x10 and x12 and not x11 and not x7 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and not x10 and x12 and not x11 and not x7 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and not x10 and not x12 and x11 and x9 and x3 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s202;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and not x10 and not x12 and x11 and x9 and not x3 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and not x10 and not x12 and x11 and not x9 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and not x10 and not x12 and x11 and not x9 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and not x10 and not x12 and x11 and not x9 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and not x10 and not x12 and x11 and not x9 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and not x10 and not x12 and not x11 and x8 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and not x10 and not x12 and not x11 and x8 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and not x10 and not x12 and not x11 and x8 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and not x10 and not x12 and not x11 and x8 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and not x10 and not x12 and not x11 and not x8 and x3 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s202;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and x16 and not x10 and not x12 and not x11 and not x8 and not x3 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and not x16 and x3 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( x66 and x65 and not x15 and not x20 and x21 and not x2 and not x16 and not x3 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and x10 and x12 and x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and x10 and x12 and not x8 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and x10 and x12 and not x8 and not x2 and x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and x10 and x12 and not x8 and not x2 and not x4 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s199;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and x10 and not x12 and x9 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and x10 and not x12 and x9 and not x2 and x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s200;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and x10 and not x12 and x9 and not x2 and not x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and x10 and not x12 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and not x10 and x12 and x7 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and not x10 and x12 and x7 and not x2 and x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and not x10 and x12 and x7 and not x2 and not x4 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s199;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and not x10 and x12 and not x7 and x11 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and not x10 and x12 and not x7 and x11 and not x2 and x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and not x10 and x12 and not x7 and x11 and not x2 and not x4 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s199;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and not x10 and x12 and not x7 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and not x10 and not x12 and x11 and x9 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and not x10 and not x12 and x11 and x9 and not x2 and x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and not x10 and not x12 and x11 and x9 and not x2 and not x4 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s199;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and not x10 and not x12 and x11 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and not x10 and not x12 and not x11 and x8 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and not x10 and not x12 and not x11 and x8 and not x2 and x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and not x10 and not x12 and not x11 and x8 and not x2 and not x4 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s199;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and x16 and not x10 and not x12 and not x11 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and not x16 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and not x16 and not x2 and x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x66 and x65 and not x15 and not x20 and not x21 and not x16 and not x2 and not x4 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s201;

      elsif ( x66 and not x65 and x62 and x16 and x15 and x14 and x9 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and not x65 and x62 and x16 and x15 and x14 and not x9 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and not x65 and x62 and x16 and x15 and not x14 and x7 and x9 ) = '1' then
         y24 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s157;

      elsif ( x66 and not x65 and x62 and x16 and x15 and not x14 and x7 and not x9 ) = '1' then
         y26 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s158;

      elsif ( x66 and not x65 and x62 and x16 and x15 and not x14 and not x7 and x9 and x12 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s65;

      elsif ( x66 and not x65 and x62 and x16 and x15 and not x14 and not x7 and x9 and not x12 and x61 and x13 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x66 and not x65 and x62 and x16 and x15 and not x14 and not x7 and x9 and not x12 and x61 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and x62 and x16 and x15 and not x14 and not x7 and x9 and not x12 and not x61 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and x62 and x16 and x15 and not x14 and not x7 and not x9 and x13 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s65;

      elsif ( x66 and not x65 and x62 and x16 and x15 and not x14 and not x7 and not x9 and not x13 and x61 and x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x66 and not x65 and x62 and x16 and x15 and not x14 and not x7 and not x9 and not x13 and x61 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and x62 and x16 and x15 and not x14 and not x7 and not x9 and not x13 and not x61 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and x62 and x16 and not x15 and x9 and x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( x66 and not x65 and x62 and x16 and not x15 and x9 and not x3 and x4 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x66 and not x65 and x62 and x16 and not x15 and x9 and not x3 and not x4 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( x66 and not x65 and x62 and x16 and not x15 and not x9 and x7 and x11 and x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( x66 and not x65 and x62 and x16 and not x15 and not x9 and x7 and x11 and not x3 and x4 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x66 and not x65 and x62 and x16 and not x15 and not x9 and x7 and x11 and not x3 and not x4 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( x66 and not x65 and x62 and x16 and not x15 and not x9 and x7 and not x11 and x3 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x66 and not x65 and x62 and x16 and not x15 and not x9 and x7 and not x11 and not x3 and x61 and x13 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x66 and not x65 and x62 and x16 and not x15 and not x9 and x7 and not x11 and not x3 and x61 and not x13 and x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x66 and not x65 and x62 and x16 and not x15 and not x9 and x7 and not x11 and not x3 and x61 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and x62 and x16 and not x15 and not x9 and x7 and not x11 and not x3 and not x61 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and x62 and x16 and not x15 and not x9 and not x7 and x10 and x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( x66 and not x65 and x62 and x16 and not x15 and not x9 and not x7 and x10 and not x3 and x4 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x66 and not x65 and x62 and x16 and not x15 and not x9 and not x7 and x10 and not x3 and not x4 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( x66 and not x65 and x62 and x16 and not x15 and not x9 and not x7 and not x10 and x3 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x66 and not x65 and x62 and x16 and not x15 and not x9 and not x7 and not x10 and not x3 and x61 and x13 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x66 and not x65 and x62 and x16 and not x15 and not x9 and not x7 and not x10 and not x3 and x61 and not x13 and x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x66 and not x65 and x62 and x16 and not x15 and not x9 and not x7 and not x10 and not x3 and x61 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and x62 and x16 and not x15 and not x9 and not x7 and not x10 and not x3 and not x61 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and x62 and not x16 and x15 and x7 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( x66 and not x65 and x62 and not x16 and x15 and not x7 and x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( x66 and not x65 and x62 and not x16 and x15 and not x7 and not x3 and x4 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x66 and not x65 and x62 and not x16 and x15 and not x7 and not x3 and not x4 and x8 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x66 and not x65 and x62 and not x16 and x15 and not x7 and not x3 and not x4 and not x8 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( x66 and not x65 and x62 and not x16 and not x15 and x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( x66 and not x65 and x62 and not x16 and not x15 and not x3 and x4 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x66 and not x65 and x62 and not x16 and not x15 and not x3 and not x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( x66 and not x65 and not x62 and x63 and x64 and x17 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and not x65 and not x62 and x63 and x64 and x17 and not x13 and x12 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and not x65 and not x62 and x63 and x64 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x62 and x63 and x64 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x62 and x63 and not x64 and x15 and x8 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x66 and not x65 and not x62 and x63 and not x64 and x15 and not x8 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x66 and not x65 and not x62 and x63 and not x64 and not x15 and x16 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x66 and not x65 and not x62 and x63 and not x64 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s135;

      elsif ( x66 and not x65 and not x62 and not x63 and x64 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x66 and not x65 and not x62 and not x63 and not x64 and x6 and x15 and x8 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and not x65 and not x62 and not x63 and not x64 and x6 and x15 and not x8 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s203;

      elsif ( x66 and not x65 and not x62 and not x63 and not x64 and x6 and not x15 and x16 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and not x65 and not x62 and not x63 and not x64 and x6 and not x15 and not x16 and x14 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s204;

      elsif ( x66 and not x65 and not x62 and not x63 and not x64 and x6 and not x15 and not x16 and not x14 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s20;

      elsif ( x66 and not x65 and not x62 and not x63 and not x64 and not x6 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x66 and x65 and x21 and x15 and x9 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x66 and x65 and x21 and x15 and not x9 and x6 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x66 and x65 and x21 and x15 and not x9 and not x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x66 and x65 and x21 and not x15 and x16 and x9 and x8 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x66 and x65 and x21 and not x15 and x16 and x9 and not x8 and x10 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x66 and x65 and x21 and not x15 and x16 and x9 and not x8 and not x10 and x18 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x66 and x65 and x21 and not x15 and x16 and x9 and not x8 and not x10 and not x18 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and x21 and not x15 and x16 and x9 and not x8 and not x10 and not x18 and x19 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and x21 and not x15 and x16 and x9 and not x8 and not x10 and not x18 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and x21 and not x15 and x16 and x9 and not x8 and not x10 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and x21 and not x15 and x16 and not x9 and x8 and x12 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x66 and x65 and x21 and not x15 and x16 and not x9 and x8 and not x12 and x18 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x66 and x65 and x21 and not x15 and x16 and not x9 and x8 and not x12 and not x18 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and x21 and not x15 and x16 and not x9 and x8 and not x12 and not x18 and x19 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and x21 and not x15 and x16 and not x9 and x8 and not x12 and not x18 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and x21 and not x15 and x16 and not x9 and x8 and not x12 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and x21 and not x15 and x16 and not x9 and not x8 and x11 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x66 and x65 and x21 and not x15 and x16 and not x9 and not x8 and not x11 and x18 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x66 and x65 and x21 and not x15 and x16 and not x9 and not x8 and not x11 and not x18 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and x21 and not x15 and x16 and not x9 and not x8 and not x11 and not x18 and x19 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and x21 and not x15 and x16 and not x9 and not x8 and not x11 and not x18 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and x21 and not x15 and x16 and not x9 and not x8 and not x11 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and x21 and not x15 and not x16 and x6 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s205;

      elsif ( not x66 and x65 and x21 and not x15 and not x16 and not x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x66 and x65 and not x21 and x22 and x18 and x14 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( not x66 and x65 and not x21 and x22 and x18 and not x14 and x13 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( not x66 and x65 and not x21 and x22 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and x22 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and x23 and x15 and x9 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and x65 and not x21 and not x22 and x23 and x15 and not x9 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x66 and x65 and not x21 and not x22 and x23 and not x15 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s205;

      elsif ( not x66 and x65 and not x21 and not x22 and not x23 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and not x65 and x68 and x20 and x15 and x8 ) = '1' then
         y2 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s206;

      elsif ( not x66 and not x65 and x68 and x20 and x15 and not x8 and x6 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s207;

      elsif ( not x66 and not x65 and x68 and x20 and x15 and not x8 and not x6 ) = '1' then
         y2 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s208;

      elsif ( not x66 and not x65 and x68 and x20 and not x15 and x16 and x7 and x8 ) = '1' then
         y2 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s208;

      elsif ( not x66 and not x65 and x68 and x20 and not x15 and x16 and x7 and not x8 ) = '1' then
         y2 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s206;

      elsif ( not x66 and not x65 and x68 and x20 and not x15 and x16 and not x7 ) = '1' then
         y2 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s206;

      elsif ( not x66 and not x65 and x68 and x20 and not x15 and not x16 and x6 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s209;

      elsif ( not x66 and not x65 and x68 and x20 and not x15 and not x16 and not x6 ) = '1' then
         y2 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s208;

      elsif ( not x66 and not x65 and x68 and not x20 and x21 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and x15 and x14 and x8 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and x15 and x14 and not x8 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s126;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and x15 and not x14 and x7 and x8 ) = '1' then
         y1 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y13 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s207;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and x15 and not x14 and x7 and not x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s210;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and x15 and not x14 and not x7 and x8 and x12 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and x15 and not x14 and not x7 and x8 and not x12 and x17 and x13 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and x15 and not x14 and not x7 and x8 and not x12 and x17 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and x15 and not x14 and not x7 and x8 and not x12 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and x15 and not x14 and not x7 and not x8 and x13 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and x15 and not x14 and not x7 and not x8 and not x13 and x17 and x12 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and x15 and not x14 and not x7 and not x8 and not x13 and x17 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and x15 and not x14 and not x7 and not x8 and not x13 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and x8 and x7 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and x8 and x7 and not x2 and x3 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and x8 and x7 and not x2 and not x3 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and x8 and not x7 and x9 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and x8 and not x7 and x9 and not x2 and x3 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and x8 and not x7 and x9 and not x2 and not x3 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and x8 and not x7 and not x9 and x2 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and x8 and not x7 and not x9 and not x2 and x17 and x13 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and x8 and not x7 and not x9 and not x2 and x17 and not x13 and x12 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and x8 and not x7 and not x9 and not x2 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and x8 and not x7 and not x9 and not x2 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and not x8 and x7 and x11 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and not x8 and x7 and x11 and not x2 and x3 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and not x8 and x7 and x11 and not x2 and not x3 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and not x8 and x7 and not x11 and x2 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and not x8 and x7 and not x11 and not x2 and x17 and x13 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and not x8 and x7 and not x11 and not x2 and x17 and not x13 and x12 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and not x8 and x7 and not x11 and not x2 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and not x8 and x7 and not x11 and not x2 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and not x8 and not x7 and x10 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and not x8 and not x7 and x10 and not x2 and x3 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and not x8 and not x7 and x10 and not x2 and not x3 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and not x8 and not x7 and not x10 and x2 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and not x8 and not x7 and not x10 and not x2 and x17 and x13 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and not x8 and not x7 and not x10 and not x2 and x17 and not x13 and x12 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and not x8 and not x7 and not x10 and not x2 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and x16 and not x15 and not x8 and not x7 and not x10 and not x2 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and not x16 and x15 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and not x16 and x15 and not x7 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and not x16 and x15 and not x7 and not x2 and x3 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and not x16 and x15 and not x7 and not x2 and not x3 and x8 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s41;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and not x16 and x15 and not x7 and not x2 and not x3 and not x8 ) = '1' then
         y2 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s206;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and not x16 and not x15 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and not x16 and not x15 and not x2 and x3 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x66 and not x65 and x68 and not x20 and not x21 and not x16 and not x15 and not x2 and not x3 ) = '1' then
         y7 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s211;

      elsif ( not x66 and not x65 and not x68 and x24 and x26 and x11 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s160;

      elsif ( not x66 and not x65 and not x68 and x24 and x26 and not x11 and x18 and x15 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x66 and not x65 and not x68 and x24 and x26 and not x11 and x18 and not x15 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x66 and not x65 and not x68 and x24 and x26 and not x11 and x18 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x68 and x24 and x26 and not x11 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x68 and x24 and not x26 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x66 and not x65 and not x68 and x24 and not x26 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x66 and not x65 and not x68 and x24 and not x26 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x68 and x24 and not x26 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x68 and not x24 and x25 and x26 and x15 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x68 and not x24 and x25 and x26 and not x15 and x3 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( not x66 and not x65 and not x68 and not x24 and x25 and x26 and not x15 and not x3 and x1 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x66 and not x65 and not x68 and not x24 and x25 and x26 and not x15 and not x3 and not x1 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and not x65 and not x68 and not x24 and x25 and not x26 and x18 and x15 and x10 and x11 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s187;

      elsif ( not x66 and not x65 and not x68 and not x24 and x25 and not x26 and x18 and x15 and x10 and not x11 and x12 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s185;

      elsif ( not x66 and not x65 and not x68 and not x24 and x25 and not x26 and x18 and x15 and x10 and not x11 and not x12 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s160;

      elsif ( not x66 and not x65 and not x68 and not x24 and x25 and not x26 and x18 and x15 and not x10 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s50;

      elsif ( not x66 and not x65 and not x68 and not x24 and x25 and not x26 and x18 and not x15 and x16 and x10 and x12 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( not x66 and not x65 and not x68 and not x24 and x25 and not x26 and x18 and not x15 and x16 and x10 and not x12 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x66 and not x65 and not x68 and not x24 and x25 and not x26 and x18 and not x15 and x16 and not x10 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( not x66 and not x65 and not x68 and not x24 and x25 and not x26 and x18 and not x15 and not x16 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x66 and not x65 and not x68 and not x24 and x25 and not x26 and not x18 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x66 and not x65 and not x68 and not x24 and not x25 and x26 and x10 and x12 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and not x65 and not x68 and not x24 and not x25 and x26 and x10 and x12 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and not x65 and not x68 and not x24 and not x25 and x26 and x10 and x12 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x68 and not x24 and not x25 and x26 and x10 and x12 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x68 and not x24 and not x25 and x26 and x10 and not x12 ) = '1' then
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s165;

      elsif ( not x66 and not x65 and not x68 and not x24 and not x25 and x26 and not x10 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and not x65 and not x68 and not x24 and not x25 and x26 and not x10 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and not x65 and not x68 and not x24 and not x25 and x26 and not x10 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x68 and not x24 and not x25 and x26 and not x10 and not x18 ) = '1' then
         current_group15m <= s1;

      else
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      end if;

   when s26 =>
      if ( x65 and x21 and x15 and x9 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( x65 and x21 and x15 and not x9 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( x65 and x21 and not x15 and x16 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x65 and x21 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s212;

      elsif ( x65 and not x21 and x23 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x23 and x22 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x21 and not x23 and not x22 and x17 and x15 and x9 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( x65 and not x21 and not x23 and not x22 and x17 and x15 and not x9 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( x65 and not x21 and not x23 and not x22 and x17 and not x15 and x16 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( x65 and not x21 and not x23 and not x22 and x17 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s205;

      elsif ( x65 and not x21 and not x23 and not x22 and not x17 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( not x65 and x62 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( not x65 and not x62 and x63 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s213;

      else
         current_group15m <= s1;

      end if;

   when s27 =>
      if ( x66 and x65 and x67 and x22 and x17 and x18 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and x65 and x67 and x22 and x17 and not x18 and x19 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and x65 and x67 and x22 and x17 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and x67 and x22 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and x67 and not x22 and x18 and x13 and x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x66 and x65 and x67 and not x22 and x18 and x13 and not x23 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and x67 and not x22 and x18 and not x13 and x12 and x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x66 and x65 and x67 and not x22 and x18 and not x13 and x12 and not x23 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and x67 and not x22 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and x67 and not x22 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x67 and x21 and x20 and x12 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and x65 and not x67 and x21 and x20 and x12 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and x65 and not x67 and x21 and x20 and x12 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x67 and x21 and x20 and x12 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x67 and x21 and x20 and not x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x67 and not x21 and x12 and x19 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and x65 and not x67 and not x21 and x12 and x19 and not x14 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and x65 and not x67 and not x21 and x12 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x67 and not x21 and x12 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x67 and not x21 and not x12 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x66 and not x65 and x67 and x62 and x15 and x8 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( x66 and not x65 and x67 and x62 and x15 and not x8 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x66 and not x65 and x67 and x62 and not x15 and x16 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x66 and not x65 and x67 and x62 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s135;

      elsif ( x66 and not x65 and x67 and not x62 and x63 and x6 and x15 and x8 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and not x65 and x67 and not x62 and x63 and x6 and x15 and not x8 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s203;

      elsif ( x66 and not x65 and x67 and not x62 and x63 and x6 and not x15 and x16 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and not x65 and x67 and not x62 and x63 and x6 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s204;

      elsif ( x66 and not x65 and x67 and not x62 and x63 and not x6 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and not x65 and x67 and not x62 and not x63 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and x21 and x16 and x15 and x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s214;

      elsif ( x66 and not x65 and not x67 and x21 and x16 and x15 and not x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s215;

      elsif ( x66 and not x65 and not x67 and x21 and x16 and not x15 and x10 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x66 and not x65 and not x67 and x21 and x16 and not x15 and not x10 ) = '1' then
         y14 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s216;

      elsif ( x66 and not x65 and not x67 and x21 and not x16 and x17 and x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s215;

      elsif ( x66 and not x65 and not x67 and x21 and not x16 and x17 and not x10 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s217;

      elsif ( x66 and not x65 and not x67 and x21 and not x16 and not x17 and x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s215;

      elsif ( x66 and not x65 and not x67 and x21 and not x16 and not x17 and not x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s218;

      elsif ( x66 and not x65 and not x67 and not x21 and x10 and x22 and x4 and x17 and x15 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s219;

      elsif ( x66 and not x65 and not x67 and not x21 and x10 and x22 and x4 and x17 and not x15 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x66 and not x65 and not x67 and not x21 and x10 and x22 and x4 and not x17 and x18 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s219;

      elsif ( x66 and not x65 and not x67 and not x21 and x10 and x22 and x4 and not x17 and not x18 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s219;

      elsif ( x66 and not x65 and not x67 and not x21 and x10 and x22 and not x4 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x66 and not x65 and not x67 and not x21 and x10 and not x22 and x7 and x16 and x15 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s219;

      elsif ( x66 and not x65 and not x67 and not x21 and x10 and not x22 and x7 and x16 and not x15 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s220;

      elsif ( x66 and not x65 and not x67 and not x21 and x10 and not x22 and x7 and not x16 and x17 and x15 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s219;

      elsif ( x66 and not x65 and not x67 and not x21 and x10 and not x22 and x7 and not x16 and x17 and not x15 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s220;

      elsif ( x66 and not x65 and not x67 and not x21 and x10 and not x22 and x7 and not x16 and not x17 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s219;

      elsif ( x66 and not x65 and not x67 and not x21 and x10 and not x22 and not x7 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s220;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and x17 and x4 and x15 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s219;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and x17 and x4 and not x15 ) = '1' then
         y2 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s221;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and x17 and not x4 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and not x17 and x18 and x15 and x12 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and not x17 and x18 and x15 and not x12 and x14 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and not x17 and x18 and x15 and not x12 and not x14 and x7 and x8 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and not x17 and x18 and x15 and not x12 and not x14 and x7 and not x8 and x9 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and not x17 and x18 and x15 and not x12 and not x14 and x7 and not x8 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and not x17 and x18 and x15 and not x12 and not x14 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and not x17 and x18 and not x15 and x14 and x13 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and not x17 and x18 and not x15 and x14 and not x13 and x7 and x8 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and not x17 and x18 and not x15 and x14 and not x13 and x7 and not x8 and x9 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and not x17 and x18 and not x15 and x14 and not x13 and x7 and not x8 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and not x17 and x18 and not x15 and x14 and not x13 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and not x17 and x18 and not x15 and not x14 and x11 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and not x17 and x18 and not x15 and not x14 and not x11 and x7 and x8 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and not x17 and x18 and not x15 and not x14 and not x11 and x7 and not x8 and x9 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and not x17 and x18 and not x15 and not x14 and not x11 and x7 and not x8 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and not x17 and x18 and not x15 and not x14 and not x11 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and not x17 and not x18 and x4 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s220;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and x22 and not x17 and not x18 and not x4 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and x16 and x7 and x15 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s222;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and x16 and x7 and not x15 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and x16 and not x7 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s220;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and not x16 and x17 and x14 and x13 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s220;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and not x16 and x17 and x14 and not x13 and x15 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s220;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and not x16 and x17 and x14 and not x13 and not x15 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and not x16 and x17 and x14 and not x13 and not x15 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and not x16 and x17 and x14 and not x13 and not x15 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and not x16 and x17 and x14 and not x13 and not x15 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and not x16 and x17 and not x14 and x15 and x12 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s220;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and not x16 and x17 and not x14 and x15 and not x12 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and not x16 and x17 and not x14 and x15 and not x12 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and not x16 and x17 and not x14 and x15 and not x12 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and not x16 and x17 and not x14 and x15 and not x12 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and not x16 and x17 and not x14 and not x15 and x11 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s220;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and not x16 and x17 and not x14 and not x15 and not x11 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and not x16 and x17 and not x14 and not x15 and not x11 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and not x16 and x17 and not x14 and not x15 and not x11 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and not x16 and x17 and not x14 and not x15 and not x11 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and not x16 and not x17 and x7 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( x66 and not x65 and not x67 and not x21 and not x10 and not x22 and not x16 and not x17 and not x7 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s220;

      elsif ( not x66 and x65 and x21 and x67 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and x21 and not x67 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and x21 and not x67 and x19 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and x21 and not x67 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and x21 and not x67 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and x22 and x67 and x23 and x18 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x66 and x65 and not x21 and x22 and x67 and x23 and not x18 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x66 and x65 and not x21 and x22 and x67 and x23 and not x18 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x66 and x65 and not x21 and x22 and x67 and x23 and not x18 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and x22 and x67 and x23 and not x18 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and x22 and x67 and not x23 ) = '1' then
         y6 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s223;

      elsif ( not x66 and x65 and not x21 and x22 and not x67 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( not x66 and x65 and not x21 and x22 and not x67 and not x19 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( not x66 and x65 and not x21 and x22 and not x67 and not x19 and x17 and not x14 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( not x66 and x65 and not x21 and x22 and not x67 and not x19 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and x22 and not x67 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and x67 and x23 ) = '1' then
         y6 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s223;

      elsif ( not x66 and x65 and not x21 and not x22 and x67 and not x23 and x19 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x66 and x65 and not x21 and not x22 and x67 and not x23 and not x19 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x66 and x65 and not x21 and not x22 and x67 and not x23 and not x19 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x66 and x65 and not x21 and not x22 and x67 and not x23 and not x19 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and x67 and not x23 and not x19 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and x7 and x23 and x9 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and x7 and x23 and not x9 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and x7 and not x23 and x9 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and x7 and not x23 and not x9 ) = '1' then
         y24 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s157;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and not x7 and x8 and x23 and x9 ) = '1' then
         y24 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s157;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and not x7 and x8 and x23 and not x9 ) = '1' then
         y26 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s158;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and not x7 and x8 and not x23 and x9 ) = '1' then
         y26 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s158;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and not x7 and x8 and not x23 and not x9 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s212;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and not x7 and not x8 and x23 and x13 and x9 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s191;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and not x7 and not x8 and x23 and x13 and not x9 and x14 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s191;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and not x7 and not x8 and x23 and x13 and not x9 and not x14 and x20 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and not x7 and not x8 and x23 and x13 and not x9 and not x14 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and not x7 and not x8 and x23 and not x13 and x14 and x9 and x20 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and not x7 and not x8 and x23 and not x13 and x14 and x9 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and not x7 and not x8 and x23 and not x13 and x14 and not x9 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s191;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and not x7 and not x8 and x23 and not x13 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and not x7 and not x8 and not x23 and x13 and x9 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s224;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and not x7 and not x8 and not x23 and x13 and not x9 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s224;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and not x7 and not x8 and not x23 and x13 and not x9 and not x14 and x18 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and not x7 and not x8 and not x23 and x13 and not x9 and not x14 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and not x7 and not x8 and not x23 and not x13 and x14 and x9 and x18 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and not x7 and not x8 and not x23 and not x13 and x14 and x9 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and not x7 and not x8 and not x23 and not x13 and x14 and not x9 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s224;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and x16 and not x7 and not x8 and not x23 and not x13 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and not x16 and x7 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and not x16 and not x7 and x8 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and not x16 and not x7 and not x8 and x5 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s22;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and not x16 and not x7 and not x8 and not x5 and x2 and x23 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and not x16 and not x7 and not x8 and not x5 and x2 and not x23 and x9 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and not x16 and not x7 and not x8 and not x5 and x2 and not x23 and not x9 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and not x16 and not x7 and not x8 and not x5 and not x2 and x9 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and not x16 and not x7 and not x8 and not x5 and not x2 and not x9 and x23 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and x15 and not x16 and not x7 and not x8 and not x5 and not x2 and not x9 and not x23 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and x5 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s22;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and x23 and x16 and x9 and x10 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and x23 and x16 and x9 and not x10 and x8 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and x23 and x16 and x9 and not x10 and not x8 and x20 and x14 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and x23 and x16 and x9 and not x10 and not x8 and x20 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and x23 and x16 and x9 and not x10 and not x8 and x20 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and x23 and x16 and x9 and not x10 and not x8 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and x23 and x16 and not x9 and x8 and x12 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and x23 and x16 and not x9 and x8 and not x12 and x20 and x14 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and x23 and x16 and not x9 and x8 and not x12 and x20 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and x23 and x16 and not x9 and x8 and not x12 and x20 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and x23 and x16 and not x9 and x8 and not x12 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and x23 and x16 and not x9 and not x8 and x11 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and x23 and x16 and not x9 and not x8 and not x11 and x20 and x14 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and x23 and x16 and not x9 and not x8 and not x11 and x20 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and x23 and x16 and not x9 and not x8 and not x11 and x20 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and x23 and x16 and not x9 and not x8 and not x11 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and x23 and not x16 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and x23 and not x16 and not x2 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s212;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and not x23 and x16 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and not x23 and x16 and x9 and not x10 and x8 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and not x23 and x16 and x9 and not x10 and not x8 and x18 and x14 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and not x23 and x16 and x9 and not x10 and not x8 and x18 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and not x23 and x16 and x9 and not x10 and not x8 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and not x23 and x16 and x9 and not x10 and not x8 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and not x23 and x16 and not x9 and x8 and x12 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and not x23 and x16 and not x9 and x8 and not x12 and x18 and x14 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and not x23 and x16 and not x9 and x8 and not x12 and x18 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and not x23 and x16 and not x9 and x8 and not x12 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and not x23 and x16 and not x9 and x8 and not x12 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and not x23 and x16 and not x9 and not x8 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and not x23 and x16 and not x9 and not x8 and not x11 and x18 and x14 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and not x23 and x16 and not x9 and not x8 and not x11 and x18 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and not x23 and x16 and not x9 and not x8 and not x11 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and not x23 and x16 and not x9 and not x8 and not x11 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and not x23 and not x16 and x2 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x66 and x65 and not x21 and not x22 and not x67 and not x15 and not x5 and not x23 and not x16 and not x2 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s205;

      elsif ( not x66 and not x65 and x67 and x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and not x20 and x21 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x66 and not x65 and x67 and not x20 and x21 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x66 and not x65 and x67 and not x20 and x21 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and not x20 and x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and not x20 and not x21 and x17 and x13 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x66 and not x65 and x67 and not x20 and not x21 and x17 and not x13 and x12 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x66 and not x65 and x67 and not x20 and not x21 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and not x20 and not x21 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x67 and x21 and x9 and x3 ) = '1' then
         current_group15m <= s40;

      elsif ( not x66 and not x65 and not x67 and x21 and x9 and not x3 and x4 ) = '1' then
         current_group15m <= s40;

      elsif ( not x66 and not x65 and not x67 and x21 and x9 and not x3 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x67 and x21 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and x12 and x19 and x15 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and x12 and x19 and not x15 ) = '1' then
         y2 <= '1' ;
         y11 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s123;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and x12 and not x19 and x20 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and x12 and not x19 and not x20 ) = '1' then
         y6 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s225;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( not x66 and not x65 and not x67 and not x21 and not x22 and x4 and x5 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and not x65 and not x67 and not x21 and not x22 and x4 and not x5 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and not x65 and not x67 and not x21 and not x22 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s28 =>
      if ( x21 and x65 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x65 and x16 and x6 and x15 and x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s214;

      elsif ( x21 and not x65 and x16 and x6 and x15 and not x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s215;

      elsif ( x21 and not x65 and x16 and x6 and not x15 and x10 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x21 and not x65 and x16 and x6 and not x15 and not x10 ) = '1' then
         y14 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s216;

      elsif ( x21 and not x65 and x16 and not x6 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s220;

      elsif ( x21 and not x65 and not x16 and x17 and x10 and x6 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s215;

      elsif ( x21 and not x65 and not x16 and x17 and x10 and not x6 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s220;

      elsif ( x21 and not x65 and not x16 and x17 and not x10 and x6 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x21 and not x65 and not x16 and x17 and not x10 and not x6 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s226;

      elsif ( x21 and not x65 and not x16 and not x17 and x6 and x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s215;

      elsif ( x21 and not x65 and not x16 and not x17 and x6 and not x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s218;

      elsif ( x21 and not x65 and not x16 and not x17 and not x6 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s220;

      elsif ( not x21 and x22 and x65 and x23 and x5 and x18 and x15 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( not x21 and x22 and x65 and x23 and x5 and x18 and not x15 ) = '1' then
         y15 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s227;

      elsif ( not x21 and x22 and x65 and x23 and x5 and not x18 and x19 and x15 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s228;

      elsif ( not x21 and x22 and x65 and x23 and x5 and not x18 and x19 and not x15 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( not x21 and x22 and x65 and x23 and x5 and not x18 and not x19 ) = '1' then
         y15 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s36;

      elsif ( not x21 and x22 and x65 and x23 and not x5 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( not x21 and x22 and x65 and not x23 ) = '1' then
         y12 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s230;

      elsif ( not x21 and x22 and not x65 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x21 and not x22 and x65 and x23 and x19 and x6 and x16 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( not x21 and not x22 and x65 and x23 and x19 and x6 and not x16 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x21 and not x22 and x65 and x23 and x19 and not x6 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( not x21 and not x22 and x65 and x23 and not x19 and x20 and x16 and x6 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s228;

      elsif ( not x21 and not x22 and x65 and x23 and not x19 and x20 and x16 and not x6 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( not x21 and not x22 and x65 and x23 and not x19 and x20 and not x16 and x17 and x18 and x6 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x21 and not x22 and x65 and x23 and not x19 and x20 and not x16 and x17 and x18 and not x6 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( not x21 and not x22 and x65 and x23 and not x19 and x20 and not x16 and x17 and not x18 and x14 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x21 and not x22 and x65 and x23 and not x19 and x20 and not x16 and x17 and not x18 and not x14 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( not x21 and not x22 and x65 and x23 and not x19 and x20 and not x16 and not x17 and x18 and x14 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x21 and not x22 and x65 and x23 and not x19 and x20 and not x16 and not x17 and x18 and not x14 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( not x21 and not x22 and x65 and x23 and not x19 and x20 and not x16 and not x17 and not x18 and x6 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x21 and not x22 and x65 and x23 and not x19 and x20 and not x16 and not x17 and not x18 and not x6 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( not x21 and not x22 and x65 and x23 and not x19 and not x20 and x6 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s231;

      elsif ( not x21 and not x22 and x65 and x23 and not x19 and not x20 and not x6 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( not x21 and not x22 and x65 and not x23 and x5 and x18 and x15 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( not x21 and not x22 and x65 and not x23 and x5 and x18 and not x15 ) = '1' then
         y15 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s227;

      elsif ( not x21 and not x22 and x65 and not x23 and x5 and not x18 and x19 and x15 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s228;

      elsif ( not x21 and not x22 and x65 and not x23 and x5 and not x18 and x19 and not x15 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( not x21 and not x22 and x65 and not x23 and x5 and not x18 and not x19 ) = '1' then
         y15 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s36;

      elsif ( not x21 and not x22 and x65 and not x23 and not x5 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      else
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s232;

      end if;

   when s29 =>
      if ( x65 and x21 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x22 and x23 and x18 and x19 and x15 and x17 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and not x21 and x22 and x23 and x18 and x19 and x15 and not x17 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x21 and x22 and x23 and x18 and x19 and not x15 and x16 and x17 ) = '1' then
         y24 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s157;

      elsif ( x65 and not x21 and x22 and x23 and x18 and x19 and not x15 and x16 and not x17 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         y20 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s227;

      elsif ( x65 and not x21 and x22 and x23 and x18 and x19 and not x15 and not x16 and x8 and x10 and x17 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and x22 and x23 and x18 and x19 and not x15 and not x16 and x8 and x10 and not x17 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x65 and not x21 and x22 and x23 and x18 and x19 and not x15 and not x16 and x8 and not x10 and x11 and x17 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x65 and not x21 and x22 and x23 and x18 and x19 and not x15 and not x16 and x8 and not x10 and x11 and not x17 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and x22 and x23 and x18 and x19 and not x15 and not x16 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x22 and x23 and x18 and x19 and not x15 and not x16 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x22 and x23 and x18 and not x19 and x16 and x15 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s203;

      elsif ( x65 and not x21 and x22 and x23 and x18 and not x19 and x16 and not x15 and x17 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x65 and not x21 and x22 and x23 and x18 and not x19 and x16 and not x15 and not x17 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s233;

      elsif ( x65 and not x21 and x22 and x23 and x18 and not x19 and not x16 and x17 and x15 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s234;

      elsif ( x65 and not x21 and x22 and x23 and x18 and not x19 and not x16 and x17 and not x15 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s235;

      elsif ( x65 and not x21 and x22 and x23 and x18 and not x19 and not x16 and not x17 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s236;

      elsif ( x65 and not x21 and x22 and x23 and x18 and not x19 and not x16 and not x17 and not x4 and x6 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x65 and not x21 and x22 and x23 and x18 and not x19 and not x16 and not x17 and not x4 and not x6 and x15 ) = '1' then
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s227;

      elsif ( x65 and not x21 and x22 and x23 and x18 and not x19 and not x16 and not x17 and not x4 and not x6 and not x15 ) = '1' then
         y16 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s227;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and x19 and x15 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s236;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and x19 and x15 and not x4 and x6 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and x19 and x15 and not x4 and not x6 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s117;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and x19 and not x15 and x17 and x13 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s236;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and x19 and not x15 and x17 and x13 and not x4 and x6 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and x19 and not x15 and x17 and x13 and not x4 and not x6 ) = '1' then
         y8 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s227;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and x19 and not x15 and x17 and not x13 and x16 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s236;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and x19 and not x15 and x17 and not x13 and x16 and not x4 and x6 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and x19 and not x15 and x17 and not x13 and x16 and not x4 and not x6 ) = '1' then
         y8 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s227;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and x19 and not x15 and x17 and not x13 and not x16 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and x19 and not x15 and not x17 and x16 and x14 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s236;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and x19 and not x15 and not x17 and x16 and x14 and not x4 and x6 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and x19 and not x15 and not x17 and x16 and x14 and not x4 and not x6 ) = '1' then
         y8 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s227;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and x19 and not x15 and not x17 and x16 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and x19 and not x15 and not x17 and not x16 and x12 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s236;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and x19 and not x15 and not x17 and not x16 and x12 and not x4 and x6 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and x19 and not x15 and not x17 and not x16 and x12 and not x4 and not x6 ) = '1' then
         y8 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s227;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and x19 and not x15 and not x17 and not x16 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and not x19 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s236;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and not x19 and not x4 and x6 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x65 and not x21 and x22 and x23 and not x18 and not x19 and not x4 and not x6 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x65 and not x21 and x22 and not x23 and x15 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      elsif ( x65 and not x21 and x22 and not x23 and not x15 and x19 and x18 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      elsif ( x65 and not x21 and x22 and not x23 and not x15 and x19 and not x18 and x8 and x9 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and x22 and not x23 and not x15 and x19 and not x18 and x8 and not x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and x22 and not x23 and not x15 and x19 and not x18 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x22 and not x23 and not x15 and x19 and not x18 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x22 and not x23 and not x15 and not x19 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      elsif ( x65 and not x21 and not x22 and x23 and x5 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s28;

      elsif ( x65 and not x21 and not x22 and x23 and not x5 and x19 and x6 and x16 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( x65 and not x21 and not x22 and x23 and not x5 and x19 and x6 and not x16 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x65 and not x21 and not x22 and x23 and not x5 and x19 and not x6 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( x65 and not x21 and not x22 and x23 and not x5 and not x19 and x20 and x16 and x6 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s228;

      elsif ( x65 and not x21 and not x22 and x23 and not x5 and not x19 and x20 and x16 and not x6 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( x65 and not x21 and not x22 and x23 and not x5 and not x19 and x20 and not x16 and x17 and x18 and x6 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( x65 and not x21 and not x22 and x23 and not x5 and not x19 and x20 and not x16 and x17 and x18 and not x6 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( x65 and not x21 and not x22 and x23 and not x5 and not x19 and x20 and not x16 and x17 and not x18 and x14 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( x65 and not x21 and not x22 and x23 and not x5 and not x19 and x20 and not x16 and x17 and not x18 and not x14 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( x65 and not x21 and not x22 and x23 and not x5 and not x19 and x20 and not x16 and not x17 and x18 and x14 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( x65 and not x21 and not x22 and x23 and not x5 and not x19 and x20 and not x16 and not x17 and x18 and not x14 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( x65 and not x21 and not x22 and x23 and not x5 and not x19 and x20 and not x16 and not x17 and not x18 and x6 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( x65 and not x21 and not x22 and x23 and not x5 and not x19 and x20 and not x16 and not x17 and not x18 and not x6 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( x65 and not x21 and not x22 and x23 and not x5 and not x19 and not x20 and x6 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s231;

      elsif ( x65 and not x21 and not x22 and x23 and not x5 and not x19 and not x20 and not x6 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and x19 and x15 and x17 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and x19 and x15 and not x17 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and x19 and not x15 and x16 and x17 ) = '1' then
         y24 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s157;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and x19 and not x15 and x16 and not x17 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         y20 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s227;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and x19 and not x15 and not x16 and x8 and x10 and x17 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and x19 and not x15 and not x16 and x8 and x10 and not x17 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and x19 and not x15 and not x16 and x8 and not x10 and x11 and x17 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and x19 and not x15 and not x16 and x8 and not x10 and x11 and not x17 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and x19 and not x15 and not x16 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and x19 and not x15 and not x16 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and not x19 and x16 and x15 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s203;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and not x19 and x16 and not x15 and x17 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and not x19 and x16 and not x15 and not x17 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s233;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and not x19 and not x16 and x17 and x15 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s234;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and not x19 and not x16 and x17 and not x15 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s235;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and not x19 and not x16 and not x17 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s236;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and not x19 and not x16 and not x17 and not x4 and x6 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and not x19 and not x16 and not x17 and not x4 and not x6 and x15 ) = '1' then
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s227;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and not x19 and not x16 and not x17 and not x4 and not x6 and not x15 ) = '1' then
         y16 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s227;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and x19 and x15 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s236;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and x19 and x15 and not x4 and x6 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and x19 and x15 and not x4 and not x6 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s117;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and x19 and not x15 and x17 and x13 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s236;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and x19 and not x15 and x17 and x13 and not x4 and x6 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and x19 and not x15 and x17 and x13 and not x4 and not x6 ) = '1' then
         y8 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s227;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and x19 and not x15 and x17 and not x13 and x16 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s236;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and x19 and not x15 and x17 and not x13 and x16 and not x4 and x6 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and x19 and not x15 and x17 and not x13 and x16 and not x4 and not x6 ) = '1' then
         y8 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s227;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and x19 and not x15 and x17 and not x13 and not x16 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and x19 and not x15 and not x17 and x16 and x14 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s236;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and x19 and not x15 and not x17 and x16 and x14 and not x4 and x6 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and x19 and not x15 and not x17 and x16 and x14 and not x4 and not x6 ) = '1' then
         y8 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s227;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and x19 and not x15 and not x17 and x16 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and x19 and not x15 and not x17 and not x16 and x12 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s236;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and x19 and not x15 and not x17 and not x16 and x12 and not x4 and x6 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and x19 and not x15 and not x17 and not x16 and x12 and not x4 and not x6 ) = '1' then
         y8 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s227;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and x19 and not x15 and not x17 and not x16 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and not x19 and x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s236;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and not x19 and not x4 and x6 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 and not x19 and not x4 and not x6 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( not x65 and x66 and x21 and x4 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s28;

      elsif ( not x65 and x66 and x21 and not x4 and x16 and x6 and x15 and x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s214;

      elsif ( not x65 and x66 and x21 and not x4 and x16 and x6 and x15 and not x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s215;

      elsif ( not x65 and x66 and x21 and not x4 and x16 and x6 and not x15 and x10 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and x66 and x21 and not x4 and x16 and x6 and not x15 and not x10 ) = '1' then
         y14 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s216;

      elsif ( not x65 and x66 and x21 and not x4 and x16 and not x6 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s220;

      elsif ( not x65 and x66 and x21 and not x4 and not x16 and x17 and x10 and x6 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s215;

      elsif ( not x65 and x66 and x21 and not x4 and not x16 and x17 and x10 and not x6 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s220;

      elsif ( not x65 and x66 and x21 and not x4 and not x16 and x17 and not x10 and x6 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( not x65 and x66 and x21 and not x4 and not x16 and x17 and not x10 and not x6 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s226;

      elsif ( not x65 and x66 and x21 and not x4 and not x16 and not x17 and x6 and x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s215;

      elsif ( not x65 and x66 and x21 and not x4 and not x16 and not x17 and x6 and not x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s218;

      elsif ( not x65 and x66 and x21 and not x4 and not x16 and not x17 and not x6 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s220;

      elsif ( not x65 and x66 and not x21 and x22 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s218;

      elsif ( not x65 and x66 and not x21 and not x22 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x24 and x26 and x16 and x18 and x15 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and not x66 and x24 and x26 and x16 and x18 and not x15 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and not x66 and x24 and x26 and x16 and x18 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x24 and x26 and x16 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x24 and x26 and not x16 ) = '1' then
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s165;

      elsif ( not x65 and not x66 and x24 and not x26 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and not x66 and x24 and not x26 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and not x66 and x24 and not x26 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x24 and not x26 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x24 and x25 and x26 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and not x24 and x25 and x26 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and not x24 and x25 and x26 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s29;

      elsif ( not x65 and not x66 and not x24 and x25 and x26 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x24 and x25 and not x26 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( not x65 and not x66 and not x24 and not x25 and x26 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      else
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s239;

      end if;

   when s30 =>
      if ( x65 and x66 and x67 and x22 and x17 and x18 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and x67 and x22 and x17 and not x18 and x19 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and x67 and x22 and x17 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x67 and x22 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x67 and not x22 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and x66 and x67 and not x22 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and x66 and x67 and not x22 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x67 and not x22 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x67 and x60 and x61 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x66 and not x67 and x60 and x61 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x66 and not x67 and x60 and x61 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x66 and not x67 and x60 and x61 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x66 and not x67 and x60 and not x61 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and not x67 and x60 and not x61 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and not x67 and x60 and not x61 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x66 and not x67 and x60 and not x61 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x66 and not x67 and not x60 and x61 and x62 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( x65 and x66 and not x67 and not x60 and x61 and not x62 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and not x67 and not x60 and x61 and not x62 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and not x67 and not x60 and x61 and not x62 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x66 and not x67 and not x60 and x61 and not x62 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and not x66 and x67 and x21 and x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x65 and not x66 and x67 and x21 and x8 and not x9 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x65 and not x66 and x67 and x21 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and x21 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and not x21 and x23 and x22 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( x65 and not x66 and x67 and not x21 and x23 and not x22 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s240;

      elsif ( x65 and not x66 and x67 and not x21 and not x23 and x22 and x3 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s240;

      elsif ( x65 and not x66 and x67 and not x21 and not x23 and x22 and not x3 and x6 and x18 and x15 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( x65 and not x66 and x67 and not x21 and not x23 and x22 and not x3 and x6 and x18 and not x15 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x65 and not x66 and x67 and not x21 and not x23 and x22 and not x3 and x6 and not x18 and x19 and x15 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x65 and not x66 and x67 and not x21 and not x23 and x22 and not x3 and x6 and not x18 and x19 and not x15 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x65 and not x66 and x67 and not x21 and not x23 and x22 and not x3 and x6 and not x18 and not x19 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( x65 and not x66 and x67 and not x21 and not x23 and x22 and not x3 and not x6 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s28;

      elsif ( x65 and not x66 and x67 and not x21 and not x23 and not x22 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( x65 and not x66 and not x67 ) = '1' then
         y6 <= '1' ;
         y8 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s1;

      else
         y6 <= '1' ;
         y21 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s1;

      end if;

   when s31 =>
      if ( x21 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s241;

      elsif ( not x21 and x23 and x22 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x23 and not x22 and x16 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x21 and x23 and not x22 and not x16 and x20 and x19 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x21 and x23 and not x22 and not x16 and x20 and not x19 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x21 and x23 and not x22 and not x16 and not x20 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x21 and not x23 and x22 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      else
         current_group15m <= s1;

      end if;

   when s32 =>
      if ( x21 and x18 and x19 and x15 and x17 ) = '1' then
         y15 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s227;

      elsif ( x21 and x18 and x19 and x15 and not x17 ) = '1' then
         y16 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s227;

      elsif ( x21 and x18 and x19 and not x15 and x16 and x17 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s203;

      elsif ( x21 and x18 and x19 and not x15 and x16 and not x17 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s233;

      elsif ( x21 and x18 and x19 and not x15 and not x16 and x17 and x10 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x21 and x18 and x19 and not x15 and not x16 and x17 and not x10 and x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and x18 and x19 and not x15 and not x16 and x17 and not x10 and x8 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x18 and x19 and not x15 and not x16 and x17 and not x10 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x18 and x19 and not x15 and not x16 and not x17 and x9 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x21 and x18 and x19 and not x15 and not x16 and not x17 and not x9 and x8 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and x18 and x19 and not x15 and not x16 and not x17 and not x9 and x8 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x18 and x19 and not x15 and not x16 and not x17 and not x9 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x18 and not x19 and x16 and x15 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s243;

      elsif ( x21 and x18 and not x19 and x16 and not x15 and x17 and x14 ) = '1' then
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s227;

      elsif ( x21 and x18 and not x19 and x16 and not x15 and x17 and not x14 ) = '1' then
         y12 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s230;

      elsif ( x21 and x18 and not x19 and x16 and not x15 and not x17 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( x21 and x18 and not x19 and not x16 and x17 and x15 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s44;

      elsif ( x21 and x18 and not x19 and not x16 and x17 and x15 and not x3 and x5 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x21 and x18 and not x19 and not x16 and x17 and x15 and not x3 and not x5 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s228;

      elsif ( x21 and x18 and not x19 and not x16 and x17 and not x15 ) = '1' then
         y6 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s223;

      elsif ( x21 and x18 and not x19 and not x16 and not x17 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s44;

      elsif ( x21 and x18 and not x19 and not x16 and not x17 and not x3 and x5 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x21 and x18 and not x19 and not x16 and not x17 and not x3 and not x5 and x15 ) = '1' then
         y2 <= '1' ;
         y6 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s244;

      elsif ( x21 and x18 and not x19 and not x16 and not x17 and not x3 and not x5 and not x15 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s234;

      elsif ( x21 and not x18 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s44;

      elsif ( x21 and not x18 and not x3 and x19 and x15 and x17 and x5 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x21 and not x18 and not x3 and x19 and x15 and x17 and not x5 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s228;

      elsif ( x21 and not x18 and not x3 and x19 and x15 and not x17 and x5 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s245;

      elsif ( x21 and not x18 and not x3 and x19 and x15 and not x17 and not x5 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x21 and not x18 and not x3 and x19 and not x15 and x16 and x17 and x5 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x21 and not x18 and not x3 and x19 and not x15 and x16 and x17 and not x5 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         y20 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s227;

      elsif ( x21 and not x18 and not x3 and x19 and not x15 and x16 and not x17 and x14 and x5 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x21 and not x18 and not x3 and x19 and not x15 and x16 and not x17 and x14 and not x5 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         y20 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s227;

      elsif ( x21 and not x18 and not x3 and x19 and not x15 and x16 and not x17 and not x14 and x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and not x18 and not x3 and x19 and not x15 and x16 and not x17 and not x14 and x8 and not x9 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and not x18 and not x3 and x19 and not x15 and x16 and not x17 and not x14 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 and not x3 and x19 and not x15 and x16 and not x17 and not x14 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 and not x3 and x19 and not x15 and not x16 and x17 and x12 and x5 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x21 and not x18 and not x3 and x19 and not x15 and not x16 and x17 and x12 and not x5 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         y20 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s227;

      elsif ( x21 and not x18 and not x3 and x19 and not x15 and not x16 and x17 and not x12 and x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and not x18 and not x3 and x19 and not x15 and not x16 and x17 and not x12 and x8 and not x9 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and not x18 and not x3 and x19 and not x15 and not x16 and x17 and not x12 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 and not x3 and x19 and not x15 and not x16 and x17 and not x12 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 and not x3 and x19 and not x15 and not x16 and not x17 and x13 and x5 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x21 and not x18 and not x3 and x19 and not x15 and not x16 and not x17 and x13 and not x5 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         y20 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s227;

      elsif ( x21 and not x18 and not x3 and x19 and not x15 and not x16 and not x17 and not x13 and x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and not x18 and not x3 and x19 and not x15 and not x16 and not x17 and not x13 and x8 and not x9 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and not x18 and not x3 and x19 and not x15 and not x16 and not x17 and not x13 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 and not x3 and x19 and not x15 and not x16 and not x17 and not x13 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 and not x3 and not x19 and x5 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( x21 and not x18 and not x3 and not x19 and not x5 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x21 and x22 and x23 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x21 and x22 and not x23 and x15 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x21 and x22 and not x23 and not x15 and x19 and x18 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x21 and x22 and not x23 and not x15 and x19 and not x18 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s189;

      elsif ( not x21 and x22 and not x23 and not x15 and not x19 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x21 and not x22 and x23 and x4 and x19 and x16 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x21 and not x22 and x23 and x4 and x19 and not x16 ) = '1' then
         y15 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s227;

      elsif ( not x21 and not x22 and x23 and x4 and not x19 and x20 and x16 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s117;

      elsif ( not x21 and not x22 and x23 and x4 and not x19 and x20 and not x16 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x21 and not x22 and x23 and x4 and not x19 and not x20 ) = '1' then
         y3 <= '1' ;
         y12 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s34;

      elsif ( not x21 and not x22 and x23 and not x4 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      else
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      end if;

   when s33 =>
      if ( x21 and x18 and x15 and x17 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and x18 and x15 and not x17 ) = '1' then
         y2 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s244;

      elsif ( x21 and x18 and not x15 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x21 and not x18 and x19 and x15 and x17 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x18 and x19 and x15 and not x17 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s246;

      elsif ( x21 and not x18 and x19 and not x15 ) = '1' then
         y8 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s227;

      elsif ( x21 and not x18 and not x19 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s31;

      elsif ( not x21 and x22 and x23 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x23 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x23 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 ) = '1' then
         current_group15m <= s1;

      else
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s161;

      end if;

   when s34 =>
      if ( x21 and x6 and x18 and x15 and x17 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and x6 and x18 and x15 and not x17 ) = '1' then
         y2 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s244;

      elsif ( x21 and x6 and x18 and not x15 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x21 and x6 and not x18 and x19 and x15 and x17 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and x6 and not x18 and x19 and x15 and not x17 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s246;

      elsif ( x21 and x6 and not x18 and x19 and not x15 ) = '1' then
         y8 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s227;

      elsif ( x21 and x6 and not x18 and not x19 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s31;

      elsif ( x21 and not x6 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s247;

      elsif ( not x21 and x23 and x22 and x18 and x15 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( not x21 and x23 and x22 and x18 and not x15 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x21 and x23 and x22 and not x18 and x19 and x15 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s247;

      elsif ( not x21 and x23 and x22 and not x18 and x19 and not x15 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      elsif ( not x21 and x23 and x22 and not x18 and not x19 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s33;

      elsif ( not x21 and x23 and not x22 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s161;

      elsif ( not x21 and not x23 and x22 ) = '1' then
         current_group15m <= s1;

      else
         y12 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s230;

      end if;

   when s35 =>
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

   when s36 =>
      if ( x21 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s240;

      elsif ( not x21 and x22 and x23 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x23 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x23 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 and x18 and x15 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( not x21 and x22 and not x23 and x18 and not x15 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x21 and x22 and not x23 and not x18 and x19 and x15 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x21 and x22 and not x23 and not x18 and x19 and not x15 ) = '1' then
         y8 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s227;

      elsif ( not x21 and x22 and not x23 and not x18 and not x19 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( not x21 and not x22 and x23 ) = '1' then
         current_group15m <= s1;

      else
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s161;

      end if;

   when s37 =>
      if ( x13 and x17 and x21 and x16 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s249;

      elsif ( x13 and x17 and x21 and not x16 and x18 and x15 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s249;

      elsif ( x13 and x17 and x21 and not x16 and x18 and not x15 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

      elsif ( x13 and x17 and x21 and not x16 and not x18 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s249;

      elsif ( x13 and x17 and not x21 and x22 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s249;

      elsif ( x13 and x17 and not x21 and not x22 and x15 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s249;

      elsif ( x13 and x17 and not x21 and not x22 and not x15 and x19 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s249;

      elsif ( x13 and x17 and not x21 and not x22 and not x15 and not x19 and x20 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s249;

      elsif ( x13 and x17 and not x21 and not x22 and not x15 and not x19 and not x20 and x16 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s249;

      elsif ( x13 and x17 and not x21 and not x22 and not x15 and not x19 and not x20 and not x16 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

      elsif ( x13 and not x17 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s249;

      else
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s249;

      end if;

   when s38 =>
      if ( x66 and x15 and x12 and x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x66 and x15 and x12 and not x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s250;

      elsif ( x66 and x15 and not x12 and x7 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x15 and not x12 and not x7 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( x66 and not x15 and x16 and x7 and x12 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s251;

      elsif ( x66 and not x15 and x16 and x7 and not x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( x66 and not x15 and x16 and not x7 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s252;

      elsif ( x66 and not x15 and not x16 and x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s253;

      elsif ( x66 and not x15 and not x16 and not x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      end if;

   when s39 =>
      if ( x65 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x20 and x21 and x15 and x8 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s254;

      elsif ( not x65 and not x20 and x21 and x15 and not x8 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s198;

      elsif ( not x65 and not x20 and x21 and not x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x65 and not x20 and x21 and not x15 and not x16 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s209;

      else
         y3 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s42;

      end if;

   when s40 =>
      if ( x66 and x65 and x60 and x61 and x15 and x2 and x12 and x7 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s67;

      elsif ( x66 and x65 and x60 and x61 and x15 and x2 and x12 and not x7 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s131;

      elsif ( x66 and x65 and x60 and x61 and x15 and x2 and not x12 and x7 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s255;

      elsif ( x66 and x65 and x60 and x61 and x15 and x2 and not x12 and not x7 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s254;

      elsif ( x66 and x65 and x60 and x61 and x15 and not x2 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s255;

      elsif ( x66 and x65 and x60 and x61 and not x15 and x16 and x7 and x12 and x2 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s256;

      elsif ( x66 and x65 and x60 and x61 and not x15 and x16 and x7 and x12 and not x2 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s255;

      elsif ( x66 and x65 and x60 and x61 and not x15 and x16 and x7 and not x12 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s255;

      elsif ( x66 and x65 and x60 and x61 and not x15 and x16 and not x7 and x12 and x9 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s255;

      elsif ( x66 and x65 and x60 and x61 and not x15 and x16 and not x7 and x12 and not x9 and x11 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s255;

      elsif ( x66 and x65 and x60 and x61 and not x15 and x16 and not x7 and x12 and not x9 and not x11 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and x65 and x60 and x61 and not x15 and x16 and not x7 and x12 and not x9 and not x11 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and x65 and x60 and x61 and not x15 and x16 and not x7 and x12 and not x9 and not x11 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x66 and x65 and x60 and x61 and not x15 and x16 and not x7 and x12 and not x9 and not x11 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x66 and x65 and x60 and x61 and not x15 and x16 and not x7 and not x12 and x11 and x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s255;

      elsif ( x66 and x65 and x60 and x61 and not x15 and x16 and not x7 and not x12 and x11 and not x10 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and x65 and x60 and x61 and not x15 and x16 and not x7 and not x12 and x11 and not x10 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and x65 and x60 and x61 and not x15 and x16 and not x7 and not x12 and x11 and not x10 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x66 and x65 and x60 and x61 and not x15 and x16 and not x7 and not x12 and x11 and not x10 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x66 and x65 and x60 and x61 and not x15 and x16 and not x7 and not x12 and not x11 and x8 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s255;

      elsif ( x66 and x65 and x60 and x61 and not x15 and x16 and not x7 and not x12 and not x11 and not x8 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and x65 and x60 and x61 and not x15 and x16 and not x7 and not x12 and not x11 and not x8 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and x65 and x60 and x61 and not x15 and x16 and not x7 and not x12 and not x11 and not x8 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x66 and x65 and x60 and x61 and not x15 and x16 and not x7 and not x12 and not x11 and not x8 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x66 and x65 and x60 and x61 and not x15 and not x16 and x2 and x7 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s257;

      elsif ( x66 and x65 and x60 and x61 and not x15 and not x16 and x2 and not x7 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      elsif ( x66 and x65 and x60 and x61 and not x15 and not x16 and not x2 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s255;

      elsif ( x66 and x65 and x60 and not x61 and x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and x60 and not x61 and not x11 and x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and x60 and not x61 and not x11 and not x7 and x16 and x15 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and x65 and x60 and not x61 and not x11 and not x7 and x16 and x15 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and x65 and x60 and not x61 and not x11 and not x7 and x16 and x15 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x66 and x65 and x60 and not x61 and not x11 and not x7 and x16 and x15 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x66 and x65 and x60 and not x61 and not x11 and not x7 and x16 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and x60 and not x61 and not x11 and not x7 and not x16 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x60 and x61 and x62 and x16 and x11 and x12 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s153;

      elsif ( x66 and x65 and not x60 and x61 and x62 and x16 and x11 and not x12 and x13 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s153;

      elsif ( x66 and x65 and not x60 and x61 and x62 and x16 and x11 and not x12 and not x13 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s154;

      elsif ( x66 and x65 and not x60 and x61 and x62 and x16 and not x11 and x13 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s63;

      elsif ( x66 and x65 and not x60 and x61 and x62 and x16 and not x11 and not x13 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( x66 and x65 and not x60 and x61 and x62 and not x16 and x17 and x11 and x13 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s258;

      elsif ( x66 and x65 and not x60 and x61 and x62 and not x16 and x17 and x11 and not x13 and x2 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x66 and x65 and not x60 and x61 and x62 and not x16 and x17 and x11 and not x13 and not x2 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( x66 and x65 and not x60 and x61 and x62 and not x16 and x17 and not x11 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s258;

      elsif ( x66 and x65 and not x60 and x61 and x62 and not x16 and not x17 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( x66 and x65 and not x60 and x61 and not x62 and x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x60 and x61 and not x62 and not x11 and x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x60 and x61 and not x62 and not x11 and not x7 and x16 and x15 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and x65 and not x60 and x61 and not x62 and not x11 and not x7 and x16 and x15 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and x65 and not x60 and x61 and not x62 and not x11 and not x7 and x16 and x15 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x66 and x65 and not x60 and x61 and not x62 and not x11 and not x7 and x16 and x15 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x66 and x65 and not x60 and x61 and not x62 and not x11 and not x7 and x16 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x60 and x61 and not x62 and not x11 and not x7 and not x16 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x60 and not x61 and x62 and x18 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and x65 and not x60 and not x61 and x62 and x18 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and x65 and not x60 and not x61 and x62 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x60 and not x61 and x62 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x60 and not x61 and not x62 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and x65 and not x60 and not x61 and not x62 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and x65 and not x60 and not x61 and not x62 and x19 and not x13 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x60 and not x61 and not x62 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and x21 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x21 and x22 and x23 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x66 and not x65 and not x21 and x22 and not x23 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x21 and not x22 and x23 and x19 and x14 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( x66 and not x65 and not x21 and not x22 and x23 and x19 and not x14 and x13 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( x66 and not x65 and not x21 and not x22 and x23 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x21 and not x22 and x23 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x21 and not x22 and not x23 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x66 and x65 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and not x20 and x21 ) = '1' then
         current_group15m <= s39;

      elsif ( not x66 and not x65 and x67 and not x20 and not x21 and x18 and x15 and x8 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x66 and not x65 and x67 and not x20 and not x21 and x18 and x15 and not x8 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s198;

      elsif ( not x66 and not x65 and x67 and not x20 and not x21 and x18 and not x15 and x16 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and not x65 and x67 and not x20 and not x21 and x18 and not x15 and not x16 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s209;

      elsif ( not x66 and not x65 and x67 and not x20 and not x21 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( not x66 and not x65 and not x67 and x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and x3 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s107;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and x3 and not x2 ) = '1' then
         current_group15m <= s40;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x3 ) = '1' then
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s179;

      elsif ( not x66 and not x65 and not x67 and not x21 and not x22 and x2 and x11 ) = '1' then
         current_group15m <= s40;

      elsif ( not x66 and not x65 and not x67 and not x21 and not x22 and x2 and not x11 ) = '1' then
         current_group15m <= s40;

      else
         y4 <= '1' ;
         current_group15m <= s43;

      end if;

   when s41 =>
      if ( x20 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x20 and x21 and x15 and x8 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s254;

      elsif ( not x20 and x21 and x15 and not x8 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s198;

      elsif ( not x20 and x21 and not x15 and x16 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s59;

      elsif ( not x20 and x21 and not x15 and not x16 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s209;

      elsif ( not x20 and not x21 and x17 and x13 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x20 and not x21 and x17 and not x13 and x12 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x20 and not x21 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s42 =>
      if ( x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x15 and x8 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x21 and x15 and not x8 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s198;

      elsif ( not x21 and not x15 and x16 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      else
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s209;

      end if;

   when s43 =>
      if ( x65 and x66 and x68 and x21 and x20 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s259;

      elsif ( x65 and x66 and x68 and x21 and not x20 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x66 and x68 and x21 and not x20 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x66 and x68 and x21 and not x20 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x68 and x21 and not x20 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x68 and not x21 and x19 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x66 and x68 and not x21 and x19 and not x14 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x66 and x68 and not x21 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x68 and not x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and x16 and x7 and x12 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and x16 and x7 and not x12 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s260;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and x16 and not x7 and x12 and x14 and x11 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         y10 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s261;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and x16 and not x7 and x12 and x14 and not x11 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and x16 and not x7 and x12 and not x14 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and x16 and not x7 and x12 and not x14 and x19 and not x13 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and x16 and not x7 and x12 and not x14 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and x16 and not x7 and not x12 and x13 and x11 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s262;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and x16 and not x7 and not x12 and x13 and not x11 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and x16 and not x7 and not x12 and not x13 and x19 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and x16 and not x7 and not x12 and not x13 and x19 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and x16 and not x7 and not x12 and not x13 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and not x16 and x11 and x7 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and not x16 and x11 and not x7 and x12 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and not x16 and x11 and not x7 and not x12 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s257;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and not x16 and not x11 and x1 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and not x16 and not x11 and not x1 and x12 and x3 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s74;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and not x16 and not x11 and not x1 and x12 and not x3 and x7 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s69;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and not x16 and not x11 and not x1 and x12 and not x3 and not x7 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s257;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and not x16 and not x11 and not x1 and not x12 and x7 and x3 ) = '1' then
         y2 <= '1' ;
         y10 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s263;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and not x16 and not x11 and not x1 and not x12 and x7 and not x3 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and not x16 and not x11 and not x1 and not x12 and not x7 and x3 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s74;

      elsif ( x65 and x66 and not x68 and x61 and x60 and x15 and not x16 and not x11 and not x1 and not x12 and not x7 and not x3 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and x1 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and x7 and x12 and x3 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s74;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and x7 and x12 and not x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s257;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and x7 and not x12 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s74;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and not x7 and x12 and x11 and x3 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s74;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and not x7 and x12 and x11 and not x3 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and not x7 and x12 and not x11 and x9 and x3 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s74;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and not x7 and x12 and not x11 and x9 and not x3 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and not x7 and x12 and not x11 and not x9 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and not x7 and x12 and not x11 and not x9 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and not x7 and x12 and not x11 and not x9 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and not x7 and x12 and not x11 and not x9 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and not x7 and not x12 and x11 and x10 and x3 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s74;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and not x7 and not x12 and x11 and x10 and not x3 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and not x7 and not x12 and x11 and not x10 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and not x7 and not x12 and x11 and not x10 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and not x7 and not x12 and x11 and not x10 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and not x7 and not x12 and x11 and not x10 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and not x7 and not x12 and not x11 and x8 and x3 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s74;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and not x7 and not x12 and not x11 and x8 and not x3 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and not x7 and not x12 and not x11 and not x8 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and not x7 and not x12 and not x11 and not x8 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and not x7 and not x12 and not x11 and not x8 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and x16 and not x7 and not x12 and not x11 and not x8 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and not x16 and x3 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s74;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and not x16 and not x3 and x7 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s257;

      elsif ( x65 and x66 and not x68 and x61 and x60 and not x15 and not x1 and not x16 and not x3 and not x7 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s264;

      elsif ( x65 and x66 and not x68 and x61 and not x60 and x62 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and x66 and not x68 and x61 and not x60 and not x62 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and not x68 and x61 and not x60 and not x62 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and not x68 and x61 and not x60 and not x62 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x66 and not x68 and x61 and not x60 and not x62 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x66 and not x68 and not x61 and x60 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and not x68 and not x61 and x60 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and not x68 and not x61 and x60 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x66 and not x68 and not x61 and x60 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x66 and not x68 and not x61 and not x60 and x62 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( x65 and x66 and not x68 and not x61 and not x60 and not x62 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and not x66 and x68 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and x68 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and x68 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x68 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x68 and x21 and x18 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x65 and not x66 and not x68 and x21 and not x18 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x68 and x21 and not x18 and x19 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x68 and x21 and not x18 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x68 and x21 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x68 and not x21 and x23 and x22 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( x65 and not x66 and not x68 and not x21 and x23 and x22 and not x19 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x66 and not x68 and not x21 and x23 and x22 and not x19 and x17 and not x14 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x66 and not x68 and not x21 and x23 and x22 and not x19 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x68 and not x21 and x23 and x22 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x68 and not x21 and x23 and not x22 and x20 and x14 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x66 and not x68 and not x21 and x23 and not x22 and x20 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x66 and not x68 and not x21 and x23 and not x22 and x20 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x68 and not x21 and x23 and not x22 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x68 and not x21 and not x23 and x18 and x14 and x22 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x68 and not x21 and not x23 and x18 and x14 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x66 and not x68 and not x21 and not x23 and x18 and not x14 and x13 and x22 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x68 and not x21 and not x23 and x18 and not x14 and x13 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x66 and not x68 and not x21 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x68 and not x21 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x20 and x18 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x67 and x20 and x18 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x67 and x20 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x20 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and x21 and x68 and x3 and x4 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( not x65 and not x67 and x21 and x68 and x3 and not x4 and x5 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( not x65 and not x67 and x21 and x68 and x3 and not x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and x21 and x68 and not x3 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and x21 and not x68 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s108;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and x19 and x12 and x17 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s246;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and x19 and x12 and not x17 ) = '1' then
         y8 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s266;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and x19 and not x12 and x17 and x8 and x16 ) = '1' then
         y8 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s267;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and x19 and not x12 and x17 and x8 and not x16 ) = '1' then
         y10 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s268;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and x19 and not x12 and x17 and not x8 and x6 and x7 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and x19 and not x12 and x17 and not x8 and x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and x19 and not x12 and x17 and not x8 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and x19 and not x12 and not x17 and x7 and x16 ) = '1' then
         y23 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s269;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and x19 and not x12 and not x17 and x7 and not x16 ) = '1' then
         y10 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s268;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and x19 and not x12 and not x17 and not x7 and x6 and x8 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and x19 and not x12 and not x17 and not x7 and x6 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and x19 and not x12 and not x17 and not x7 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and not x19 and x16 and x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s270;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and not x19 and x16 and not x12 and x17 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s109;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and not x19 and x16 and not x12 and not x17 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s271;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and not x19 and not x16 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and not x19 and not x16 and not x2 and x3 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and not x19 and not x16 and not x2 and not x3 and x17 and x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s272;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and not x19 and not x16 and not x2 and not x3 and x17 and not x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s272;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and not x19 and not x16 and not x2 and not x3 and not x17 and x12 ) = '1' then
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s273;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and x18 and not x19 and not x16 and not x2 and not x3 and not x17 and not x12 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s273;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and x12 and x3 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and x12 and not x3 and x17 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s271;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and x12 and not x3 and not x17 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and not x12 and x16 and x17 and x3 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and not x12 and x16 and x17 and not x3 ) = '1' then
         y10 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s273;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and not x12 and x16 and not x17 and x15 and x3 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and not x12 and x16 and not x17 and x15 and not x3 ) = '1' then
         y10 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s273;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and not x12 and x16 and not x17 and not x15 and x6 and x7 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and not x12 and x16 and not x17 and not x15 and x6 and not x7 and x8 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and not x12 and x16 and not x17 and not x15 and x6 and not x7 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and not x12 and x16 and not x17 and not x15 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and not x12 and not x16 and x17 and x14 and x3 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and not x12 and not x16 and x17 and x14 and not x3 ) = '1' then
         y10 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s273;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and not x12 and not x16 and x17 and not x14 and x6 and x7 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and not x12 and not x16 and x17 and not x14 and x6 and not x7 and x8 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and not x12 and not x16 and x17 and not x14 and x6 and not x7 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and not x12 and not x16 and x17 and not x14 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and not x12 and not x16 and not x17 and x13 and x6 and x7 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and not x12 and not x16 and not x17 and x13 and x6 and not x7 and x8 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and not x12 and not x16 and not x17 and x13 and x6 and not x7 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and not x12 and not x16 and not x17 and x13 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and not x12 and not x16 and not x17 and not x13 and x3 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and x19 and not x12 and not x16 and not x17 and not x13 and not x3 ) = '1' then
         y10 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s273;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and not x19 and x3 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and not x19 and not x3 and x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s271;

      elsif ( not x65 and not x67 and not x21 and x22 and x68 and not x18 and not x2 and not x19 and not x3 and not x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s272;

      elsif ( not x65 and not x67 and not x21 and x22 and not x68 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s126;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and x18 and x19 and x15 and x17 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s246;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and x18 and x19 and x15 and not x17 ) = '1' then
         y8 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s266;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and x18 and x19 and not x15 and x16 and x17 ) = '1' then
         y8 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s267;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and x18 and x19 and not x15 and x16 and not x17 ) = '1' then
         y23 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s269;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and x18 and x19 and not x15 and not x16 and x17 and x10 ) = '1' then
         y10 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s273;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and x18 and x19 and not x15 and not x16 and x17 and not x10 and x9 and x8 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and x18 and x19 and not x15 and not x16 and x17 and not x10 and x9 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and x18 and x19 and not x15 and not x16 and x17 and not x10 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and x18 and x19 and not x15 and not x16 and not x17 and x9 ) = '1' then
         y10 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s273;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and x18 and x19 and not x15 and not x16 and not x17 and not x9 and x8 and x10 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and x18 and x19 and not x15 and not x16 and not x17 and not x9 and x8 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and x18 and x19 and not x15 and not x16 and not x17 and not x9 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and x18 and not x19 and x16 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s274;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and x18 and not x19 and not x16 and x2 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s173;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and x18 and not x19 and not x16 and not x2 and x5 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s275;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and x18 and not x19 and not x16 and not x2 and not x5 and x15 ) = '1' then
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s273;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and x18 and not x19 and not x16 and not x2 and not x5 and not x15 ) = '1' then
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s273;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and x2 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s173;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and x15 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s275;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and not x15 and x16 and x17 and x5 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s275;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and not x15 and x16 and x17 and not x5 ) = '1' then
         y10 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s273;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and not x15 and x16 and not x17 and x14 and x5 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s275;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and not x15 and x16 and not x17 and x14 and not x5 ) = '1' then
         y10 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s273;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and not x15 and x16 and not x17 and not x14 and x8 and x9 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and not x15 and x16 and not x17 and not x14 and x8 and not x9 and x10 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and not x15 and x16 and not x17 and not x14 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and not x15 and x16 and not x17 and not x14 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and not x15 and not x16 and x17 and x13 and x5 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s275;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and not x15 and not x16 and x17 and x13 and not x5 ) = '1' then
         y10 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s273;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and not x15 and not x16 and x17 and not x13 and x8 and x9 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and not x15 and not x16 and x17 and not x13 and x8 and not x9 and x10 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and not x15 and not x16 and x17 and not x13 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and not x15 and not x16 and x17 and not x13 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and not x15 and not x16 and not x17 and x12 and x5 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s275;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and not x15 and not x16 and not x17 and x12 and not x5 ) = '1' then
         y10 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s273;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and not x15 and not x16 and not x17 and not x12 and x8 and x9 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and not x15 and not x16 and not x17 and not x12 and x8 and not x9 and x10 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and not x15 and not x16 and not x17 and not x12 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and x19 and not x15 and not x16 and not x17 and not x12 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and not x19 and x5 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s275;

      elsif ( not x65 and not x67 and not x21 and not x22 and x68 and not x18 and not x2 and not x19 and not x5 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s274;

      else
         current_group15m <= s1;

      end if;

   when s44 =>
      if ( x65 and x66 and x67 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x65 and x66 and not x67 and x21 and x20 ) = '1' then
         y9 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s276;

      elsif ( x65 and x66 and not x67 and x21 and not x20 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( x65 and x66 and not x67 and not x21 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( x65 and not x66 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( not x65 and x20 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( not x65 and not x20 and x21 ) = '1' then
         y4 <= '1' ;
         y16 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s45;

      else
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      end if;

   when s45 =>
      if ( x20 ) = '1' then
         current_group15m <= s1;

      else
         y2 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s277;

      end if;

   when s46 =>
      if ( x24 and x26 and x19 ) = '1' then
         current_group15m <= s46;

      elsif ( x24 and x26 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x24 and not x26 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      elsif ( not x24 and x25 and x26 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and not x26 and x15 and x6 and x10 and x11 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s188;

      elsif ( not x24 and x25 and not x26 and x15 and x6 and x10 and not x11 and x12 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s172;

      elsif ( not x24 and x25 and not x26 and x15 and x6 and x10 and not x11 and not x12 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x24 and x25 and not x26 and x15 and x6 and not x10 ) = '1' then
         y8 <= '1' ;
         y17 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s164;

      elsif ( not x24 and x25 and not x26 and x15 and not x6 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and x12 and x10 and x8 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and x12 and x10 and not x8 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and x12 and x10 and not x8 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and x12 and x10 and not x8 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and x12 and x10 and not x8 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and x12 and not x10 and x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and x12 and not x10 and not x7 and x11 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and x12 and not x10 and not x7 and not x11 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and x12 and not x10 and not x7 and not x11 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and x12 and not x10 and not x7 and not x11 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and x12 and not x10 and not x7 and not x11 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and not x12 and x10 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and not x12 and not x10 and x11 and x9 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and not x12 and not x10 and x11 and not x9 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and not x12 and not x10 and x11 and not x9 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and not x12 and not x10 and x11 and not x9 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and not x12 and not x10 and x11 and not x9 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and not x12 and not x10 and not x11 and x8 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and not x12 and not x10 and not x11 and x8 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and not x12 and not x10 and not x11 and x8 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and not x12 and not x10 and not x11 and x8 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and not x26 and not x15 and x16 and not x12 and not x10 and not x11 and not x8 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x24 and x25 and not x26 and not x15 and not x16 and x6 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x24 and x25 and not x26 and not x15 and not x16 and not x6 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x24 and not x25 and x26 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      elsif ( not x24 and not x25 and not x26 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x24 and not x25 and not x26 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x24 and not x25 and not x26 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s47 =>
      if ( x68 and x20 and x18 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x68 and x20 and x18 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x68 and x20 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x68 and x20 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x68 and not x20 and x21 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( x68 and not x20 and x21 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( x68 and not x20 and x21 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x68 and not x20 and x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x68 and not x20 and not x21 and x17 and x13 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( x68 and not x20 and not x21 and x17 and not x13 and x12 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( x68 and not x20 and not x21 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x68 and not x20 and not x21 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x68 and x24 and x26 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s279;

      elsif ( not x68 and x24 and not x26 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x68 and x24 and not x26 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x68 and x24 and not x26 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x68 and x24 and not x26 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x68 and not x24 and x25 and x26 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x68 and not x24 and x25 and not x26 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x68 and not x24 and not x25 and x26 ) = '1' then
         current_group15m <= s1;

      elsif ( not x68 and not x24 and not x25 and not x26 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x68 and not x24 and not x25 and not x26 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x68 and not x24 and not x25 and not x26 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s48 =>
      if ( x66 and x21 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x66 and x21 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x66 and x21 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x21 and x22 and x23 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x66 and not x21 and x22 and not x23 and x18 and x14 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and not x21 and x22 and not x23 and x18 and not x14 and x13 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and not x21 and x22 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x21 and x22 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x21 and not x22 and x23 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      elsif ( x66 and not x21 and not x22 and not x23 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s180;

      elsif ( not x66 and x24 and x26 and x18 and x15 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x66 and x24 and x26 and x18 and not x15 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x66 and x24 and x26 and x18 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x24 and x26 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x24 and not x26 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x24 and x25 and x26 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x66 and not x24 and x25 and x26 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x66 and not x24 and x25 and x26 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s48;

      elsif ( not x66 and not x24 and x25 and x26 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x24 and x25 and not x26 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x24 and not x25 and x26 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and not x24 and not x25 and x26 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and not x24 and not x25 and x26 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x24 and not x25 and x26 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x24 and not x25 and not x26 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x66 and not x24 and not x25 and not x26 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x66 and not x24 and not x25 and not x26 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s49 =>
      if ( x24 and x26 and x18 and x15 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( x24 and x26 and x18 and not x15 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( x24 and x26 and x18 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x24 and x26 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x24 and not x26 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x25 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x25 and x19 and not x14 and not x13 and x26 ) = '1' then
         current_group15m <= s49;

      elsif ( not x24 and x25 and x19 and not x14 and not x13 and not x26 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and x26 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x24 and not x25 and x26 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x24 and not x25 and x26 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and x26 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and not x26 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x24 and not x25 and not x26 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x24 and not x25 and not x26 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s50 =>
      if ( x65 and x22 and x17 and x18 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x22 and x17 and not x18 and x19 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x22 and x17 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x22 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x22 and x18 and x13 and x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and not x22 and x18 and x13 and not x23 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and not x22 and x18 and not x13 and x12 and x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and not x22 and x18 and not x13 and x12 and not x23 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and not x22 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x22 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x26 and x24 ) = '1' then
         y12 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s49;

      elsif ( not x65 and x26 and not x24 and x25 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x26 and not x24 and not x25 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x65 and x26 and not x24 and not x25 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x65 and x26 and not x24 and not x25 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x26 and not x24 and not x25 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x26 and x24 ) = '1' then
         y15 <= '1' ;
         y112 <= '1' ;
         current_group15m <= s280;

      elsif ( not x65 and not x26 and not x24 and x25 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x26 and not x24 and x25 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x26 and not x24 and x25 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x26 and not x24 and x25 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x26 and not x24 and not x25 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x65 and not x26 and not x24 and not x25 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x65 and not x26 and not x24 and not x25 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s51 =>
      if ( x65 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x24 and x26 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x24 and not x26 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and x24 and not x26 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and x24 and not x26 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x24 and not x26 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x24 and x25 and x26 ) = '1' then
         y11 <= '1' ;
         y16 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s281;

      elsif ( not x65 and not x24 and x25 and not x26 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and not x24 and not x25 and x26 and x3 and x16 and x11 ) = '1' then
         y15 <= '1' ;
         y112 <= '1' ;
         current_group15m <= s46;

      elsif ( not x65 and not x24 and not x25 and x26 and x3 and x16 and not x11 and x12 ) = '1' then
         y15 <= '1' ;
         y112 <= '1' ;
         current_group15m <= s46;

      elsif ( not x65 and not x24 and not x25 and x26 and x3 and x16 and not x11 and not x12 and x10 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x65 and not x24 and not x25 and x26 and x3 and x16 and not x11 and not x12 and not x10 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s50;

      elsif ( not x65 and not x24 and not x25 and x26 and x3 and not x16 and x17 and x10 and x12 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( not x65 and not x24 and not x25 and x26 and x3 and not x16 and x17 and x10 and not x12 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s17;

      elsif ( not x65 and not x24 and not x25 and x26 and x3 and not x16 and x17 and not x10 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( not x65 and not x24 and not x25 and x26 and x3 and not x16 and not x17 ) = '1' then
         y15 <= '1' ;
         y112 <= '1' ;
         current_group15m <= s46;

      elsif ( not x65 and not x24 and not x25 and x26 and not x3 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x65 and not x24 and not x25 and not x26 and x4 and x15 and x11 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      elsif ( not x65 and not x24 and not x25 and not x26 and x4 and x15 and not x11 and x12 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      elsif ( not x65 and not x24 and not x25 and not x26 and x4 and x15 and not x11 and not x12 and x10 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x65 and not x24 and not x25 and not x26 and x4 and x15 and not x11 and not x12 and not x10 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s50;

      elsif ( not x65 and not x24 and not x25 and not x26 and x4 and not x15 and x16 and x10 and x12 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( not x65 and not x24 and not x25 and not x26 and x4 and not x15 and x16 and x10 and not x12 ) = '1' then
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s239;

      elsif ( not x65 and not x24 and not x25 and not x26 and x4 and not x15 and x16 and not x10 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( not x65 and not x24 and not x25 and not x26 and x4 and not x15 and not x16 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      else
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s165;

      end if;

   when s52 =>
      if ( x66 and x21 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( x66 and not x21 and x22 and x10 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s219;

      elsif ( x66 and not x21 and x22 and not x10 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s28;

      elsif ( x66 and not x21 and not x22 ) = '1' then
         y8 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s82;

      elsif ( not x66 and x24 and x11 and x26 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x66 and x24 and x11 and not x26 and x13 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x66 and x24 and x11 and not x26 and x13 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x66 and x24 and x11 and not x26 and x13 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x24 and x11 and not x26 and x13 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x24 and x11 and not x26 and not x13 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s282;

      elsif ( not x66 and x24 and not x11 and x26 and x12 and x13 and x16 and x18 and x15 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x66 and x24 and not x11 and x26 and x12 and x13 and x16 and x18 and not x15 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x66 and x24 and not x11 and x26 and x12 and x13 and x16 and x18 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x24 and not x11 and x26 and x12 and x13 and x16 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x24 and not x11 and x26 and x12 and x13 and not x16 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x66 and x24 and not x11 and x26 and x12 and not x13 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x66 and x24 and not x11 and x26 and not x12 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x66 and x24 and not x11 and not x26 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x66 and x24 and not x11 and not x26 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x66 and x24 and not x11 and not x26 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x24 and not x11 and not x26 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x24 and x25 and x26 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x66 and not x24 and x25 and not x26 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x24 and not x25 and x26 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and not x24 and not x25 and x26 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and not x24 and not x25 and x26 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x24 and not x25 and x26 and not x18 ) = '1' then
         current_group15m <= s1;

      else
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      end if;

   when s53 =>
      if ( x66 and x67 and x65 and x22 ) = '1' then
         y9 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s111;

      elsif ( x66 and x67 and x65 and not x22 and x23 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x66 and x67 and x65 and not x22 and not x23 and x18 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x67 and x65 and not x22 and not x23 and x18 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x67 and x65 and not x22 and not x23 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x67 and x65 and not x22 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x67 and not x65 and x63 and x15 and x64 and x8 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( x66 and x67 and not x65 and x63 and x15 and x64 and not x8 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x66 and x67 and not x65 and x63 and x15 and not x64 and x16 and x8 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x67 and not x65 and x63 and x15 and not x64 and x16 and x8 and not x14 and x7 ) = '1' then
         y24 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s157;

      elsif ( x66 and x67 and not x65 and x63 and x15 and not x64 and x16 and x8 and not x14 and not x7 and x12 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s65;

      elsif ( x66 and x67 and not x65 and x63 and x15 and not x64 and x16 and x8 and not x14 and not x7 and not x12 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( x66 and x67 and not x65 and x63 and x15 and not x64 and x16 and not x8 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and x67 and not x65 and x63 and x15 and not x64 and x16 and not x8 and not x14 and x7 ) = '1' then
         y26 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s158;

      elsif ( x66 and x67 and not x65 and x63 and x15 and not x64 and x16 and not x8 and not x14 and not x7 and x13 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s65;

      elsif ( x66 and x67 and not x65 and x63 and x15 and not x64 and x16 and not x8 and not x14 and not x7 and not x13 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( x66 and x67 and not x65 and x63 and x15 and not x64 and not x16 and x7 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s159;

      elsif ( x66 and x67 and not x65 and x63 and x15 and not x64 and not x16 and not x7 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( x66 and x67 and not x65 and x63 and x15 and not x64 and not x16 and not x7 and not x3 and x5 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( x66 and x67 and not x65 and x63 and x15 and not x64 and not x16 and not x7 and not x3 and not x5 and x8 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( x66 and x67 and not x65 and x63 and x15 and not x64 and not x16 and not x7 and not x3 and not x5 and not x8 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and x16 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s151;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and x16 and not x64 and x8 and x7 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and x16 and not x64 and x8 and x7 and not x3 and x5 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and x16 and not x64 and x8 and x7 and not x3 and not x5 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s151;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and x16 and not x64 and x8 and not x7 and x9 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and x16 and not x64 and x8 and not x7 and x9 and not x3 and x5 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and x16 and not x64 and x8 and not x7 and x9 and not x3 and not x5 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s151;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and x16 and not x64 and x8 and not x7 and not x9 and x3 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and x16 and not x64 and x8 and not x7 and not x9 and not x3 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and x16 and not x64 and not x8 and x7 and x11 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and x16 and not x64 and not x8 and x7 and x11 and not x3 and x5 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and x16 and not x64 and not x8 and x7 and x11 and not x3 and not x5 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s151;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and x16 and not x64 and not x8 and x7 and not x11 and x3 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and x16 and not x64 and not x8 and x7 and not x11 and not x3 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and x16 and not x64 and not x8 and not x7 and x10 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and x16 and not x64 and not x8 and not x7 and x10 and not x3 and x5 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and x16 and not x64 and not x8 and not x7 and x10 and not x3 and not x5 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s151;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and x16 and not x64 and not x8 and not x7 and not x10 and x3 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and x16 and not x64 and not x8 and not x7 and not x10 and not x3 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and not x16 and x64 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s135;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and not x16 and not x64 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and not x16 and not x64 and not x3 and x5 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( x66 and x67 and not x65 and x63 and not x15 and not x16 and not x64 and not x3 and not x5 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s135;

      elsif ( x66 and x67 and not x65 and not x63 and x64 and x19 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x66 and x67 and not x65 and not x63 and x64 and x19 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x66 and x67 and not x65 and not x63 and x64 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x67 and not x65 and not x63 and x64 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x67 and not x65 and not x63 and not x64 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and x65 and x61 and x60 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and not x67 and x65 and x61 and x60 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and not x67 and x65 and x61 and x60 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x66 and not x67 and x65 and x61 and x60 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x66 and not x67 and x65 and x61 and not x60 and x62 and x11 and x13 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x66 and not x67 and x65 and x61 and not x60 and x62 and x11 and x13 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x66 and not x67 and x65 and x61 and not x60 and x62 and x11 and x13 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and x65 and x61 and not x60 and x62 and x11 and x13 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and x65 and x61 and not x60 and x62 and x11 and not x13 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( x66 and not x67 and x65 and x61 and not x60 and x62 and not x11 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x66 and not x67 and x65 and x61 and not x60 and x62 and not x11 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x66 and not x67 and x65 and x61 and not x60 and x62 and not x11 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and x65 and x61 and not x60 and x62 and not x11 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and x65 and x61 and not x60 and not x62 and x7 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x66 and not x67 and x65 and x61 and not x60 and not x62 and not x7 ) = '1' then
         current_group15m <= s39;

      elsif ( x66 and not x67 and x65 and not x61 and x60 and x7 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x66 and not x67 and x65 and not x61 and x60 and not x7 ) = '1' then
         current_group15m <= s39;

      elsif ( x66 and not x67 and x65 and not x61 and not x60 and x62 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( x66 and not x67 and x65 and not x61 and not x60 and not x62 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s258;

      elsif ( x66 and not x67 and not x65 and x21 and x68 and x9 and x8 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x66 and not x67 and not x65 and x21 and x68 and x9 and not x8 and x7 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x66 and not x67 and not x65 and x21 and x68 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and x21 and x68 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and x21 and not x68 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x66 and not x67 and not x65 and x21 and not x68 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x66 and not x67 and not x65 and x21 and not x68 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and x21 and not x68 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and x68 and x5 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and x68 and not x5 and x17 and x10 and x15 and x6 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s283;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and x68 and not x5 and x17 and x10 and x15 and not x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and x68 and not x5 and x17 and x10 and not x15 and x16 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and x68 and not x5 and x17 and x10 and not x15 and not x16 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and x68 and not x5 and x17 and not x10 and x6 ) = '1' then
         y13 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s284;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and x68 and not x5 and x17 and not x10 and not x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and x68 and not x5 and not x17 and x18 and x6 and x10 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s219;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and x68 and not x5 and not x17 and x18 and x6 and not x10 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and x68 and not x5 and not x17 and x18 and not x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and x68 and not x5 and not x17 and not x18 and x6 and x10 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s219;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and x68 and not x5 and not x17 and not x18 and x6 and not x10 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s28;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and x68 and not x5 and not x17 and not x18 and not x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and not x68 and x23 and x18 and x15 and x10 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and not x68 and x23 and x18 and x15 and not x10 and x12 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and not x68 and x23 and x18 and x15 and not x10 and not x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s285;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and not x68 and x23 and x18 and not x15 and x16 and x10 and x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s286;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and not x68 and x23 and x18 and not x15 and x16 and x10 and not x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and not x68 and x23 and x18 and not x15 and x16 and not x10 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s286;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and not x68 and x23 and x18 and not x15 and not x16 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and not x68 and x23 and not x18 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and not x68 and not x23 and x18 and x14 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and not x68 and not x23 and x18 and not x14 and x13 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and not x68 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and x22 and not x68 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and x17 and x10 and x15 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and x17 and x10 and not x15 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and x17 and not x10 and x15 and x6 and x14 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and x17 and not x10 and x15 and x6 and not x14 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s287;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and x17 and not x10 and x15 and not x6 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and x17 and not x10 and x15 and not x6 and x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and x17 and not x10 and x15 and not x6 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and x17 and not x10 and not x15 and x5 and x14 ) = '1' then
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s288;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and x17 and not x10 and not x15 and x5 and not x14 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s287;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and x17 and not x10 and not x15 and not x5 and x4 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and x17 and not x10 and not x15 and not x5 and x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and x17 and not x10 and not x15 and not x5 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and not x17 and x14 and x10 ) = '1' then
         y13 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s289;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and not x17 and x14 and not x10 and x15 ) = '1' then
         y13 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s284;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and not x17 and x14 and not x10 and not x15 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s290;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and not x17 and not x14 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and not x17 and not x14 and not x2 and x15 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and not x17 and not x14 and not x2 and x15 and not x3 and x10 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s291;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and not x17 and not x14 and not x2 and x15 and not x3 and not x10 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s292;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and not x17 and not x14 and not x2 and not x15 and x10 and x3 ) = '1' then
         y2 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s221;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and not x17 and not x14 and not x2 and not x15 and x10 and not x3 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and not x17 and not x14 and not x2 and not x15 and not x10 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and x16 and not x17 and not x14 and not x2 and not x15 and not x10 and not x3 ) = '1' then
         y14 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s216;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and x10 and x15 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and x10 and x15 and not x3 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s290;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and x10 and not x15 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and not x10 and x14 and x15 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and not x10 and x14 and x15 and not x3 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and not x10 and x14 and not x15 and x13 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and not x10 and x14 and not x15 and x13 and not x3 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and not x10 and x14 and not x15 and not x13 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and not x10 and x14 and not x15 and not x13 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and not x10 and x14 and not x15 and not x13 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and not x10 and x14 and not x15 and not x13 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and x15 and x12 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and x15 and x12 and not x3 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and x15 and not x12 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and x15 and not x12 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and x15 and not x12 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and x15 and not x12 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and not x15 and x11 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and not x15 and x11 and not x3 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and not x15 and not x11 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and not x15 and not x11 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and not x15 and not x11 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and not x15 and not x11 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and not x17 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and not x17 and not x3 and x10 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s293;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and x68 and not x16 and not x2 and not x17 and not x3 and not x10 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s231;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and not x68 and x23 and x19 and x14 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and not x68 and x23 and x19 and not x14 and x13 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and not x68 and x23 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and not x68 and x23 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x67 and not x65 and not x21 and not x22 and not x68 and not x23 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x66 and x65 and x15 and x9 and x21 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x66 and x65 and x15 and x9 and not x21 and x23 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x66 and x65 and x15 and x9 and not x21 and not x23 ) = '1' then
         y15 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_group15m <= s294;

      elsif ( not x66 and x65 and x15 and not x9 and x21 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x66 and x65 and x15 and not x9 and not x21 and x23 and x6 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( not x66 and x65 and x15 and not x9 and not x21 and x23 and not x6 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x66 and x65 and x15 and not x9 and not x21 and not x23 and x6 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x66 and x65 and x15 and not x9 and not x21 and not x23 and not x6 ) = '1' then
         y15 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_group15m <= s294;

      elsif ( not x66 and x65 and not x15 and x21 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s212;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and x8 and x23 and x9 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and x8 and x23 and not x9 and x12 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and x8 and x23 and not x9 and not x12 and x20 and x14 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and x8 and x23 and not x9 and not x12 and x20 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and x8 and x23 and not x9 and not x12 and x20 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and x8 and x23 and not x9 and not x12 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and x8 and not x23 and x9 ) = '1' then
         y15 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_group15m <= s294;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and x8 and not x23 and not x9 and x12 ) = '1' then
         y15 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_group15m <= s294;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and x8 and not x23 and not x9 and not x12 and x18 and x14 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and x8 and not x23 and not x9 and not x12 and x18 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and x8 and not x23 and not x9 and not x12 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and x8 and not x23 and not x9 and not x12 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and not x8 and x23 and x9 and x10 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and not x8 and x23 and x9 and not x10 and x20 and x14 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and not x8 and x23 and x9 and not x10 and x20 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and not x8 and x23 and x9 and not x10 and x20 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and not x8 and x23 and x9 and not x10 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and not x8 and x23 and not x9 and x11 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and not x8 and x23 and not x9 and not x11 and x20 and x14 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and not x8 and x23 and not x9 and not x11 and x20 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and not x8 and x23 and not x9 and not x11 and x20 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and not x8 and x23 and not x9 and not x11 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and not x8 and not x23 and x9 and x10 ) = '1' then
         y15 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_group15m <= s294;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and not x8 and not x23 and x9 and not x10 and x18 and x14 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and not x8 and not x23 and x9 and not x10 and x18 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and not x8 and not x23 and x9 and not x10 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and not x8 and not x23 and x9 and not x10 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and not x8 and not x23 and not x9 and x11 ) = '1' then
         y15 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_group15m <= s294;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and not x8 and not x23 and not x9 and not x11 and x18 and x14 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and not x8 and not x23 and not x9 and not x11 and x18 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and not x8 and not x23 and not x9 and not x11 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x15 and not x21 and x16 and not x8 and not x23 and not x9 and not x11 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x15 and not x21 and not x16 and x23 and x6 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s205;

      elsif ( not x66 and x65 and not x15 and not x21 and not x16 and x23 and not x6 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x66 and x65 and not x15 and not x21 and not x16 and not x23 and x6 ) = '1' then
         y31 <= '1' ;
         current_group15m <= s96;

      elsif ( not x66 and x65 and not x15 and not x21 and not x16 and not x23 and not x6 ) = '1' then
         y15 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_group15m <= s294;

      elsif ( not x66 and not x65 and x24 and x26 and x18 and x15 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x66 and not x65 and x24 and x26 and x18 and not x15 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x66 and not x65 and x24 and x26 and x18 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x24 and x26 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x24 and not x26 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x66 and not x65 and not x24 and x25 and x26 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x66 and not x65 and not x24 and x25 and x26 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x66 and not x65 and not x24 and x25 and x26 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s53;

      elsif ( not x66 and not x65 and not x24 and x25 and x26 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x24 and x25 and not x26 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s189;

      elsif ( not x66 and not x65 and not x24 and not x25 and x26 and x16 and x10 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and not x65 and not x24 and not x25 and x26 and x16 and not x10 and x11 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and not x65 and not x24 and not x25 and x26 and x16 and not x10 and not x11 and x12 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and not x65 and not x24 and not x25 and x26 and x16 and not x10 and not x11 and not x12 ) = '1' then
         y12 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s49;

      elsif ( not x66 and not x65 and not x24 and not x25 and x26 and not x16 and x17 and x10 and x12 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s282;

      elsif ( not x66 and not x65 and not x24 and not x25 and x26 and not x16 and x17 and x10 and not x12 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s204;

      elsif ( not x66 and not x65 and not x24 and not x25 and x26 and not x16 and x17 and not x10 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s282;

      elsif ( not x66 and not x65 and not x24 and not x25 and x26 and not x16 and not x17 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      else
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      end if;

   when s54 =>
      if ( x65 and x21 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s139;

      elsif ( x65 and not x21 and x22 and x23 and x15 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      elsif ( x65 and not x21 and x22 and x23 and not x15 and x19 and x18 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      elsif ( x65 and not x21 and x22 and x23 and not x15 and x19 and not x18 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s295;

      elsif ( x65 and not x21 and x22 and x23 and not x15 and not x19 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      elsif ( x65 and not x21 and x22 and not x23 and x11 and x18 and x15 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x65 and not x21 and x22 and not x23 and x11 and x18 and not x15 ) = '1' then
         y15 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s227;

      elsif ( x65 and not x21 and x22 and not x23 and x11 and not x18 and x19 and x15 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s247;

      elsif ( x65 and not x21 and x22 and not x23 and x11 and not x18 and x19 and not x15 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x65 and not x21 and x22 and not x23 and x11 and not x18 and not x19 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s231;

      elsif ( x65 and not x21 and x22 and not x23 and not x11 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x65 and not x21 and not x22 and x23 and x16 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      elsif ( x65 and not x21 and not x22 and x23 and not x16 and x20 and x19 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      elsif ( x65 and not x21 and not x22 and x23 and not x16 and x20 and not x19 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and not x22 and x23 and not x16 and x20 and not x19 and x9 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and not x22 and x23 and not x16 and x20 and not x19 and x9 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x22 and x23 and not x16 and x20 and not x19 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x22 and x23 and not x16 and not x20 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      elsif ( x65 and not x21 and not x22 and not x23 and x15 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      elsif ( x65 and not x21 and not x22 and not x23 and not x15 and x19 and x18 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      elsif ( x65 and not x21 and not x22 and not x23 and not x15 and x19 and not x18 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s295;

      elsif ( x65 and not x21 and not x22 and not x23 and not x15 and not x19 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      elsif ( not x65 and x24 and x16 and x26 and x11 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s171;

      elsif ( not x65 and x24 and x16 and x26 and not x11 and x7 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and x24 and x16 and x26 and not x11 and not x7 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s171;

      elsif ( not x65 and x24 and x16 and not x26 and x6 and x11 and x12 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s296;

      elsif ( not x65 and x24 and x16 and not x26 and x6 and x11 and not x12 and x13 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s297;

      elsif ( not x65 and x24 and x16 and not x26 and x6 and x11 and not x12 and not x13 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s160;

      elsif ( not x65 and x24 and x16 and not x26 and x6 and not x11 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and x24 and x16 and not x26 and not x6 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x65 and x24 and not x16 and x26 and x7 and x17 and x13 and x11 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and x24 and not x16 and x26 and x7 and x17 and x13 and not x11 and x12 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( not x65 and x24 and not x16 and x26 and x7 and x17 and x13 and not x11 and not x12 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and x24 and not x16 and x26 and x7 and x17 and not x13 and x11 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s183;

      elsif ( not x65 and x24 and not x16 and x26 and x7 and x17 and not x13 and not x11 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and x24 and not x16 and x26 and x7 and not x17 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x65 and x24 and not x16 and x26 and not x7 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s171;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and x13 and x11 and x9 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and x13 and x11 and not x9 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and x13 and x11 and not x9 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and x13 and x11 and not x9 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and x13 and x11 and not x9 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and x13 and not x11 and x7 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and x13 and not x11 and not x7 and x12 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and x13 and not x11 and not x7 and not x12 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and x13 and not x11 and not x7 and not x12 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and x13 and not x11 and not x7 and not x12 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and x13 and not x11 and not x7 and not x12 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and not x13 and x11 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and not x13 and not x11 and x12 and x10 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and not x13 and not x11 and x12 and not x10 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and not x13 and not x11 and x12 and not x10 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and not x13 and not x11 and x12 and not x10 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and not x13 and not x11 and x12 and not x10 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and not x13 and not x11 and not x12 and x8 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and not x13 and not x11 and not x12 and not x8 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and not x13 and not x11 and not x12 and not x8 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and not x13 and not x11 and not x12 and not x8 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x24 and not x16 and not x26 and x17 and not x13 and not x11 and not x12 and not x8 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x24 and not x16 and not x26 and not x17 and x6 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x24 and not x16 and not x26 and not x17 and not x6 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x65 and not x24 and x25 and x26 and x1 ) = '1' then
         y8 <= '1' ;
         y17 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s164;

      elsif ( not x65 and not x24 and x25 and x26 and not x1 and x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x24 and x25 and x26 and not x1 and not x18 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x65 and not x24 and x25 and not x26 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( not x65 and not x24 and x25 and not x26 and not x2 and x18 and x15 and x10 and x11 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s187;

      elsif ( not x65 and not x24 and x25 and not x26 and not x2 and x18 and x15 and x10 and not x11 and x12 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s185;

      elsif ( not x65 and not x24 and x25 and not x26 and not x2 and x18 and x15 and x10 and not x11 and not x12 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s160;

      elsif ( not x65 and not x24 and x25 and not x26 and not x2 and x18 and x15 and not x10 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s50;

      elsif ( not x65 and not x24 and x25 and not x26 and not x2 and x18 and not x15 and x16 and x10 and x12 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( not x65 and not x24 and x25 and not x26 and not x2 and x18 and not x15 and x16 and x10 and not x12 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and not x24 and x25 and not x26 and not x2 and x18 and not x15 and x16 and not x10 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( not x65 and not x24 and x25 and not x26 and not x2 and x18 and not x15 and not x16 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x65 and not x24 and x25 and not x26 and not x2 and not x18 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      else
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      end if;

   when s55 =>
      if ( x65 and x21 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x22 and x23 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x22 and not x23 and x15 and x9 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x21 and x22 and not x23 and x15 and not x9 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x65 and not x21 and x22 and not x23 and not x15 and x16 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and x22 and not x23 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s205;

      elsif ( x65 and not x21 and not x22 and x23 and x17 and x15 and x9 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( x65 and not x21 and not x22 and x23 and x17 and x15 and not x9 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x65 and not x21 and not x22 and x23 and x17 and not x15 and x16 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and not x22 and x23 and x17 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s205;

      elsif ( x65 and not x21 and not x22 and x23 and not x17 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x21 and not x22 and not x23 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( not x65 and x66 and x63 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x63 and x62 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x63 and not x62 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s298;

      elsif ( not x65 and not x66 and x25 ) = '1' then
         y2 <= '1' ;
         y14 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s56 =>
      if ( x66 and x65 and x67 and x22 and x17 and x18 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and x65 and x67 and x22 and x17 and not x18 and x19 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and x65 and x67 and x22 and x17 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and x67 and x22 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and x67 and not x22 and x18 and x13 and x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x66 and x65 and x67 and not x22 and x18 and x13 and not x23 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and x67 and not x22 and x18 and not x13 and x12 and x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x66 and x65 and x67 and not x22 and x18 and not x13 and x12 and not x23 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and x67 and not x22 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and x67 and not x22 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x67 and x21 and x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and x3 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x3 and x18 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s299;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x3 and not x18 and x15 and x10 and x11 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s192;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x3 and not x18 and x15 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s193;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x3 and not x18 and x15 and x10 and not x11 and not x12 ) = '1' then
         y1 <= '1' ;
         y8 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s192;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x3 and not x18 and x15 and not x10 and x12 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s300;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x3 and not x18 and x15 and not x10 and not x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s192;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x3 and not x18 and not x15 and x16 and x10 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x3 and not x18 and not x15 and x16 and x10 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x3 and not x18 and not x15 and x16 and x10 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x3 and not x18 and not x15 and x16 and x10 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x3 and not x18 and not x15 and x16 and not x10 and x12 and x11 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s199;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x3 and not x18 and not x15 and x16 and not x10 and x12 and not x11 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x3 and not x18 and not x15 and x16 and not x10 and x12 and not x11 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x3 and not x18 and not x15 and x16 and not x10 and x12 and not x11 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x3 and not x18 and not x15 and x16 and not x10 and x12 and not x11 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x3 and not x18 and not x15 and x16 and not x10 and not x12 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x3 and not x18 and not x15 and x16 and not x10 and not x12 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x3 and not x18 and not x15 and x16 and not x10 and not x12 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x3 and not x18 and not x15 and x16 and not x10 and not x12 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and not x67 and x21 and not x20 and not x3 and not x18 and not x15 and not x16 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s201;

      elsif ( x66 and x65 and not x67 and not x21 and x15 and x10 and x11 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x66 and x65 and not x67 and not x21 and x15 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s301;

      elsif ( x66 and x65 and not x67 and not x21 and x15 and x10 and not x11 and not x12 ) = '1' then
         y8 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s195;

      elsif ( x66 and x65 and not x67 and not x21 and x15 and not x10 and x12 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      elsif ( x66 and x65 and not x67 and not x21 and x15 and not x10 and not x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s192;

      elsif ( x66 and x65 and not x67 and not x21 and not x15 and x16 and x10 and x12 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s259;

      elsif ( x66 and x65 and not x67 and not x21 and not x15 and x16 and x10 and not x12 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s302;

      elsif ( x66 and x65 and not x67 and not x21 and not x15 and x16 and not x10 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s259;

      elsif ( x66 and x65 and not x67 and not x21 and not x15 and not x16 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s303;

      elsif ( x66 and not x65 and x21 and x15 and x4 and x10 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x66 and not x65 and x21 and x15 and x4 and not x10 and x12 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x66 and not x65 and x21 and x15 and x4 and not x10 and not x12 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      elsif ( x66 and not x65 and x21 and x15 and not x4 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( x66 and not x65 and x21 and not x15 and x16 and x10 and x12 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( x66 and not x65 and x21 and not x15 and x16 and x10 and not x12 ) = '1' then
         y4 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s304;

      elsif ( x66 and not x65 and x21 and not x15 and x16 and not x10 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( x66 and not x65 and x21 and not x15 and not x16 and x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( x66 and not x65 and x21 and not x15 and not x16 and not x4 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( x66 and not x65 and not x21 and x22 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( x66 and not x65 and not x21 and not x22 and x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s250;

      elsif ( x66 and not x65 and not x21 and not x22 and not x23 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s85;

      elsif ( not x66 and x65 and x68 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x66 and x65 and x68 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x66 and x65 and x68 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and x68 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x68 and x21 and x18 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x66 and x65 and not x68 and x21 and not x18 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and not x68 and x21 and not x18 and x19 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and not x68 and x21 and not x18 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x68 and x21 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and x15 and x16 and x7 and x9 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and x15 and x16 and x7 and not x9 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and x15 and x16 and not x7 and x8 and x9 ) = '1' then
         y24 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s157;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and x15 and x16 and not x7 and x8 and not x9 ) = '1' then
         y26 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s158;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and x15 and x16 and not x7 and not x8 and x9 and x13 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s191;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and x15 and x16 and not x7 and not x8 and x9 and not x13 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and x15 and x16 and not x7 and not x8 and x9 and not x13 and not x19 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and x15 and x16 and not x7 and not x8 and x9 and not x13 and not x19 and x17 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and x15 and x16 and not x7 and not x8 and x9 and not x13 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and x15 and x16 and not x7 and not x8 and not x9 and x14 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s191;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and x15 and x16 and not x7 and not x8 and not x9 and not x14 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and x15 and x16 and not x7 and not x8 and not x9 and not x14 and not x19 and x17 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and x15 and x16 and not x7 and not x8 and not x9 and not x14 and not x19 and x17 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and x15 and x16 and not x7 and not x8 and not x9 and not x14 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and x15 and not x16 and x7 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s147;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and x15 and not x16 and not x7 and x8 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s147;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and x15 and not x16 and not x7 and not x8 and x4 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s22;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and x15 and not x16 and not x7 and not x8 and not x4 and x5 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and x15 and not x16 and not x7 and not x8 and not x4 and not x5 and x9 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and x15 and not x16 and not x7 and not x8 and not x4 and not x5 and not x9 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and x4 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s22;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and x16 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and x16 and x9 and not x10 and x8 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and x16 and x9 and not x10 and not x8 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and x16 and x9 and not x10 and not x8 and not x19 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and x16 and x9 and not x10 and not x8 and not x19 and x17 and not x14 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and x16 and x9 and not x10 and not x8 and not x19 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and x16 and x9 and not x10 and not x8 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and x16 and not x9 and x8 and x12 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and x16 and not x9 and x8 and not x12 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and x16 and not x9 and x8 and not x12 and not x19 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and x16 and not x9 and x8 and not x12 and not x19 and x17 and not x14 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and x16 and not x9 and x8 and not x12 and not x19 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and x16 and not x9 and x8 and not x12 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and x16 and not x9 and not x8 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and x16 and not x9 and not x8 and not x11 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and x16 and not x9 and not x8 and not x11 and not x19 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and x16 and not x9 and not x8 and not x11 and not x19 and x17 and not x14 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and x16 and not x9 and not x8 and not x11 and not x19 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and x16 and not x9 and not x8 and not x11 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and not x16 and x5 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and x65 and not x68 and not x21 and x22 and not x15 and not x4 and not x16 and not x5 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s212;

      elsif ( not x66 and x65 and not x68 and not x21 and not x22 and x2 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( not x66 and x65 and not x68 and not x21 and not x22 and not x2 and x17 and x15 and x9 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and x65 and not x68 and not x21 and not x22 and not x2 and x17 and x15 and not x9 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x66 and x65 and not x68 and not x21 and not x22 and not x2 and x17 and not x15 and x16 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x66 and x65 and not x68 and not x21 and not x22 and not x2 and x17 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s205;

      elsif ( not x66 and x65 and not x68 and not x21 and not x22 and not x2 and not x17 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( not x66 and not x65 and x20 and x15 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s198;

      elsif ( not x66 and not x65 and x20 and not x15 ) = '1' then
         y7 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s211;

      elsif ( not x66 and not x65 and not x20 and x21 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x66 and not x65 and not x20 and x21 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x66 and not x65 and not x20 and x21 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x20 and x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x20 and not x21 and x17 and x13 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x66 and not x65 and not x20 and not x21 and x17 and not x13 and x12 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x66 and not x65 and not x20 and not x21 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s57 =>
      if ( x21 ) = '1' then
         current_group15m <= s1;

      else
         y2 <= '1' ;
         current_group15m <= s56;

      end if;

   when s58 =>
      if ( x68 and x21 and x20 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s191;

      elsif ( x68 and x21 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x68 and not x21 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s59;

      else
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      end if;

   when s59 =>
      if ( x65 and x21 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s60;

      elsif ( not x65 and x20 and x18 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x20 and x18 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x20 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x20 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x20 and x21 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x20 and x21 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x20 and x21 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x20 and x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x20 and not x21 and x17 and x13 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x65 and not x20 and not x21 and x17 and not x13 and x12 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x65 and not x20 and not x21 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s60 =>
      if ( x21 and x20 and x2 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s306;

      elsif ( x21 and x20 and not x2 and x18 and x15 and x10 and x11 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s192;

      elsif ( x21 and x20 and not x2 and x18 and x15 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s193;

      elsif ( x21 and x20 and not x2 and x18 and x15 and x10 and not x11 and not x12 ) = '1' then
         y1 <= '1' ;
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s194;

      elsif ( x21 and x20 and not x2 and x18 and x15 and not x10 and x12 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s300;

      elsif ( x21 and x20 and not x2 and x18 and x15 and not x10 and not x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s192;

      elsif ( x21 and x20 and not x2 and x18 and not x15 and x16 and x10 and x12 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s259;

      elsif ( x21 and x20 and not x2 and x18 and not x15 and x16 and x10 and not x12 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( x21 and x20 and not x2 and x18 and not x15 and x16 and not x10 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s259;

      elsif ( x21 and x20 and not x2 and x18 and not x15 and not x16 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x21 and x20 and not x2 and not x18 ) = '1' then
         y4 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s307;

      elsif ( x21 and not x20 ) = '1' then
         y4 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s307;

      else
         y4 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s307;

      end if;

   when s61 =>
      if ( x21 and x20 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x20 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x20 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x20 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x20 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x20 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x20 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x20 and not x19 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s62 =>
      if ( x65 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( not x65 and x66 and x21 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s232;

      elsif ( not x65 and x66 and not x21 and x22 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s262;

      elsif ( not x65 and x66 and not x21 and not x22 and x10 and x16 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s219;

      elsif ( not x65 and x66 and not x21 and not x22 and x10 and not x16 and x17 and x15 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s219;

      elsif ( not x65 and x66 and not x21 and not x22 and x10 and not x16 and x17 and not x15 and x3 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s214;

      elsif ( not x65 and x66 and not x21 and not x22 and x10 and not x16 and x17 and not x15 and not x3 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s308;

      elsif ( not x65 and x66 and not x21 and not x22 and x10 and not x16 and not x17 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s219;

      elsif ( not x65 and x66 and not x21 and not x22 and not x10 and x16 and x15 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s309;

      elsif ( not x65 and x66 and not x21 and not x22 and not x10 and x16 and not x15 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s310;

      elsif ( not x65 and x66 and not x21 and not x22 and not x10 and not x16 and x17 and x15 and x14 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s217;

      elsif ( not x65 and x66 and not x21 and not x22 and not x10 and not x16 and x17 and x15 and not x14 ) = '1' then
         y2 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s79;

      elsif ( not x65 and x66 and not x21 and not x22 and not x10 and not x16 and x17 and not x15 ) = '1' then
         y2 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s79;

      elsif ( not x65 and x66 and not x21 and not x22 and not x10 and not x16 and not x17 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s311;

      elsif ( not x65 and not x66 and x68 and x21 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x66 and x68 and not x21 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( not x65 and not x66 and not x68 and x22 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and not x66 and not x68 and not x22 and x21 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      else
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      end if;

   when s63 =>
      if ( x61 and x60 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x61 and not x60 and x62 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x61 and not x60 and not x62 ) = '1' then
         current_group15m <= s40;

      elsif ( not x61 and x60 ) = '1' then
         current_group15m <= s40;

      elsif ( not x61 and not x60 and x62 ) = '1' then
         current_group15m <= s40;

      else
         current_group15m <= s1;

      end if;

   when s64 =>
      if ( x60 and x61 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s286;

      elsif ( x60 and not x61 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s154;

      elsif ( not x60 and x62 and x61 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x60 and x62 and x61 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x60 and x62 and x61 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( not x60 and x62 and x61 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x60 and x62 and not x61 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s312;

      else
         y3 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s154;

      end if;

   when s65 =>
      if ( x65 and x66 and x61 and x60 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( x65 and x66 and x61 and not x60 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s258;

      elsif ( x65 and x66 and not x61 and x60 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s258;

      elsif ( x65 and x66 and not x61 and not x60 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and not x66 ) = '1' then
         y15 <= '1' ;
         y21 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s313;

      elsif ( not x65 and x66 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and not x66 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s65;

      else
         current_group15m <= s1;

      end if;

   when s66 =>
      if ( x61 and x60 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s68;

      elsif ( x61 and not x60 and x62 ) = '1' then
         current_group15m <= s1;

      elsif ( x61 and not x60 and not x62 ) = '1' then
         current_group15m <= s39;

      elsif ( not x61 and x60 ) = '1' then
         current_group15m <= s39;

      elsif ( not x61 and not x60 and x62 and x4 and x15 and x12 and x7 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s314;

      elsif ( not x61 and not x60 and x62 and x4 and x15 and x12 and not x7 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s315;

      elsif ( not x61 and not x60 and x62 and x4 and x15 and not x12 and x7 ) = '1' then
         current_group15m <= s316;

      elsif ( not x61 and not x60 and x62 and x4 and x15 and not x12 and not x7 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x61 and not x60 and x62 and x4 and not x15 and x16 and x7 and x12 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s315;

      elsif ( not x61 and not x60 and x62 and x4 and not x15 and x16 and x7 and not x12 ) = '1' then
         current_group15m <= s316;

      elsif ( not x61 and not x60 and x62 and x4 and not x15 and x16 and not x7 ) = '1' then
         current_group15m <= s316;

      elsif ( not x61 and not x60 and x62 and x4 and not x15 and not x16 and x7 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s252;

      elsif ( not x61 and not x60 and x62 and x4 and not x15 and not x16 and not x7 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( not x61 and not x60 and x62 and not x4 ) = '1' then
         current_group15m <= s316;

      elsif ( not x61 and not x60 and not x62 and x15 and x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( not x61 and not x60 and not x62 and x15 and not x7 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x61 and not x60 and not x62 and x15 and not x7 and not x11 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s254;

      elsif ( not x61 and not x60 and not x62 and not x15 and x16 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      end if;

   when s67 =>
      if ( x65 and x60 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s68;

      elsif ( x65 and not x60 and x61 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x60 and not x61 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s118;

      elsif ( not x65 and x21 and x3 ) = '1' then
         y13 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s141;

      elsif ( not x65 and x21 and not x3 and x20 and x16 and x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s113;

      elsif ( not x65 and x21 and not x3 and x20 and x16 and not x10 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and x21 and not x3 and x20 and not x16 and x17 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x65 and x21 and not x3 and x20 and not x16 and not x17 ) = '1' then
         y5 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s115;

      elsif ( not x65 and x21 and not x3 and not x20 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s317;

      elsif ( not x65 and not x21 and x20 and x15 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( not x65 and not x21 and x20 and not x15 and x14 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( not x65 and not x21 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s68 =>
      if ( x60 and x61 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x60 and x61 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x60 and x61 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x60 and x61 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x60 and not x61 and x15 and x5 and x12 and x7 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s318;

      elsif ( x60 and not x61 and x15 and x5 and x12 and not x7 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s318;

      elsif ( x60 and not x61 and x15 and x5 and not x12 and x7 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( x60 and not x61 and x15 and x5 and not x12 and not x7 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s254;

      elsif ( x60 and not x61 and x15 and not x5 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( x60 and not x61 and not x15 and x16 and x7 and x12 and x5 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s75;

      elsif ( x60 and not x61 and not x15 and x16 and x7 and x12 and not x5 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( x60 and not x61 and not x15 and x16 and x7 and not x12 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( x60 and not x61 and not x15 and x16 and not x7 and x12 and x9 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( x60 and not x61 and not x15 and x16 and not x7 and x12 and not x9 and x11 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( x60 and not x61 and not x15 and x16 and not x7 and x12 and not x9 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x60 and not x61 and not x15 and x16 and not x7 and not x12 and x11 and x10 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( x60 and not x61 and not x15 and x16 and not x7 and not x12 and x11 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x60 and not x61 and not x15 and x16 and not x7 and not x12 and not x11 and x8 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( x60 and not x61 and not x15 and x16 and not x7 and not x12 and not x11 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x60 and not x61 and not x15 and not x16 and x5 and x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s253;

      elsif ( x60 and not x61 and not x15 and not x16 and x5 and not x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x60 and not x61 and not x15 and not x16 and not x5 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( not x60 and x61 and x62 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s286;

      elsif ( not x60 and x61 and not x62 and x15 and x5 and x12 and x7 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s318;

      elsif ( not x60 and x61 and not x62 and x15 and x5 and x12 and not x7 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s318;

      elsif ( not x60 and x61 and not x62 and x15 and x5 and not x12 and x7 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( not x60 and x61 and not x62 and x15 and x5 and not x12 and not x7 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s254;

      elsif ( not x60 and x61 and not x62 and x15 and not x5 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( not x60 and x61 and not x62 and not x15 and x16 and x7 and x12 and x5 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s75;

      elsif ( not x60 and x61 and not x62 and not x15 and x16 and x7 and x12 and not x5 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( not x60 and x61 and not x62 and not x15 and x16 and x7 and not x12 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( not x60 and x61 and not x62 and not x15 and x16 and not x7 and x12 and x9 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( not x60 and x61 and not x62 and not x15 and x16 and not x7 and x12 and not x9 and x11 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( not x60 and x61 and not x62 and not x15 and x16 and not x7 and x12 and not x9 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x60 and x61 and not x62 and not x15 and x16 and not x7 and not x12 and x11 and x10 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( not x60 and x61 and not x62 and not x15 and x16 and not x7 and not x12 and x11 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x60 and x61 and not x62 and not x15 and x16 and not x7 and not x12 and not x11 and x8 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( not x60 and x61 and not x62 and not x15 and x16 and not x7 and not x12 and not x11 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x60 and x61 and not x62 and not x15 and not x16 and x5 and x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s253;

      elsif ( not x60 and x61 and not x62 and not x15 and not x16 and x5 and not x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( not x60 and x61 and not x62 and not x15 and not x16 and not x5 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( not x60 and not x61 and x62 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      else
         y3 <= '1' ;
         current_group15m <= s320;

      end if;

   when s69 =>
      if ( x65 and x60 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s68;

      elsif ( x65 and not x60 and x61 ) = '1' then
         y2 <= '1' ;
         y19 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s321;

      elsif ( x65 and not x60 and not x61 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      else
         y14 <= '1' ;
         current_group15m <= s286;

      end if;

   when s70 =>
      if ( x60 ) = '1' then
         current_group15m <= s316;

      elsif ( not x60 and x61 ) = '1' then
         current_group15m <= s316;

      else
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      end if;

   when s71 =>
      if ( x60 ) = '1' then
         current_group15m <= s316;

      elsif ( not x60 and x61 ) = '1' then
         current_group15m <= s316;

      elsif ( not x60 and not x61 and x17 and x62 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s255;

      elsif ( not x60 and not x61 and x17 and not x62 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s63;

      else
         current_group15m <= s39;

      end if;

   when s72 =>
      if ( x65 and x66 and x61 and x60 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x61 and not x60 and x62 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x66 and x61 and not x60 and x62 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x66 and x61 and not x60 and x62 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x61 and not x60 and x62 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x61 and not x60 and not x62 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( x65 and x66 and not x61 and x60 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( x65 and x66 and not x61 and not x60 and x62 and x7 and x15 and x12 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s292;

      elsif ( x65 and x66 and not x61 and not x60 and x62 and x7 and x15 and not x12 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s63;

      elsif ( x65 and x66 and not x61 and not x60 and x62 and x7 and not x15 and x16 and x12 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s290;

      elsif ( x65 and x66 and not x61 and not x60 and x62 and x7 and not x15 and x16 and not x12 and x2 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         y10 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s322;

      elsif ( x65 and x66 and not x61 and not x60 and x62 and x7 and not x15 and x16 and not x12 and not x2 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s262;

      elsif ( x65 and x66 and not x61 and not x60 and x62 and x7 and not x15 and not x16 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and x66 and not x61 and not x60 and x62 and not x7 and x15 and x12 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s290;

      elsif ( x65 and x66 and not x61 and not x60 and x62 and not x7 and x15 and not x12 ) = '1' then
         y2 <= '1' ;
         y10 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s263;

      elsif ( x65 and x66 and not x61 and not x60 and x62 and not x7 and not x15 and x16 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x65 and x66 and not x61 and not x60 and x62 and not x7 and not x15 and not x16 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x66 and not x61 and not x60 and not x62 and x4 and x15 and x7 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and x66 and not x61 and not x60 and not x62 and x4 and x15 and not x7 and x11 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and x66 and not x61 and not x60 and not x62 and x4 and x15 and not x7 and not x11 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x66 and not x61 and not x60 and not x62 and x4 and not x15 and x16 ) = '1' then
         current_group15m <= s70;

      elsif ( x65 and x66 and not x61 and not x60 and not x62 and x4 and not x15 and not x16 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( x65 and x66 and not x61 and not x60 and not x62 and not x4 ) = '1' then
         current_group15m <= s70;

      elsif ( x65 and not x66 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( not x65 and x21 and x66 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x21 and x66 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x21 and x66 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and x66 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and not x66 and x19 and x20 and x12 and x17 ) = '1' then
         y8 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s266;

      elsif ( not x65 and x21 and not x66 and x19 and x20 and x12 and not x17 ) = '1' then
         y8 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s267;

      elsif ( not x65 and x21 and not x66 and x19 and x20 and not x12 and x16 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x65 and x21 and not x66 and x19 and x20 and not x12 and not x16 and x17 and x5 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s181;

      elsif ( not x65 and x21 and not x66 and x19 and x20 and not x12 and not x16 and x17 and not x5 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s246;

      elsif ( not x65 and x21 and not x66 and x19 and x20 and not x12 and not x16 and not x17 and x4 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s181;

      elsif ( not x65 and x21 and not x66 and x19 and x20 and not x12 and not x16 and not x17 and not x4 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s246;

      elsif ( not x65 and x21 and not x66 and x19 and not x20 and x16 and x12 ) = '1' then
         y8 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s323;

      elsif ( not x65 and x21 and not x66 and x19 and not x20 and x16 and not x12 and x17 ) = '1' then
         y8 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s82;

      elsif ( not x65 and x21 and not x66 and x19 and not x20 and x16 and not x12 and not x17 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x65 and x21 and not x66 and x19 and not x20 and not x16 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x65 and x21 and not x66 and not x19 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x65 and not x21 and x66 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      else
         y3 <= '1' ;
         current_group15m <= s89;

      end if;

   when s73 =>
      if ( x60 and x15 and x12 and x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x60 and x15 and x12 and not x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s250;

      elsif ( x60 and x15 and not x12 and x7 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x60 and x15 and not x12 and not x7 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s262;

      elsif ( x60 and not x15 and x16 and x7 and x12 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s251;

      elsif ( x60 and not x15 and x16 and x7 and not x12 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x60 and not x15 and x16 and not x7 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x60 and not x15 and not x16 and x7 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s318;

      elsif ( x60 and not x15 and not x16 and not x7 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s74;

      elsif ( not x60 and x61 and x15 and x12 and x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( not x60 and x61 and x15 and x12 and not x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s250;

      elsif ( not x60 and x61 and x15 and not x12 and x7 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( not x60 and x61 and x15 and not x12 and not x7 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s262;

      elsif ( not x60 and x61 and not x15 and x16 and x7 and x12 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s251;

      elsif ( not x60 and x61 and not x15 and x16 and x7 and not x12 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x60 and x61 and not x15 and x16 and not x7 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x60 and x61 and not x15 and not x16 and x7 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s318;

      elsif ( not x60 and x61 and not x15 and not x16 and not x7 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s74;

      elsif ( not x60 and not x61 and x62 ) = '1' then
         y4 <= '1' ;
         y13 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s64;

      else
         y25 <= '1' ;
         current_group15m <= s324;

      end if;

   when s74 =>
      if ( x61 and x60 and x7 and x15 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x61 and x60 and x7 and not x15 and x16 and x12 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s251;

      elsif ( x61 and x60 and x7 and not x15 and x16 and not x12 and x3 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s258;

      elsif ( x61 and x60 and x7 and not x15 and x16 and not x12 and not x3 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( x61 and x60 and x7 and not x15 and not x16 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s253;

      elsif ( x61 and x60 and not x7 and x15 and x12 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s250;

      elsif ( x61 and x60 and not x7 and x15 and not x12 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( x61 and x60 and not x7 and not x15 and x16 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x61 and x60 and not x7 and not x15 and not x16 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x61 and not x60 and x62 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x61 and not x60 and not x62 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      elsif ( not x61 and x60 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      elsif ( not x61 and not x60 and x62 and x16 and x15 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( not x61 and not x60 and x62 and x16 and not x15 and x11 and x12 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      elsif ( not x61 and not x60 and x62 and x16 and not x15 and x11 and not x12 and x7 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      elsif ( not x61 and not x60 and x62 and x16 and not x15 and x11 and not x12 and not x7 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x61 and not x60 and x62 and x16 and not x15 and not x11 and x7 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      elsif ( not x61 and not x60 and x62 and x16 and not x15 and not x11 and not x7 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x61 and not x60 and x62 and not x16 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      elsif ( not x61 and not x60 and not x62 and x15 and x16 and x9 and x11 ) = '1' then
         current_group15m <= s40;

      elsif ( not x61 and not x60 and not x62 and x15 and x16 and x9 and not x11 and x7 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x61 and not x60 and not x62 and x15 and x16 and x9 and not x11 and not x7 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         y10 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s261;

      elsif ( not x61 and not x60 and not x62 and x15 and x16 and not x9 and x11 and x7 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s262;

      elsif ( not x61 and not x60 and not x62 and x15 and x16 and not x9 and x11 and not x7 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s260;

      elsif ( not x61 and not x60 and not x62 and x15 and x16 and not x9 and not x11 and x7 and x14 ) = '1' then
         current_group15m <= s316;

      elsif ( not x61 and not x60 and not x62 and x15 and x16 and not x9 and not x11 and x7 and not x14 ) = '1' then
         current_group15m <= s40;

      elsif ( not x61 and not x60 and not x62 and x15 and x16 and not x9 and not x11 and not x7 and x13 ) = '1' then
         current_group15m <= s316;

      elsif ( not x61 and not x60 and not x62 and x15 and x16 and not x9 and not x11 and not x7 and not x13 ) = '1' then
         current_group15m <= s40;

      elsif ( not x61 and not x60 and not x62 and x15 and not x16 and x9 and x3 ) = '1' then
         current_group15m <= s40;

      elsif ( not x61 and not x60 and not x62 and x15 and not x16 and x9 and not x3 and x7 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s325;

      elsif ( not x61 and not x60 and not x62 and x15 and not x16 and x9 and not x3 and not x7 and x11 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s325;

      elsif ( not x61 and not x60 and not x62 and x15 and not x16 and x9 and not x3 and not x7 and not x11 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( not x61 and not x60 and not x62 and x15 and not x16 and not x9 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s69;

      elsif ( not x61 and not x60 and not x62 and x15 and not x16 and not x9 and not x3 and x5 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      elsif ( not x61 and not x60 and not x62 and x15 and not x16 and not x9 and not x3 and not x5 and x7 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s326;

      elsif ( not x61 and not x60 and not x62 and x15 and not x16 and not x9 and not x3 and not x5 and not x7 and x11 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( not x61 and not x60 and not x62 and x15 and not x16 and not x9 and not x3 and not x5 and not x7 and not x11 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( not x61 and not x60 and not x62 and not x15 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s69;

      elsif ( not x61 and not x60 and not x62 and not x15 and not x3 and x16 and x11 and x9 ) = '1' then
         current_group15m <= s40;

      elsif ( not x61 and not x60 and not x62 and not x15 and not x3 and x16 and x11 and not x9 and x7 and x5 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      elsif ( not x61 and not x60 and not x62 and not x15 and not x3 and x16 and x11 and not x9 and x7 and not x5 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s326;

      elsif ( not x61 and not x60 and not x62 and not x15 and not x3 and x16 and x11 and not x9 and not x7 and x5 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s131;

      elsif ( not x61 and not x60 and not x62 and not x15 and not x3 and x16 and x11 and not x9 and not x7 and not x5 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s67;

      elsif ( not x61 and not x60 and not x62 and not x15 and not x3 and x16 and not x11 and x7 and x9 and x5 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s256;

      elsif ( not x61 and not x60 and not x62 and not x15 and not x3 and x16 and not x11 and x7 and x9 and not x5 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s252;

      elsif ( not x61 and not x60 and not x62 and not x15 and not x3 and x16 and not x11 and x7 and not x9 and x8 and x5 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s256;

      elsif ( not x61 and not x60 and not x62 and not x15 and not x3 and x16 and not x11 and x7 and not x9 and x8 and not x5 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s252;

      elsif ( not x61 and not x60 and not x62 and not x15 and not x3 and x16 and not x11 and x7 and not x9 and not x8 ) = '1' then
         current_group15m <= s40;

      elsif ( not x61 and not x60 and not x62 and not x15 and not x3 and x16 and not x11 and not x7 and x9 and x10 and x5 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s256;

      elsif ( not x61 and not x60 and not x62 and not x15 and not x3 and x16 and not x11 and not x7 and x9 and x10 and not x5 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s252;

      elsif ( not x61 and not x60 and not x62 and not x15 and not x3 and x16 and not x11 and not x7 and x9 and not x10 ) = '1' then
         current_group15m <= s40;

      elsif ( not x61 and not x60 and not x62 and not x15 and not x3 and x16 and not x11 and not x7 and not x9 and x12 and x5 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s256;

      elsif ( not x61 and not x60 and not x62 and not x15 and not x3 and x16 and not x11 and not x7 and not x9 and x12 and not x5 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s252;

      elsif ( not x61 and not x60 and not x62 and not x15 and not x3 and x16 and not x11 and not x7 and not x9 and not x12 ) = '1' then
         current_group15m <= s40;

      elsif ( not x61 and not x60 and not x62 and not x15 and not x3 and not x16 and x5 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      else
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s68;

      end if;

   when s75 =>
      if ( x65 and x60 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      elsif ( x65 and not x60 and x61 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      elsif ( x65 and not x60 and not x61 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( not x65 and x21 and x16 and x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s113;

      elsif ( not x65 and x21 and x16 and not x10 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and x21 and not x16 and x17 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x65 and x21 and not x16 and not x17 ) = '1' then
         y5 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s115;

      elsif ( not x65 and not x21 and x3 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s14;

      elsif ( not x65 and not x21 and not x3 and x19 and x16 and x10 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s67;

      elsif ( not x65 and not x21 and not x3 and x19 and x16 and not x10 ) = '1' then
         y5 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s113;

      elsif ( not x65 and not x21 and not x3 and x19 and not x16 and x17 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x65 and not x21 and not x3 and x19 and not x16 and not x17 ) = '1' then
         y5 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s115;

      else
         y13 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s141;

      end if;

   when s76 =>
      if ( x65 and x61 and x60 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x61 and x60 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x61 and x60 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x61 and x60 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x61 and not x60 and x62 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and x16 and x7 and x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and x16 and x7 and not x12 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and x16 and not x7 and x12 and x14 and x11 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s260;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and x16 and not x7 and x12 and x14 and not x11 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and x16 and not x7 and x12 and not x14 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and x16 and not x7 and x12 and not x14 and x18 and not x13 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and x16 and not x7 and x12 and not x14 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and x16 and not x7 and not x12 and x13 and x11 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         y10 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s261;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and x16 and not x7 and not x12 and x13 and not x11 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and x16 and not x7 and not x12 and not x13 and x18 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and x16 and not x7 and not x12 and not x13 and x18 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and x16 and not x7 and not x12 and not x13 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and not x16 and x11 and x7 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s327;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and not x16 and x11 and not x7 and x12 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and not x16 and x11 and not x7 and not x12 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s318;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and not x16 and not x11 and x4 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s328;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and not x16 and not x11 and not x4 and x2 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and not x16 and not x11 and not x4 and not x2 and x12 and x7 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s329;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and not x16 and not x11 and not x4 and not x2 and x12 and not x7 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s318;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and not x16 and not x11 and not x4 and not x2 and not x12 and x7 ) = '1' then
         y2 <= '1' ;
         y10 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s263;

      elsif ( x65 and x61 and not x60 and not x62 and x15 and not x16 and not x11 and not x4 and not x2 and not x12 and not x7 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x61 and not x60 and not x62 and not x15 and x4 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s328;

      elsif ( x65 and x61 and not x60 and not x62 and not x15 and not x4 and x16 and x7 and x12 and x2 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x61 and not x60 and not x62 and not x15 and not x4 and x16 and x7 and x12 and not x2 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s318;

      elsif ( x65 and x61 and not x60 and not x62 and not x15 and not x4 and x16 and x7 and not x12 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s65;

      elsif ( x65 and x61 and not x60 and not x62 and not x15 and not x4 and x16 and not x7 and x12 and x11 and x2 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x61 and not x60 and not x62 and not x15 and not x4 and x16 and not x7 and x12 and x11 and not x2 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and x61 and not x60 and not x62 and not x15 and not x4 and x16 and not x7 and x12 and not x11 and x9 and x2 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x61 and not x60 and not x62 and not x15 and not x4 and x16 and not x7 and x12 and not x11 and x9 and not x2 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and x61 and not x60 and not x62 and not x15 and not x4 and x16 and not x7 and x12 and not x11 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x61 and not x60 and not x62 and not x15 and not x4 and x16 and not x7 and not x12 and x11 and x10 and x2 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x61 and not x60 and not x62 and not x15 and not x4 and x16 and not x7 and not x12 and x11 and x10 and not x2 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and x61 and not x60 and not x62 and not x15 and not x4 and x16 and not x7 and not x12 and x11 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x61 and not x60 and not x62 and not x15 and not x4 and x16 and not x7 and not x12 and not x11 and x8 and x2 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x61 and not x60 and not x62 and not x15 and not x4 and x16 and not x7 and not x12 and not x11 and x8 and not x2 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and x61 and not x60 and not x62 and not x15 and not x4 and x16 and not x7 and not x12 and not x11 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x61 and not x60 and not x62 and not x15 and not x4 and not x16 and x2 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x61 and not x60 and not x62 and not x15 and not x4 and not x16 and not x2 and x7 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s318;

      elsif ( x65 and x61 and not x60 and not x62 and not x15 and not x4 and not x16 and not x2 and not x7 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s191;

      elsif ( x65 and not x61 and x60 and x15 and x16 and x7 and x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( x65 and not x61 and x60 and x15 and x16 and x7 and not x12 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( x65 and not x61 and x60 and x15 and x16 and not x7 and x12 and x14 and x11 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s260;

      elsif ( x65 and not x61 and x60 and x15 and x16 and not x7 and x12 and x14 and not x11 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( x65 and not x61 and x60 and x15 and x16 and not x7 and x12 and not x14 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x61 and x60 and x15 and x16 and not x7 and x12 and not x14 and x18 and not x13 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and not x61 and x60 and x15 and x16 and not x7 and x12 and not x14 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and not x61 and x60 and x15 and x16 and not x7 and not x12 and x13 and x11 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         y10 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s261;

      elsif ( x65 and not x61 and x60 and x15 and x16 and not x7 and not x12 and x13 and not x11 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( x65 and not x61 and x60 and x15 and x16 and not x7 and not x12 and not x13 and x18 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x61 and x60 and x15 and x16 and not x7 and not x12 and not x13 and x18 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and not x61 and x60 and x15 and x16 and not x7 and not x12 and not x13 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and not x61 and x60 and x15 and not x16 and x11 and x7 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s327;

      elsif ( x65 and not x61 and x60 and x15 and not x16 and x11 and not x7 and x12 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( x65 and not x61 and x60 and x15 and not x16 and x11 and not x7 and not x12 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s318;

      elsif ( x65 and not x61 and x60 and x15 and not x16 and not x11 and x4 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s328;

      elsif ( x65 and not x61 and x60 and x15 and not x16 and not x11 and not x4 and x2 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and not x61 and x60 and x15 and not x16 and not x11 and not x4 and not x2 and x12 and x7 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s329;

      elsif ( x65 and not x61 and x60 and x15 and not x16 and not x11 and not x4 and not x2 and x12 and not x7 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s318;

      elsif ( x65 and not x61 and x60 and x15 and not x16 and not x11 and not x4 and not x2 and not x12 and x7 ) = '1' then
         y2 <= '1' ;
         y10 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s263;

      elsif ( x65 and not x61 and x60 and x15 and not x16 and not x11 and not x4 and not x2 and not x12 and not x7 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x61 and x60 and not x15 and x4 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s328;

      elsif ( x65 and not x61 and x60 and not x15 and not x4 and x16 and x7 and x12 and x2 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and not x61 and x60 and not x15 and not x4 and x16 and x7 and x12 and not x2 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s318;

      elsif ( x65 and not x61 and x60 and not x15 and not x4 and x16 and x7 and not x12 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s65;

      elsif ( x65 and not x61 and x60 and not x15 and not x4 and x16 and not x7 and x12 and x11 and x2 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and not x61 and x60 and not x15 and not x4 and x16 and not x7 and x12 and x11 and not x2 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and not x61 and x60 and not x15 and not x4 and x16 and not x7 and x12 and not x11 and x9 and x2 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and not x61 and x60 and not x15 and not x4 and x16 and not x7 and x12 and not x11 and x9 and not x2 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and not x61 and x60 and not x15 and not x4 and x16 and not x7 and x12 and not x11 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x61 and x60 and not x15 and not x4 and x16 and not x7 and not x12 and x11 and x10 and x2 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and not x61 and x60 and not x15 and not x4 and x16 and not x7 and not x12 and x11 and x10 and not x2 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and not x61 and x60 and not x15 and not x4 and x16 and not x7 and not x12 and x11 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x61 and x60 and not x15 and not x4 and x16 and not x7 and not x12 and not x11 and x8 and x2 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and not x61 and x60 and not x15 and not x4 and x16 and not x7 and not x12 and not x11 and x8 and not x2 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and not x61 and x60 and not x15 and not x4 and x16 and not x7 and not x12 and not x11 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x61 and x60 and not x15 and not x4 and not x16 and x2 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and not x61 and x60 and not x15 and not x4 and not x16 and not x2 and x7 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s318;

      elsif ( x65 and not x61 and x60 and not x15 and not x4 and not x16 and not x2 and not x7 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s191;

      elsif ( x65 and not x61 and not x60 and x62 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and not x61 and not x60 and not x62 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s74;

      elsif ( not x65 and x15 and x66 and x21 and x10 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s330;

      elsif ( not x65 and x15 and x66 and x21 and not x10 and x12 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x65 and x15 and x66 and x21 and not x10 and not x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s48;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and x10 and x23 and x16 and x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s331;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and x10 and x23 and x16 and not x12 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and x10 and x23 and not x16 and x11 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s332;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and x10 and x23 and not x16 and not x11 and x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s48;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and x10 and x23 and not x16 and not x11 and not x12 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and x10 and x23 and not x16 and not x11 and not x12 and not x2 and x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and x10 and x23 and not x16 and not x11 and not x12 and not x2 and not x4 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s333;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and x10 and not x23 and x11 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s334;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and x10 and not x23 and not x11 and x12 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s334;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and x10 and not x23 and not x11 and not x12 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and not x10 and x23 and x11 and x16 and x12 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s330;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and not x10 and x23 and x11 and x16 and not x12 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and not x10 and x23 and x11 and not x16 and x12 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s22;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and not x10 and x23 and x11 and not x16 and not x12 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and not x10 and x23 and not x11 and x16 and x12 and x13 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s335;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and not x10 and x23 and not x11 and x16 and x12 and not x13 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and not x10 and x23 and not x11 and x16 and x12 and not x13 and x17 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and not x10 and x23 and not x11 and x16 and x12 and not x13 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and not x10 and x23 and not x11 and x16 and not x12 and x14 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s335;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and not x10 and x23 and not x11 and x16 and not x12 and not x14 and x17 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and not x10 and x23 and not x11 and x16 and not x12 and not x14 and x17 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and not x10 and x23 and not x11 and x16 and not x12 and not x14 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and not x10 and x23 and not x11 and not x16 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and not x10 and x23 and not x11 and not x16 and not x2 and x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and not x10 and x23 and not x11 and not x16 and not x2 and not x4 and x12 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and not x10 and x23 and not x11 and not x16 and not x2 and not x4 and not x12 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s336;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and not x10 and not x23 and x12 and x11 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and not x10 and not x23 and x12 and not x11 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x65 and x15 and x66 and not x21 and x22 and not x10 and not x23 and not x12 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and x16 and x9 and x7 and x23 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and x16 and x9 and x7 and not x23 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and x16 and x9 and not x7 and x8 and x23 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and x16 and x9 and not x7 and x8 and not x23 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s126;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and x16 and x9 and not x7 and not x8 and x13 and x23 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s337;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and x16 and x9 and not x7 and not x8 and x13 and not x23 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s338;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and x16 and x9 and not x7 and not x8 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and x16 and not x9 and x7 and x23 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and x16 and not x9 and x7 and not x23 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and x16 and not x9 and not x7 and x8 and x23 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s126;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and x16 and not x9 and not x7 and x8 and not x23 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s332;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and x16 and not x9 and not x7 and not x8 and x14 and x23 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s337;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and x16 and not x9 and not x7 and not x8 and x14 and not x23 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s338;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and x16 and not x9 and not x7 and not x8 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and not x16 and x8 and x9 and x7 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and not x16 and x8 and x9 and not x7 and x23 ) = '1' then
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s339;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and not x16 and x8 and x9 and not x7 and not x23 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s331;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and not x16 and x8 and not x9 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and not x16 and not x8 and x7 and x9 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and not x16 and not x8 and x7 and not x9 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and not x16 and not x8 and x7 and not x9 and not x2 and x3 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and not x16 and not x8 and x7 and not x9 and not x2 and not x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s340;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and not x16 and not x8 and not x7 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and not x16 and not x8 and not x7 and not x2 and x3 and x23 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and not x16 and not x8 and not x7 and not x2 and x3 and not x23 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and not x16 and not x8 and not x7 and not x2 and not x3 and x9 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s286;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and not x16 and not x8 and not x7 and not x2 and not x3 and not x9 and x23 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s341;

      elsif ( not x65 and x15 and x66 and not x21 and not x22 and not x16 and not x8 and not x7 and not x2 and not x3 and not x9 and not x23 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x15 and not x66 and x8 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and x15 and not x66 and not x8 and x6 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s207;

      elsif ( not x65 and x15 and not x66 and not x8 and not x6 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and not x15 and x16 and x66 and x21 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s286;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and x10 and x23 and x12 and x8 and x2 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s341;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and x10 and x23 and x12 and x8 and not x2 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and x10 and x23 and x12 and x8 and not x2 and x17 and not x14 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and x10 and x23 and x12 and x8 and not x2 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and x10 and x23 and x12 and x8 and not x2 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and x10 and x23 and x12 and not x8 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and x10 and x23 and x12 and not x8 and not x2 and x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and x10 and x23 and x12 and not x8 and not x2 and not x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and x10 and x23 and not x12 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and x10 and x23 and not x12 and not x2 and x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s342;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and x10 and x23 and not x12 and not x2 and not x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and x10 and not x23 and x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s286;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and x10 and not x23 and not x12 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s341;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and x12 and x7 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and x12 and x7 and not x2 and x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and x12 and x7 and not x2 and not x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and x12 and not x7 and x11 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and x12 and not x7 and x11 and not x2 and x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and x12 and not x7 and x11 and not x2 and not x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and x12 and not x7 and not x11 and x2 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s341;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and x12 and not x7 and not x11 and not x2 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and x12 and not x7 and not x11 and not x2 and x17 and not x14 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and x12 and not x7 and not x11 and not x2 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and x12 and not x7 and not x11 and not x2 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and not x12 and x11 and x9 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and not x12 and x11 and x9 and not x2 and x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and not x12 and x11 and x9 and not x2 and not x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and not x12 and x11 and not x9 and x2 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s341;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and not x12 and x11 and not x9 and not x2 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and not x12 and x11 and not x9 and not x2 and x17 and not x14 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and not x12 and x11 and not x9 and not x2 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and not x12 and x11 and not x9 and not x2 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and not x12 and not x11 and x8 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and not x12 and not x11 and x8 and not x2 and x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and not x12 and not x11 and x8 and not x2 and not x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and not x12 and not x11 and not x8 and x2 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s341;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and not x12 and not x11 and not x8 and not x2 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and not x12 and not x11 and not x8 and not x2 and x17 and not x14 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and not x12 and not x11 and not x8 and not x2 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and x23 and not x12 and not x11 and not x8 and not x2 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and x22 and not x10 and not x23 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s286;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and x9 and x7 and x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and x9 and x7 and not x11 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and x9 and x7 and not x11 and not x2 and x23 and x3 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and x9 and x7 and not x11 and not x2 and x23 and not x3 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s331;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and x9 and x7 and not x11 and not x2 and not x23 and x3 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and x9 and x7 and not x11 and not x2 and not x23 and not x3 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and x9 and not x7 and x10 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and x9 and not x7 and x10 and not x2 and x23 and x3 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and x9 and not x7 and x10 and not x2 and x23 and not x3 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s331;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and x9 and not x7 and x10 and not x2 and not x23 and x3 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and x9 and not x7 and x10 and not x2 and not x23 and not x3 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and x9 and not x7 and not x10 and x8 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and x9 and not x7 and not x10 and x8 and not x2 and x23 and x3 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and x9 and not x7 and not x10 and x8 and not x2 and x23 and not x3 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s331;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and x9 and not x7 and not x10 and x8 and not x2 and not x23 and x3 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and x9 and not x7 and not x10 and x8 and not x2 and not x23 and not x3 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and x9 and not x7 and not x10 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and x7 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and x7 and not x2 and x23 and x3 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s342;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and x7 and not x2 and x23 and not x3 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and x7 and not x2 and not x23 and x3 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s343;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and x7 and not x2 and not x23 and not x3 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and not x7 and x8 and x12 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and not x7 and x8 and x12 and not x2 and x23 and x3 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and not x7 and x8 and x12 and not x2 and x23 and not x3 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s331;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and not x7 and x8 and x12 and not x2 and not x23 and x3 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and not x7 and x8 and x12 and not x2 and not x23 and not x3 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and not x7 and x8 and not x12 and x23 and x19 and x14 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and not x7 and x8 and not x12 and x23 and x19 and not x14 and x13 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and not x7 and x8 and not x12 and x23 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and not x7 and x8 and not x12 and x23 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and not x7 and x8 and not x12 and not x23 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and not x7 and not x8 and x11 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and not x7 and not x8 and x11 and not x2 and x23 and x3 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and not x7 and not x8 and x11 and not x2 and x23 and not x3 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s331;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and not x7 and not x8 and x11 and not x2 and not x23 and x3 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and not x7 and not x8 and x11 and not x2 and not x23 and not x3 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x15 and x16 and x66 and not x21 and not x22 and not x9 and not x7 and not x8 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x15 and x16 and not x66 and x8 and x7 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and not x15 and x16 and not x66 and x8 and not x7 and x9 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and not x15 and x16 and not x66 and x8 and not x7 and not x9 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x15 and x16 and not x66 and x8 and not x7 and not x9 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x15 and x16 and not x66 and x8 and not x7 and not x9 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x15 and x16 and not x66 and x8 and not x7 and not x9 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x15 and x16 and not x66 and not x8 and x7 and x11 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and not x15 and x16 and not x66 and not x8 and x7 and not x11 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x15 and x16 and not x66 and not x8 and x7 and not x11 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x15 and x16 and not x66 and not x8 and x7 and not x11 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x15 and x16 and not x66 and not x8 and x7 and not x11 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x15 and x16 and not x66 and not x8 and not x7 and x10 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and not x15 and x16 and not x66 and not x8 and not x7 and not x10 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x15 and x16 and not x66 and not x8 and not x7 and not x10 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x15 and x16 and not x66 and not x8 and not x7 and not x10 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x15 and x16 and not x66 and not x8 and not x7 and not x10 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x15 and not x16 and x66 and x21 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s340;

      elsif ( not x65 and not x15 and not x16 and x66 and not x21 and x22 and x23 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( not x65 and not x15 and not x16 and x66 and not x21 and x22 and x23 and not x2 and x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( not x65 and not x15 and not x16 and x66 and not x21 and x22 and x23 and not x2 and not x4 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and not x15 and not x16 and x66 and not x21 and x22 and not x23 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s81;

      elsif ( not x65 and not x15 and not x16 and x66 and not x21 and not x22 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( not x65 and not x15 and not x16 and x66 and not x21 and not x22 and not x2 and x23 and x3 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( not x65 and not x15 and not x16 and x66 and not x21 and not x22 and not x2 and x23 and not x3 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s332;

      elsif ( not x65 and not x15 and not x16 and x66 and not x21 and not x22 and not x2 and not x23 and x3 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and not x15 and not x16 and x66 and not x21 and not x22 and not x2 and not x23 and not x3 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s48;

      elsif ( not x65 and not x15 and not x16 and not x66 and x6 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      else
         y8 <= '1' ;
         current_group15m <= s92;

      end if;

   when s77 =>
      if ( x65 and x66 and x67 and x22 and x17 and x18 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and x67 and x22 and x17 and not x18 and x19 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and x67 and x22 and x17 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x67 and x22 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x67 and not x22 and x18 and x13 and x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and x66 and x67 and not x22 and x18 and x13 and not x23 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x66 and x67 and not x22 and x18 and not x13 and x12 and x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and x66 and x67 and not x22 and x18 and not x13 and x12 and not x23 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x66 and x67 and not x22 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x67 and not x22 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x67 and x21 and x20 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and not x67 and x21 and x20 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and not x67 and x21 and x20 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x67 and x21 and x20 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x67 and x21 and not x20 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x66 and not x67 and x21 and not x20 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x66 and not x67 and x21 and not x20 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x67 and x21 and not x20 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x67 and not x21 and x19 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x66 and not x67 and not x21 and x19 and not x14 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x66 and not x67 and not x21 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x67 and not x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x21 and x18 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x65 and not x66 and x21 and not x18 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x21 and not x18 and x19 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x21 and not x18 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x21 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and x23 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( x65 and not x66 and not x21 and x22 and x23 and not x19 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x66 and not x21 and x22 and x23 and not x19 and x17 and not x14 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x66 and not x21 and x22 and x23 and not x19 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and x23 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x23 and x18 and x14 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x21 and x22 and not x23 and x18 and not x14 and x13 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x21 and x22 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x22 and x23 and x20 and x14 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x66 and not x21 and not x22 and x23 and x20 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x66 and not x21 and not x22 and x23 and x20 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x22 and x23 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x22 and not x23 and x15 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( x65 and not x66 and not x21 and not x22 and not x23 and not x15 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s205;

      elsif ( not x65 and x66 and x67 and x68 and x21 and x19 and x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and x66 and x67 and x68 and x21 and x19 and not x15 and x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and x66 and x67 and x68 and x21 and x19 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and x68 and x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and x68 and not x21 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s344;

      elsif ( not x65 and x66 and x67 and not x68 and x62 and x61 and x13 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and x66 and x67 and not x68 and x62 and x61 and not x13 and x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and x66 and x67 and not x68 and x62 and x61 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x68 and x62 and not x61 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and x63 and x17 and x13 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and x63 and x17 and x13 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and x63 and x17 and not x13 and x12 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and x63 and x17 and not x13 and x12 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and x63 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and x63 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and not x63 and x19 and x13 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and not x63 and x19 and x13 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and not x63 and x19 and not x13 and x12 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and not x63 and x19 and not x13 and x12 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and not x63 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x68 and not x62 and not x63 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and x21 and x68 ) = '1' then
         y8 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s82;

      elsif ( not x65 and x66 and not x67 and x21 and not x68 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s143;

      elsif ( not x65 and x66 and not x67 and not x21 and x68 and x22 and x7 and x8 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and x66 and not x67 and not x21 and x68 and x22 and x7 and not x8 and x9 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and x66 and not x67 and not x21 and x68 and x22 and x7 and not x8 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and not x21 and x68 and x22 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and not x21 and x68 and not x22 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x66 and not x67 and not x21 and x68 and not x22 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x66 and not x67 and not x21 and x68 and not x22 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and not x21 and x68 and not x22 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and not x21 and not x68 and x23 and x22 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x65 and x66 and not x67 and not x21 and not x68 and x23 and not x22 and x19 and x14 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x65 and x66 and not x67 and not x21 and not x68 and x23 and not x22 and x19 and not x14 and x13 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x65 and x66 and not x67 and not x21 and not x68 and x23 and not x22 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and not x21 and not x68 and x23 and not x22 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and not x21 and not x68 and not x23 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and not x66 and x68 and x20 and x18 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x66 and x68 and x20 and x18 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x66 and x68 and x20 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x68 and x20 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x68 and not x20 and x21 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x66 and x68 and not x20 and x21 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x66 and x68 and not x20 and x21 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x68 and not x20 and x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x68 and not x20 and not x21 and x17 and x13 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x65 and not x66 and x68 and not x20 and not x21 and x17 and not x13 and x12 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x65 and not x66 and x68 and not x20 and not x21 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x68 and not x20 and not x21 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x68 and x24 and x26 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( not x65 and not x66 and not x68 and x24 and not x26 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and not x66 and not x68 and x24 and not x26 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and not x66 and not x68 and x24 and not x26 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x68 and x24 and not x26 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x68 and not x24 and x25 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and not x68 and not x24 and x25 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and not x68 and not x24 and x25 and x19 and not x14 and not x13 and x26 ) = '1' then
         current_group15m <= s77;

      elsif ( not x65 and not x66 and not x68 and not x24 and x25 and x19 and not x14 and not x13 and not x26 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x68 and not x24 and x25 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x68 and not x24 and not x25 and x26 and x4 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x65 and not x66 and not x68 and not x24 and not x25 and x26 and not x4 and x19 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and not x66 and not x68 and not x24 and not x25 and x26 and not x4 and not x19 and x20 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and not x66 and not x68 and not x24 and not x25 and x26 and not x4 and not x19 and not x20 and x21 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and not x66 and not x68 and not x24 and not x25 and x26 and not x4 and not x19 and not x20 and not x21 and x22 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and not x66 and not x68 and not x24 and not x25 and x26 and not x4 and not x19 and not x20 and not x21 and not x22 and x16 and x11 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x66 and not x68 and not x24 and not x25 and x26 and not x4 and not x19 and not x20 and not x21 and not x22 and x16 and not x11 and x12 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x66 and not x68 and not x24 and not x25 and x26 and not x4 and not x19 and not x20 and not x21 and not x22 and x16 and not x11 and not x12 and x10 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and not x66 and not x68 and not x24 and not x25 and x26 and not x4 and not x19 and not x20 and not x21 and not x22 and x16 and not x11 and not x12 and not x10 ) = '1' then
         y12 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s49;

      elsif ( not x65 and not x66 and not x68 and not x24 and not x25 and x26 and not x4 and not x19 and not x20 and not x21 and not x22 and not x16 and x17 and x10 and x12 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( not x65 and not x66 and not x68 and not x24 and not x25 and x26 and not x4 and not x19 and not x20 and not x21 and not x22 and not x16 and x17 and x10 and not x12 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and not x66 and not x68 and not x24 and not x25 and x26 and not x4 and not x19 and not x20 and not x21 and not x22 and not x16 and x17 and not x10 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( not x65 and not x66 and not x68 and not x24 and not x25 and x26 and not x4 and not x19 and not x20 and not x21 and not x22 and not x16 and not x17 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x66 and not x68 and not x24 and not x25 and not x26 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x65 and not x66 and not x68 and not x24 and not x25 and not x26 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x65 and not x66 and not x68 and not x24 and not x25 and not x26 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s78 =>
      if ( x65 and x66 and x61 and x60 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x66 and x61 and x60 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x66 and x61 and x60 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x66 and x61 and x60 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x66 and x61 and not x60 and x62 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x66 and x61 and not x60 and x62 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x66 and x61 and not x60 and x62 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x61 and not x60 and x62 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x61 and not x60 and not x62 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and x61 and not x60 and not x62 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and x61 and not x60 and not x62 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x66 and x61 and not x60 and not x62 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x66 and not x61 and x60 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and not x61 and x60 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and not x61 and x60 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x66 and not x61 and x60 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x66 and not x61 and not x60 and x62 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and x66 and not x61 and not x60 and not x62 ) = '1' then
         y2 <= '1' ;
         y10 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s263;

      elsif ( x65 and not x66 and x67 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x67 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x67 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and not x68 and x22 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and not x68 and not x22 ) = '1' then
         y28 <= '1' ;
         current_group15m <= s94;

      elsif ( not x65 and x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x7 and x8 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and not x21 and x7 and not x8 and x9 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and not x21 and x7 and not x8 and not x9 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s79 =>
      if ( x21 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( not x21 and x22 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x10 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s226;

      elsif ( not x21 and not x22 and not x10 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x21 and not x22 and not x10 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x21 and not x22 and not x10 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s80 =>
      if ( x22 ) = '1' then
         current_group15m <= s1;

      elsif ( not x22 and x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x22 and not x21 and x23 and x15 and x7 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s81;

      elsif ( not x22 and not x21 and x23 and x15 and not x7 and x9 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x22 and not x21 and x23 and x15 and not x7 and not x9 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x22 and not x21 and x23 and not x15 and x7 and x9 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s330;

      elsif ( not x22 and not x21 and x23 and not x15 and x7 and not x9 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( not x22 and not x21 and x23 and not x15 and not x7 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s330;

      else
         y14 <= '1' ;
         current_group15m <= s285;

      end if;

   when s81 =>
      if ( x21 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s336;

      elsif ( not x21 and x22 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x21 and not x22 and x23 and x19 and x14 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x21 and not x22 and x23 and x19 and not x14 and x13 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x21 and not x22 and x23 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and not x19 ) = '1' then
         current_group15m <= s1;

      else
         y12 <= '1' ;
         current_group15m <= s100;

      end if;

   when s82 =>
      if ( x21 and x66 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( x21 and not x66 and x3 and x4 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( x21 and not x66 and x3 and not x4 and x5 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( x21 and not x66 and x3 and not x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x66 and not x3 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x66 and x22 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s232;

      elsif ( not x21 and x66 and not x22 and x16 and x15 and x10 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s219;

      elsif ( not x21 and x66 and not x22 and x16 and x15 and not x10 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s309;

      elsif ( not x21 and x66 and not x22 and x16 and not x15 and x10 ) = '1' then
         y2 <= '1' ;
         y16 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s124;

      elsif ( not x21 and x66 and not x22 and x16 and not x15 and not x10 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s310;

      elsif ( not x21 and x66 and not x22 and not x16 and x17 and x10 and x15 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s219;

      elsif ( not x21 and x66 and not x22 and not x16 and x17 and x10 and not x15 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s308;

      elsif ( not x21 and x66 and not x22 and not x16 and x17 and not x10 ) = '1' then
         y2 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s79;

      elsif ( not x21 and x66 and not x22 and not x16 and not x17 and x10 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s219;

      elsif ( not x21 and x66 and not x22 and not x16 and not x17 and not x10 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s311;

      elsif ( not x21 and not x66 and x8 and x9 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x21 and not x66 and x8 and not x9 and x10 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x21 and not x66 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s83 =>
      if ( x65 and x66 and x68 and x21 and x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x68 and x21 and not x20 and x18 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s299;

      elsif ( x65 and x66 and x68 and x21 and not x20 and not x18 and x15 and x10 and x11 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s192;

      elsif ( x65 and x66 and x68 and x21 and not x20 and not x18 and x15 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s193;

      elsif ( x65 and x66 and x68 and x21 and not x20 and not x18 and x15 and x10 and not x11 and not x12 ) = '1' then
         y1 <= '1' ;
         y8 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s192;

      elsif ( x65 and x66 and x68 and x21 and not x20 and not x18 and x15 and not x10 and x12 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s300;

      elsif ( x65 and x66 and x68 and x21 and not x20 and not x18 and x15 and not x10 and not x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s192;

      elsif ( x65 and x66 and x68 and x21 and not x20 and not x18 and not x15 and x16 and x10 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x66 and x68 and x21 and not x20 and not x18 and not x15 and x16 and x10 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x66 and x68 and x21 and not x20 and not x18 and not x15 and x16 and x10 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x68 and x21 and not x20 and not x18 and not x15 and x16 and x10 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x68 and x21 and not x20 and not x18 and not x15 and x16 and not x10 and x12 and x11 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s199;

      elsif ( x65 and x66 and x68 and x21 and not x20 and not x18 and not x15 and x16 and not x10 and x12 and not x11 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x66 and x68 and x21 and not x20 and not x18 and not x15 and x16 and not x10 and x12 and not x11 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x66 and x68 and x21 and not x20 and not x18 and not x15 and x16 and not x10 and x12 and not x11 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x68 and x21 and not x20 and not x18 and not x15 and x16 and not x10 and x12 and not x11 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x68 and x21 and not x20 and not x18 and not x15 and x16 and not x10 and not x12 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x66 and x68 and x21 and not x20 and not x18 and not x15 and x16 and not x10 and not x12 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x66 and x68 and x21 and not x20 and not x18 and not x15 and x16 and not x10 and not x12 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x68 and x21 and not x20 and not x18 and not x15 and x16 and not x10 and not x12 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x68 and x21 and not x20 and not x18 and not x15 and not x16 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s201;

      elsif ( x65 and x66 and x68 and not x21 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and x60 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and x16 and x4 and x11 and x12 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s15;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and x16 and x4 and x11 and not x12 and x13 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s345;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and x16 and x4 and x11 and not x12 and not x13 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and x16 and x4 and not x11 and x13 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and x16 and x4 and not x11 and not x13 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and x16 and not x4 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and x13 and x11 and x9 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and x13 and x11 and not x9 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and x13 and x11 and not x9 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and x13 and x11 and not x9 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and x13 and x11 and not x9 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and x13 and not x11 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and x13 and not x11 and not x8 and x12 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and x13 and not x11 and not x8 and not x12 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and x13 and not x11 and not x8 and not x12 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and x13 and not x11 and not x8 and not x12 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and x13 and not x11 and not x8 and not x12 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and not x13 and x11 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and not x13 and not x11 and x12 and x10 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and not x13 and not x11 and x12 and not x10 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and not x13 and not x11 and x12 and not x10 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and not x13 and not x11 and x12 and not x10 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and not x13 and not x11 and x12 and not x10 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and not x13 and not x11 and not x12 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and not x13 and not x11 and not x12 and not x7 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and not x13 and not x11 and not x12 and not x7 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and not x13 and not x11 and not x12 and not x7 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and x17 and not x13 and not x11 and not x12 and not x7 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and not x17 and x45 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x16 and not x17 and not x45 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and x66 and not x68 and not x60 and not x61 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and x21 and x68 and x18 ) = '1' then
         y14 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s116;

      elsif ( x65 and not x66 and x67 and x21 and x68 and not x18 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s117;

      elsif ( x65 and not x66 and x67 and x21 and not x68 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x67 and x21 and not x68 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x67 and x21 and not x68 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and x21 and not x68 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and not x21 and x22 and x68 and x8 and x23 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x66 and x67 and not x21 and x22 and x68 and x8 and x23 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x66 and x67 and not x21 and x22 and x68 and x8 and x23 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and not x21 and x22 and x68 and x8 and not x23 and x9 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x66 and x67 and not x21 and x22 and x68 and x8 and not x23 and not x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x66 and x67 and not x21 and x22 and x68 and x8 and not x23 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and not x21 and x22 and x68 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and not x21 and x22 and not x68 and x19 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x67 and not x21 and x22 and not x68 and x19 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x67 and not x21 and x22 and not x68 and x19 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and not x21 and x22 and not x68 and x19 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and not x21 and x22 and not x68 and not x19 and x18 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x67 and not x21 and x22 and not x68 and not x19 and x18 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x67 and not x21 and x22 and not x68 and not x19 and x18 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and not x21 and x22 and not x68 and not x19 and x18 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and not x21 and x22 and not x68 and not x19 and not x18 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and x67 and not x21 and not x22 and x68 and x23 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x66 and x67 and not x21 and not x22 and x68 and x23 and x9 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x66 and x67 and not x21 and not x22 and x68 and x23 and x9 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and not x21 and not x22 and x68 and x23 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and not x21 and not x22 and x68 and not x23 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x66 and x67 and not x21 and not x22 and x68 and not x23 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x66 and x67 and not x21 and not x22 and x68 and not x23 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and not x21 and not x22 and x68 and not x23 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and not x21 and not x22 and not x68 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x67 and not x21 and not x22 and not x68 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x67 and not x21 and not x22 and not x68 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and not x21 and not x22 and not x68 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and x14 and x17 and x20 and x16 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and x14 and x17 and x20 and not x16 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s346;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and x14 and x17 and not x20 and x16 ) = '1' then
         y13 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s347;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and x14 and x17 and not x20 and not x16 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and x14 and not x17 and x16 and x4 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s348;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and x14 and not x17 and x16 and not x4 ) = '1' then
         y10 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s349;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and x14 and not x17 and not x16 and x20 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and x14 and not x17 and not x16 and x20 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and x14 and not x17 and not x16 and x20 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and x14 and not x17 and not x16 and x20 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and x14 and not x17 and not x16 and not x20 ) = '1' then
         y15 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s350;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and x15 and x17 and x20 and x16 ) = '1' then
         y9 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and x15 and x17 and x20 and not x16 ) = '1' then
         y4 <= '1' ;
         y12 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and x15 and x17 and not x20 and x16 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s346;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and x15 and x17 and not x20 and not x16 ) = '1' then
         y9 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and x15 and not x17 and x16 ) = '1' then
         y15 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s350;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and x15 and not x17 and not x16 and x13 ) = '1' then
         y15 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s350;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and x15 and not x17 and not x16 and not x13 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and x15 and not x17 and not x16 and not x13 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and x15 and not x17 and not x16 and not x13 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and x15 and not x17 and not x16 and not x13 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and not x15 and x17 and x6 and x16 and x7 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and not x15 and x17 and x6 and x16 and not x7 and x5 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and not x15 and x17 and x6 and x16 and not x7 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and not x15 and x17 and x6 and not x16 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and not x15 and x17 and not x6 and x7 and x16 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and not x15 and x17 and not x6 and x7 and not x16 and x5 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and not x15 and x17 and not x6 and x7 and not x16 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and not x15 and x17 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and not x15 and not x17 and x16 and x12 ) = '1' then
         y15 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s350;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and not x15 and not x17 and x16 and not x12 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and not x15 and not x17 and x16 and not x12 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and not x15 and not x17 and x16 and not x12 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and not x15 and not x17 and x16 and not x12 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and not x15 and not x17 and not x16 and x11 ) = '1' then
         y15 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s350;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and not x15 and not x17 and not x16 and not x11 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and not x15 and not x17 and not x16 and not x11 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and not x15 and not x17 and not x16 and not x11 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and x19 and not x14 and not x15 and not x17 and not x16 and not x11 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and x17 and x20 and x14 and x13 ) = '1' then
         y10 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s349;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and x17 and x20 and x14 and not x13 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and x17 and x20 and not x14 and x13 ) = '1' then
         y2 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s349;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and x17 and x20 and not x14 and not x13 and x6 ) = '1' then
         y6 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s102;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and x17 and x20 and not x14 and not x13 and not x6 and x5 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and x17 and x20 and not x14 and not x13 and not x6 and x5 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and x17 and x20 and not x14 and not x13 and not x6 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and x17 and not x20 and x15 and x14 ) = '1' then
         y10 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s349;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and x17 and not x20 and x15 and not x14 ) = '1' then
         y6 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s102;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and x17 and not x20 and not x15 and x14 ) = '1' then
         y15 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s350;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and x17 and not x20 and not x15 and not x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and x20 and x13 and x12 and x14 ) = '1' then
         y15 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s350;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and x20 and x13 and x12 and not x14 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and x20 and x13 and x12 and not x14 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and x20 and x13 and x12 and not x14 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and x20 and x13 and x12 and not x14 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and x20 and x13 and not x12 ) = '1' then
         y15 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s350;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and x20 and not x13 and x11 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and x20 and not x13 and x11 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and x20 and not x13 and x11 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and x20 and not x13 and x11 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and x20 and not x13 and not x11 ) = '1' then
         y15 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s350;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and not x20 and x14 and x13 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s348;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and not x20 and x14 and not x13 and x15 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s348;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and not x20 and x14 and not x13 and not x15 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and not x20 and x14 and not x13 and not x15 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and not x20 and x14 and not x13 and not x15 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and not x20 and x14 and not x13 and not x15 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and not x20 and not x14 and x15 and x12 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s348;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and not x20 and not x14 and x15 and not x12 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and not x20 and not x14 and x15 and not x12 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and not x20 and not x14 and x15 and not x12 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and not x20 and not x14 and x15 and not x12 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and not x20 and not x14 and not x15 and x11 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s348;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and not x20 and not x14 and not x15 and not x11 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and not x20 and not x14 and not x15 and not x11 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and not x20 and not x14 and not x15 and not x11 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and x18 and not x19 and not x17 and not x20 and not x14 and not x15 and not x11 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and x20 and x19 and x14 and x15 ) = '1' then
         y29 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and x20 and x19 and x14 and not x15 and x16 ) = '1' then
         y29 <= '1' ;
         y31 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and x20 and x19 and x14 and not x15 and not x16 and x4 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s348;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and x20 and x19 and x14 and not x15 and not x16 and not x4 ) = '1' then
         y4 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and x20 and x19 and not x14 and x16 and x15 and x13 ) = '1' then
         y29 <= '1' ;
         y31 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and x20 and x19 and not x14 and x16 and x15 and not x13 ) = '1' then
         y29 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and x20 and x19 and not x14 and x16 and not x15 and x4 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s348;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and x20 and x19 and not x14 and x16 and not x15 and not x4 ) = '1' then
         y4 <= '1' ;
         y17 <= '1' ;
         y29 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and x20 and x19 and not x14 and not x16 and x15 ) = '1' then
         y4 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and x20 and x19 and not x14 and not x16 and not x15 and x4 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and x20 and x19 and not x14 and not x16 and not x15 and not x4 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and x20 and not x19 and x16 and x14 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and x20 and not x19 and x16 and not x14 and x4 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and x20 and not x19 and x16 and not x14 and not x4 ) = '1' then
         y16 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s352;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and x20 and not x19 and not x16 and x13 and x14 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and x20 and not x19 and not x16 and x13 and x14 and not x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and x20 and not x19 and not x16 and x13 and not x14 and x4 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and x20 and not x19 and not x16 and x13 and not x14 and not x4 ) = '1' then
         y4 <= '1' ;
         y12 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and x20 and not x19 and not x16 and not x13 and x4 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and x20 and not x19 and not x16 and not x13 and not x4 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s346;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and not x20 and x14 and x19 and x15 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and not x20 and x14 and x19 and not x15 and x16 ) = '1' then
         y29 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and not x20 and x14 and x19 and not x15 and not x16 and x4 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s348;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and not x20 and x14 and x19 and not x15 and not x16 and not x4 ) = '1' then
         y4 <= '1' ;
         y29 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and not x20 and x14 and not x19 and x16 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s346;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and not x20 and x14 and not x19 and not x16 and x15 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and not x20 and x14 and not x19 and not x16 and x15 and not x13 ) = '1' then
         y4 <= '1' ;
         y12 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and not x20 and x14 and not x19 and not x16 and not x15 ) = '1' then
         y9 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and not x20 and not x14 and x15 and x16 and x19 and x13 ) = '1' then
         y29 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and not x20 and not x14 and x15 and x16 and x19 and not x13 ) = '1' then
         y4 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and not x20 and not x14 and x15 and x16 and not x19 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and not x20 and not x14 and x15 and not x16 and x4 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s348;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and not x20 and not x14 and x15 and not x16 and not x4 and x19 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and not x20 and not x14 and x15 and not x16 and not x4 and not x19 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and not x20 and not x14 and not x15 and x4 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s348;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and not x20 and not x14 and not x15 and not x4 and x19 and x16 ) = '1' then
         y29 <= '1' ;
         y31 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and not x20 and not x14 and not x15 and not x4 and x19 and not x16 ) = '1' then
         y4 <= '1' ;
         y12 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and not x20 and not x14 and not x15 and not x4 and not x19 and x16 ) = '1' then
         y16 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s352;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and x17 and not x20 and not x14 and not x15 and not x4 and not x19 and not x16 ) = '1' then
         y13 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s347;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and not x17 and x4 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s348;

      elsif ( x65 and not x66 and not x67 and x68 and not x3 and not x18 and not x17 and not x4 ) = '1' then
         y4 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s353;

      elsif ( x65 and not x66 and not x67 and not x68 and x21 and x18 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x65 and not x66 and not x67 and not x68 and x21 and not x18 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x67 and not x68 and x21 and not x18 and x19 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x67 and not x68 and x21 and not x18 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and not x68 and x21 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and not x68 and not x21 and x23 and x22 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( x65 and not x66 and not x67 and not x68 and not x21 and x23 and x22 and not x19 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x66 and not x67 and not x68 and not x21 and x23 and x22 and not x19 and x17 and not x14 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x66 and not x67 and not x68 and not x21 and x23 and x22 and not x19 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and not x68 and not x21 and x23 and x22 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and not x68 and not x21 and x23 and not x22 and x20 and x14 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x66 and not x67 and not x68 and not x21 and x23 and not x22 and x20 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x66 and not x67 and not x68 and not x21 and x23 and not x22 and x20 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and not x68 and not x21 and x23 and not x22 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and not x68 and not x21 and not x23 and x18 and x14 and x22 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x67 and not x68 and not x21 and not x23 and x18 and x14 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x66 and not x67 and not x68 and not x21 and not x23 and x18 and not x14 and x13 and x22 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x67 and not x68 and not x21 and not x23 and x18 and not x14 and x13 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x66 and not x67 and not x68 and not x21 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and not x68 and not x21 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x62 and x61 and x13 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and x67 and x62 and x61 and not x13 and x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and x67 and x62 and x61 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x62 and not x61 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and not x62 and x63 and x17 and x13 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and x67 and not x62 and x63 and x17 and x13 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and x67 and not x62 and x63 and x17 and not x13 and x12 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and x67 and not x62 and x63 and x17 and not x13 and x12 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and x67 and not x62 and x63 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and not x62 and x63 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and not x62 and not x63 and x19 and x13 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x67 and not x62 and not x63 and x19 and x13 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x67 and not x62 and not x63 and x19 and not x13 and x12 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x67 and not x62 and not x63 and x19 and not x13 and x12 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x67 and not x62 and not x63 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and not x62 and not x63 and not x19 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s84 =>
      if ( x21 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x21 and x23 and x22 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s354;

      elsif ( not x21 and x23 and not x22 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s80;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s80;

      end if;

   when s85 =>
      if ( x65 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x65 and x22 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s340;

      else
         y3 <= '1' ;
         y4 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s337;

      end if;

   when s86 =>
      if ( x65 and x66 and x67 and x23 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x67 and not x23 and x6 and x15 and x8 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x66 and x67 and not x23 and x6 and x15 and not x8 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x65 and x66 and x67 and not x23 and x6 and not x15 and x16 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x66 and x67 and not x23 and x6 and not x15 and not x16 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s122;

      elsif ( x65 and x66 and x67 and not x23 and not x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x66 and not x67 and x60 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      elsif ( x65 and x66 and not x67 and not x60 and x61 and x62 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and x66 and not x67 and not x60 and x61 and not x62 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and x15 and x16 and x12 and x7 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s254;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and x15 and x16 and x12 and not x7 and x14 and x11 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and x15 and x16 and x12 and not x7 and x14 and not x11 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s355;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and x15 and x16 and x12 and not x7 and not x14 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and x15 and x16 and not x12 and x7 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and x15 and x16 and not x12 and not x7 and x13 and x11 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and x15 and x16 and not x12 and not x7 and x13 and not x11 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s355;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and x15 and x16 and not x12 and not x7 and not x13 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and x15 and not x16 and x11 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s291;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and x15 and not x16 and x11 and not x7 and x12 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s231;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and x15 and not x16 and x11 and not x7 and not x12 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s210;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and x15 and not x16 and not x11 and x6 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s74;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and x15 and not x16 and not x11 and not x6 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and x15 and not x16 and not x11 and not x6 and not x2 and x12 and x7 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s356;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and x15 and not x16 and not x11 and not x6 and not x2 and x12 and not x7 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s357;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and x15 and not x16 and not x11 and not x6 and not x2 and not x12 and x7 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and x15 and not x16 and not x11 and not x6 and not x2 and not x12 and not x7 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and not x15 and x6 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s74;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and not x15 and not x6 and x16 and x7 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and not x15 and not x6 and x16 and x7 and not x2 and x12 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s357;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and not x15 and not x6 and x16 and x7 and not x2 and not x12 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and not x15 and not x6 and x16 and not x7 and x12 and x11 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and not x15 and not x6 and x16 and not x7 and x12 and x11 and not x2 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s260;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and not x15 and not x6 and x16 and not x7 and x12 and not x11 and x9 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and not x15 and not x6 and x16 and not x7 and x12 and not x11 and x9 and not x2 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s260;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and not x15 and not x6 and x16 and not x7 and x12 and not x11 and not x9 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and not x15 and not x6 and x16 and not x7 and not x12 and x11 and x10 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and not x15 and not x6 and x16 and not x7 and not x12 and x11 and x10 and not x2 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s260;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and not x15 and not x6 and x16 and not x7 and not x12 and x11 and not x10 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and not x15 and not x6 and x16 and not x7 and not x12 and not x11 and x8 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and not x15 and not x6 and x16 and not x7 and not x12 and not x11 and x8 and not x2 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s260;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and not x15 and not x6 and x16 and not x7 and not x12 and not x11 and not x8 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and not x15 and not x6 and not x16 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and not x15 and not x6 and not x16 and not x2 and x7 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and x62 and not x15 and not x6 and not x16 and not x2 and not x7 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s68;

      elsif ( x65 and x66 and not x67 and not x60 and not x61 and not x62 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s65;

      elsif ( x65 and not x66 and x21 and x17 and x16 and x13 and x18 and x15 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and x21 and x17 and x16 and x13 and x18 and not x15 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x65 and not x66 and x21 and x17 and x16 and x13 and not x18 and x14 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x65 and not x66 and x21 and x17 and x16 and x13 and not x18 and not x14 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x65 and not x66 and x21 and x17 and x16 and not x13 and x14 and x18 and x15 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x65 and not x66 and x21 and x17 and x16 and not x13 and x14 and x18 and not x15 ) = '1' then
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s288;

      elsif ( x65 and not x66 and x21 and x17 and x16 and not x13 and x14 and not x18 ) = '1' then
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s288;

      elsif ( x65 and not x66 and x21 and x17 and x16 and not x13 and not x14 and x18 and x15 and x6 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and x21 and x17 and x16 and not x13 and not x14 and x18 and x15 and not x6 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x21 and x17 and x16 and not x13 and not x14 and x18 and x15 and not x6 and x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x21 and x17 and x16 and not x13 and not x14 and x18 and x15 and not x6 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x21 and x17 and x16 and not x13 and not x14 and x18 and not x15 and x5 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and x21 and x17 and x16 and not x13 and not x14 and x18 and not x15 and not x5 and x4 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x21 and x17 and x16 and not x13 and not x14 and x18 and not x15 and not x5 and x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x21 and x17 and x16 and not x13 and not x14 and x18 and not x15 and not x5 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x21 and x17 and x16 and not x13 and not x14 and not x18 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and x13 and x18 and x15 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and x13 and x18 and not x15 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and x13 and x18 and not x15 and not x2 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and x13 and not x18 and x14 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and x13 and not x18 and x14 and not x2 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and x13 and not x18 and x14 and not x2 and not x3 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and x13 and not x18 and not x14 and x12 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and x13 and not x18 and not x14 and x12 and not x2 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and x13 and not x18 and not x14 and x12 and not x2 and not x3 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and x13 and not x18 and not x14 and not x12 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and x13 and not x18 and not x14 and not x12 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and x13 and not x18 and not x14 and not x12 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and x13 and not x18 and not x14 and not x12 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and x14 and x18 and x15 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and x14 and x18 and x15 and not x2 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and x14 and x18 and not x15 and x12 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and x14 and x18 and not x15 and x12 and not x2 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and x14 and x18 and not x15 and not x12 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and x14 and x18 and not x15 and not x12 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and x14 and x18 and not x15 and not x12 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and x14 and x18 and not x15 and not x12 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and x14 and not x18 and x11 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and x14 and not x18 and x11 and not x2 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and x14 and not x18 and x11 and not x2 and not x3 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and x14 and not x18 and not x11 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and x14 and not x18 and not x11 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and x14 and not x18 and not x11 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and x14 and not x18 and not x11 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and not x14 and x18 and x15 and x11 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and not x14 and x18 and x15 and x11 and not x2 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and not x14 and x18 and x15 and not x11 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and not x14 and x18 and x15 and not x11 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and not x14 and x18 and x15 and not x11 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and not x14 and x18 and x15 and not x11 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and not x14 and x18 and not x15 and x10 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and not x14 and x18 and not x15 and x10 and not x2 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and not x14 and x18 and not x15 and not x10 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and not x14 and x18 and not x15 and not x10 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and not x14 and x18 and not x15 and not x10 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and not x14 and x18 and not x15 and not x10 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and not x14 and not x18 and x10 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and not x14 and not x18 and x10 and not x2 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and not x14 and not x18 and x10 and not x2 and not x3 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and not x14 and not x18 and not x10 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and not x14 and not x18 and not x10 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and not x14 and not x18 and not x10 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x21 and x17 and not x16 and not x13 and not x14 and not x18 and not x10 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x21 and not x17 and x16 and x14 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x66 and x21 and not x17 and x16 and x14 and not x13 and x15 and x18 and x12 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( x65 and not x66 and x21 and not x17 and x16 and x14 and not x13 and x15 and x18 and not x12 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s169;

      elsif ( x65 and not x66 and x21 and not x17 and x16 and x14 and not x13 and x15 and not x18 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( x65 and not x66 and x21 and not x17 and x16 and x14 and not x13 and not x15 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s174;

      elsif ( x65 and not x66 and x21 and not x17 and x16 and not x14 and x15 and x18 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( x65 and not x66 and x21 and not x17 and x16 and not x14 and x15 and x18 and not x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s346;

      elsif ( x65 and not x66 and x21 and not x17 and x16 and not x14 and x15 and not x18 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s346;

      elsif ( x65 and not x66 and x21 and not x17 and x16 and not x14 and x15 and not x18 and not x13 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s169;

      elsif ( x65 and not x66 and x21 and not x17 and x16 and not x14 and not x15 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and x21 and not x17 and x16 and not x14 and not x15 and not x2 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and x21 and not x17 and x16 and not x14 and not x15 and not x2 and not x3 and x13 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and x21 and not x17 and x16 and not x14 and not x15 and not x2 and not x3 and not x13 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s300;

      elsif ( x65 and not x66 and x21 and not x17 and not x16 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and x21 and not x17 and not x16 and not x2 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and x21 and not x17 and not x16 and not x2 and not x3 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s51;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and x19 and x10 and x15 ) = '1' then
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s288;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and x19 and x10 and not x15 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s300;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and x19 and not x10 and x15 and x6 and x14 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s360;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and x19 and not x10 and x15 and x6 and not x14 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and x19 and not x10 and x15 and not x6 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and x19 and not x10 and x15 and not x6 and x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and x19 and not x10 and x15 and not x6 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and x19 and not x10 and not x15 and x5 and x14 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and x19 and not x10 and not x15 and x5 and not x14 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and x19 and not x10 and not x15 and not x5 and x4 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and x19 and not x10 and not x15 and not x5 and x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and x19 and not x10 and not x15 and not x5 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and not x19 and x13 and x15 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s300;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and not x19 and x13 and not x15 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s360;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and not x19 and not x13 and x15 and x6 and x14 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and not x19 and not x13 and x15 and x6 and not x14 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and not x19 and not x13 and x15 and not x6 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and not x19 and not x13 and x15 and not x6 and x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and not x19 and not x13 and x15 and not x6 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and not x19 and not x13 and not x15 and x5 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and not x19 and not x13 and not x15 and x5 and not x14 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and not x19 and not x13 and not x15 and not x5 and x4 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and not x19 and not x13 and not x15 and not x5 and x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and x18 and not x19 and not x13 and not x15 and not x5 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and not x18 and x13 and x15 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and not x18 and x13 and not x15 ) = '1' then
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s288;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and not x18 and not x13 and x14 and x19 and x15 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s300;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and not x18 and not x13 and x14 and x19 and not x15 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s360;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and not x18 and not x13 and x14 and not x19 and x15 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s360;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and not x18 and not x13 and x14 and not x19 and not x15 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and not x18 and not x13 and not x14 and x15 and x6 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and not x18 and not x13 and not x14 and x15 and not x6 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and not x18 and not x13 and not x14 and x15 and not x6 and x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and not x18 and not x13 and not x14 and x15 and not x6 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and not x18 and not x13 and not x14 and not x15 and x5 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and not x18 and not x13 and not x14 and not x15 and not x5 and x4 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and not x18 and not x13 and not x14 and not x15 and not x5 and x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and x16 and not x18 and not x13 and not x14 and not x15 and not x5 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and x15 and x19 and x10 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and x15 and x19 and not x10 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and x15 and x19 and not x10 and not x2 and x14 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and x15 and x19 and not x10 and not x2 and x14 and not x3 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and x15 and x19 and not x10 and not x2 and not x14 and x12 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and x15 and x19 and not x10 and not x2 and not x14 and x12 and not x3 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and x15 and x19 and not x10 and not x2 and not x14 and not x12 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and x15 and x19 and not x10 and not x2 and not x14 and not x12 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and x15 and x19 and not x10 and not x2 and not x14 and not x12 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and x15 and x19 and not x10 and not x2 and not x14 and not x12 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and x15 and not x19 and x13 ) = '1' then
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s288;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and x15 and not x19 and not x13 and x14 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and x15 and not x19 and not x13 and x14 and not x2 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and x15 and not x19 and not x13 and x14 and not x2 and not x3 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and x15 and not x19 and not x13 and not x14 and x11 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and x15 and not x19 and not x13 and not x14 and not x11 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and x15 and not x19 and not x13 and not x14 and not x11 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and x15 and not x19 and not x13 and not x14 and not x11 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and x15 and not x19 and not x13 and not x14 and not x11 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and x19 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and x19 and not x2 and x10 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and x19 and not x2 and not x10 and x14 and x13 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and x19 and not x2 and not x10 and x14 and x13 and not x3 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and x19 and not x2 and not x10 and x14 and not x13 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and x19 and not x2 and not x10 and x14 and not x13 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and x19 and not x2 and not x10 and x14 and not x13 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and x19 and not x2 and not x10 and x14 and not x13 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and x19 and not x2 and not x10 and not x14 and x11 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and x19 and not x2 and not x10 and not x14 and x11 and not x3 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and x19 and not x2 and not x10 and not x14 and not x11 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and x19 and not x2 and not x10 and not x14 and not x11 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and x19 and not x2 and not x10 and not x14 and not x11 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and x19 and not x2 and not x10 and not x14 and not x11 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and not x19 and x13 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and not x19 and x13 and not x2 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and not x19 and not x13 and x14 and x12 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and not x19 and not x13 and x14 and not x12 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and not x19 and not x13 and x14 and not x12 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and not x19 and not x13 and x14 and not x12 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and not x19 and not x13 and x14 and not x12 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and not x19 and not x13 and not x14 and x10 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and not x19 and not x13 and not x14 and not x10 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and not x19 and not x13 and not x14 and not x10 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and not x19 and not x13 and not x14 and not x10 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and x18 and not x15 and not x19 and not x13 and not x14 and not x10 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and x13 and x15 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and x13 and not x15 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and x13 and not x15 and not x2 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and x14 and x15 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and x14 and x15 and not x3 and x19 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and x14 and x15 and not x3 and not x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and x14 and not x15 and x12 and x19 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and x14 and not x15 and x12 and x19 and not x3 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and x14 and not x15 and x12 and not x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and x14 and not x15 and not x12 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and x14 and not x15 and not x12 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and x14 and not x15 and not x12 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and x14 and not x15 and not x12 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and not x14 and x15 and x11 and x19 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and not x14 and x15 and x11 and x19 and not x3 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and not x14 and x15 and x11 and not x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and not x14 and x15 and not x11 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and not x14 and x15 and not x11 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and not x14 and x15 and not x11 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and not x14 and x15 and not x11 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and not x14 and not x15 and x10 and x19 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and not x14 and not x15 and x10 and x19 and not x3 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and not x14 and not x15 and x10 and not x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and not x14 and not x15 and not x10 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and not x14 and not x15 and not x10 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and not x14 and not x15 and not x10 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and x22 and not x16 and not x18 and not x13 and not x2 and not x14 and not x15 and not x10 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and x18 and x13 and x15 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and x18 and x13 and not x15 ) = '1' then
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s288;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and x18 and not x13 and x15 and x6 and x14 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s300;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and x18 and not x13 and x15 and x6 and not x14 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and x18 and not x13 and x15 and not x6 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and x18 and not x13 and x15 and not x6 and x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and x18 and not x13 and x15 and not x6 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and x18 and not x13 and not x15 and x5 and x14 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s360;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and x18 and not x13 and not x15 and x5 and not x14 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and x18 and not x13 and not x15 and not x5 and x4 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and x18 and not x13 and not x15 and not x5 and x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and x18 and not x13 and not x15 and not x5 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and not x18 and x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and not x18 and x14 and not x13 and x15 and x16 ) = '1' then
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and not x18 and x14 and not x13 and x15 and not x16 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and not x18 and x14 and not x13 and not x15 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and not x18 and not x14 and x15 and x13 ) = '1' then
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and not x18 and not x14 and x15 and not x13 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and not x18 and not x14 and not x15 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and not x18 and not x14 and not x15 and not x2 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and not x18 and not x14 and not x15 and not x2 and not x3 and x13 ) = '1' then
         y5 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s361;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and x19 and not x18 and not x14 and not x15 and not x2 and not x3 and not x13 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and x16 and x13 and x20 and x14 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and x16 and x13 and x20 and not x14 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and x16 and x13 and not x20 and x15 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and x16 and x13 and not x20 and not x15 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and x16 and not x13 and x14 and x20 ) = '1' then
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s288;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and x16 and not x13 and x14 and not x20 and x15 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and x16 and not x13 and x14 and not x20 and not x15 ) = '1' then
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s288;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and x16 and not x13 and not x14 and x20 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and x16 and not x13 and not x14 and not x20 and x15 and x6 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and x16 and not x13 and not x14 and not x20 and x15 and not x6 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and x16 and not x13 and not x14 and not x20 and x15 and not x6 and x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and x16 and not x13 and not x14 and not x20 and x15 and not x6 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and x16 and not x13 and not x14 and not x20 and not x15 and x5 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and x16 and not x13 and not x14 and not x20 and not x15 and not x5 and x4 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and x16 and not x13 and not x14 and not x20 and not x15 and not x5 and x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and x16 and not x13 and not x14 and not x20 and not x15 and not x5 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and x13 and x20 and x14 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and x13 and x20 and x14 and not x2 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and x13 and x20 and x14 and not x2 and not x3 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and x13 and x20 and not x14 and x12 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and x13 and x20 and not x14 and x12 and not x2 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and x13 and x20 and not x14 and x12 and not x2 and not x3 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and x13 and x20 and not x14 and not x12 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and x13 and x20 and not x14 and not x12 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and x13 and x20 and not x14 and not x12 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and x13 and x20 and not x14 and not x12 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and x13 and not x20 and x15 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and x13 and not x20 and not x15 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and x13 and not x20 and not x15 and not x2 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and x14 and x20 and x11 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and x14 and x20 and x11 and not x2 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and x14 and x20 and x11 and not x2 and not x3 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and x14 and x20 and not x11 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and x14 and x20 and not x11 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and x14 and x20 and not x11 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and x14 and x20 and not x11 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and x14 and not x20 and x15 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and x14 and not x20 and x15 and not x2 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and x14 and not x20 and not x15 and x12 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and x14 and not x20 and not x15 and x12 and not x2 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and x14 and not x20 and not x15 and not x12 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and x14 and not x20 and not x15 and not x12 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and x14 and not x20 and not x15 and not x12 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and x14 and not x20 and not x15 and not x12 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and not x14 and x20 and x10 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and not x14 and x20 and x10 and not x2 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and not x14 and x20 and x10 and not x2 and not x3 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and not x14 and x20 and not x10 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and not x14 and x20 and not x10 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and not x14 and x20 and not x10 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and not x14 and x20 and not x10 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and not x14 and not x20 and x15 and x11 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and not x14 and not x20 and x15 and x11 and not x2 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and not x14 and not x20 and x15 and not x11 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and not x14 and not x20 and x15 and not x11 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and not x14 and not x20 and x15 and not x11 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and not x14 and not x20 and x15 and not x11 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and not x14 and not x20 and not x15 and x10 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and not x14 and not x20 and not x15 and x10 and not x2 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and not x14 and not x20 and not x15 and not x10 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and not x14 and not x20 and not x15 and not x10 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and not x14 and not x20 and not x15 and not x10 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x17 and not x22 and not x19 and not x16 and not x13 and not x14 and not x20 and not x15 and not x10 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and x14 and x18 and x19 and x10 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and x14 and x18 and x19 and not x10 and x15 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and x14 and x18 and x19 and not x10 and not x15 ) = '1' then
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and x14 and x18 and not x19 and x13 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and x14 and x18 and not x19 and not x13 and x15 ) = '1' then
         y5 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s361;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and x14 and x18 and not x19 and not x13 and not x15 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and x14 and not x18 and x19 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and x14 and not x18 and x19 and not x13 and x15 ) = '1' then
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and x14 and not x18 and x19 and not x13 and not x15 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and x14 and not x18 and not x19 and x13 ) = '1' then
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and x14 and not x18 and not x19 and not x13 and x15 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and x14 and not x18 and not x19 and not x13 and not x15 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and x15 and x19 and x18 and x10 ) = '1' then
         y5 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s361;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and x15 and x19 and x18 and not x10 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and x15 and x19 and not x18 and x13 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and x15 and x19 and not x18 and not x13 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and x15 and not x19 and x13 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and x15 and not x19 and not x13 and x18 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and x15 and not x19 and not x13 and x18 and not x3 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and x15 and not x19 and not x13 and not x18 and x3 ) = '1' then
         y5 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s361;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and x15 and not x19 and not x13 and not x18 and not x3 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and not x15 and x2 and x18 and x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and not x15 and x2 and x18 and not x19 and x13 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and not x15 and x2 and x18 and not x19 and not x13 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s362;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and not x15 and x2 and not x18 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and not x15 and not x2 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and not x15 and not x2 and not x3 and x19 and x18 and x10 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and not x15 and not x2 and not x3 and x19 and x18 and not x10 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and not x15 and not x2 and not x3 and x19 and not x18 and x13 ) = '1' then
         y5 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s361;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and not x15 and not x2 and not x3 and x19 and not x18 and not x13 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and not x15 and not x2 and not x3 and not x19 and x13 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s363;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and not x15 and not x2 and not x3 and not x19 and not x13 and x18 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and x16 and not x14 and not x15 and not x2 and not x3 and not x19 and not x13 and not x18 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s362;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and not x16 and x18 and x19 and x10 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and not x16 and x18 and x19 and not x10 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and not x16 and x18 and x19 and not x10 and not x2 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and not x16 and x18 and x19 and not x10 and not x2 and not x3 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s51;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and not x16 and x18 and not x19 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and not x16 and x18 and not x19 and not x2 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and not x16 and x18 and not x19 and not x2 and not x3 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s51;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and not x16 and not x18 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and not x16 and not x18 and not x2 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and not x17 and x22 and not x16 and not x18 and not x2 and not x3 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s51;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and x15 and x13 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and x15 and not x13 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and x15 and not x13 and not x2 and x14 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and x15 and not x13 and not x2 and x14 and not x3 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and x15 and not x13 and not x2 and not x14 and x11 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and x15 and not x13 and not x2 and not x14 and x11 and not x3 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and x15 and not x13 and not x2 and not x14 and not x11 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and x15 and not x13 and not x2 and not x14 and not x11 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and x15 and not x13 and not x2 and not x14 and not x11 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and x15 and not x13 and not x2 and not x14 and not x11 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and not x15 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and not x15 and not x2 and x13 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and not x15 and not x2 and not x13 and x14 and x12 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and not x15 and not x2 and not x13 and x14 and x12 and not x3 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and not x15 and not x2 and not x13 and x14 and not x12 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and not x15 and not x2 and not x13 and x14 and not x12 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and not x15 and not x2 and not x13 and x14 and not x12 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and not x15 and not x2 and not x13 and x14 and not x12 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and not x15 and not x2 and not x13 and not x14 and x10 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and not x15 and not x2 and not x13 and not x14 and x10 and not x3 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and not x15 and not x2 and not x13 and not x14 and not x10 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and not x15 and not x2 and not x13 and not x14 and not x10 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and not x15 and not x2 and not x13 and not x14 and not x10 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and x18 and not x15 and not x2 and not x13 and not x14 and not x10 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and not x18 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and not x18 and not x2 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and x19 and not x18 and not x2 and not x3 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s51;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and not x19 and x16 and x14 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and not x19 and x16 and x14 and not x13 and x15 and x20 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and not x19 and x16 and x14 and not x13 and x15 and not x20 and x12 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and not x19 and x16 and x14 and not x13 and x15 and not x20 and not x12 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and not x19 and x16 and x14 and not x13 and not x15 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s362;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and not x19 and x16 and not x14 and x15 and x20 and x13 ) = '1' then
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and not x19 and x16 and not x14 and x15 and x20 and not x13 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and not x19 and x16 and not x14 and x15 and not x20 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and not x19 and x16 and not x14 and x15 and not x20 and not x13 ) = '1' then
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and not x19 and x16 and not x14 and not x15 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and not x19 and x16 and not x14 and not x15 and not x2 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and not x19 and x16 and not x14 and not x15 and not x2 and not x3 and x13 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and not x19 and x16 and not x14 and not x15 and not x2 and not x3 and not x13 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s300;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and not x19 and not x16 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and not x19 and not x16 and not x2 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s359;

      elsif ( x65 and not x66 and not x21 and not x17 and not x22 and not x19 and not x16 and not x2 and not x3 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s51;

      elsif ( not x65 and x21 and x68 and x16 and x17 and x10 and x15 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and x21 and x68 and x16 and x17 and x10 and not x15 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x65 and x21 and x68 and x16 and x17 and not x10 and x15 and x7 and x14 ) = '1' then
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s288;

      elsif ( not x65 and x21 and x68 and x16 and x17 and not x10 and x15 and x7 and not x14 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( not x65 and x21 and x68 and x16 and x17 and not x10 and x15 and not x7 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x21 and x68 and x16 and x17 and not x10 and x15 and not x7 and x9 and not x8 and x14 ) = '1' then
         current_group15m <= s86;

      elsif ( not x65 and x21 and x68 and x16 and x17 and not x10 and x15 and not x7 and x9 and not x8 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and x68 and x16 and x17 and not x10 and x15 and not x7 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and x68 and x16 and x17 and not x10 and not x15 and x8 and x14 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s310;

      elsif ( not x65 and x21 and x68 and x16 and x17 and not x10 and not x15 and x8 and not x14 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s305;

      elsif ( not x65 and x21 and x68 and x16 and x17 and not x10 and not x15 and not x8 and x9 and x14 ) = '1' then
         current_group15m <= s86;

      elsif ( not x65 and x21 and x68 and x16 and x17 and not x10 and not x15 and not x8 and x9 and not x14 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x21 and x68 and x16 and x17 and not x10 and not x15 and not x8 and x9 and not x14 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and x68 and x16 and x17 and not x10 and not x15 and not x8 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and x68 and x16 and not x17 and x14 and x10 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x21 and x68 and x16 and not x17 and x14 and not x10 and x15 and x13 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s8;

      elsif ( not x65 and x21 and x68 and x16 and not x17 and x14 and not x10 and x15 and not x13 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s122;

      elsif ( not x65 and x21 and x68 and x16 and not x17 and x14 and not x10 and not x15 ) = '1' then
         y2 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s221;

      elsif ( not x65 and x21 and x68 and x16 and not x17 and not x14 and x2 ) = '1' then
         y2 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s322;

      elsif ( not x65 and x21 and x68 and x16 and not x17 and not x14 and not x2 and x4 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x21 and x68 and x16 and not x17 and not x14 and not x2 and not x4 and x15 and x10 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s357;

      elsif ( not x65 and x21 and x68 and x16 and not x17 and not x14 and not x2 and not x4 and x15 and not x10 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s357;

      elsif ( not x65 and x21 and x68 and x16 and not x17 and not x14 and not x2 and not x4 and not x15 and x10 ) = '1' then
         y2 <= '1' ;
         y16 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s124;

      elsif ( not x65 and x21 and x68 and x16 and not x17 and not x14 and not x2 and not x4 and not x15 and not x10 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x65 and x21 and x68 and not x16 and x2 ) = '1' then
         y2 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s322;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and x10 and x4 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and x10 and not x4 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s297;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and not x10 and x14 and x15 and x4 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and not x10 and x14 and x15 and not x4 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and not x10 and x14 and not x15 and x13 and x4 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and not x10 and x14 and not x15 and x13 and not x4 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and not x10 and x14 and not x15 and not x13 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and not x10 and x14 and not x15 and not x13 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and not x10 and x14 and not x15 and not x13 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and not x10 and x14 and not x15 and not x13 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and x15 and x12 and x4 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and x15 and x12 and not x4 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and x15 and not x12 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and x15 and not x12 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and x15 and not x12 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and x15 and not x12 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and not x15 and x11 and x4 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and not x15 and x11 and not x4 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and not x15 and not x11 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and not x15 and not x11 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and not x15 and not x11 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and x17 and not x10 and not x14 and not x15 and not x11 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and not x17 and x4 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and not x17 and not x4 and x10 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s296;

      elsif ( not x65 and x21 and x68 and not x16 and not x2 and not x17 and not x4 and not x10 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s356;

      elsif ( not x65 and x21 and not x68 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s143;

      elsif ( not x65 and not x21 and x22 and x68 and x7 and x8 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and not x21 and x22 and x68 and x7 and not x8 and x9 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and not x21 and x22 and x68 and x7 and not x8 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and x68 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and not x68 and x23 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and not x21 and x22 and not x68 and x23 and x17 and not x14 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and not x21 and x22 and not x68 and x23 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and not x68 and x23 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and not x68 and not x23 and x18 and x14 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x21 and x22 and not x68 and not x23 and x18 and not x14 and x13 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x21 and x22 and not x68 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and not x68 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and not x22 and x68 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and not x21 and not x22 and not x68 and x23 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s330;

      else
         y3 <= '1' ;
         y4 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s333;

      end if;

   when s87 =>
      if ( x21 and x19 and x15 and x10 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s330;

      elsif ( x21 and x19 and x15 and not x10 and x12 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( x21 and x19 and x15 and not x10 and not x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s48;

      elsif ( x21 and x19 and not x15 and x16 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x21 and x19 and not x15 and not x16 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s340;

      elsif ( x21 and not x19 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s84;

      elsif ( not x21 and x23 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x23 and x22 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s84;

      else
         current_group15m <= s1;

      end if;

   when s88 =>
      if ( x21 and x66 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x21 and x66 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x21 and x66 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x66 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x66 and x19 and x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s272;

      elsif ( x21 and not x66 and x19 and not x12 and x17 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s272;

      elsif ( x21 and not x66 and x19 and not x12 and not x17 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s273;

      elsif ( x21 and not x66 and not x19 and x20 and x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s272;

      elsif ( x21 and not x66 and not x19 and x20 and not x12 ) = '1' then
         y10 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s273;

      elsif ( x21 and not x66 and not x19 and not x20 and x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s270;

      elsif ( x21 and not x66 and not x19 and not x20 and not x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s109;

      elsif ( not x21 and x66 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x66 and x22 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      else
         current_group15m <= s1;

      end if;

   when s89 =>
      if ( x66 and x65 and x61 and x60 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and x65 and x61 and not x60 and x62 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and x61 and not x60 and not x62 and x15 and x12 and x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x66 and x65 and x61 and not x60 and not x62 and x15 and x12 and not x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s250;

      elsif ( x66 and x65 and x61 and not x60 and not x62 and x15 and not x12 and x7 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x66 and x65 and x61 and not x60 and not x62 and x15 and not x12 and not x7 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s262;

      elsif ( x66 and x65 and x61 and not x60 and not x62 and not x15 and x16 and x7 and x12 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s251;

      elsif ( x66 and x65 and x61 and not x60 and not x62 and not x15 and x16 and x7 and not x12 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s252;

      elsif ( x66 and x65 and x61 and not x60 and not x62 and not x15 and x16 and not x7 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s252;

      elsif ( x66 and x65 and x61 and not x60 and not x62 and not x15 and not x16 and x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s253;

      elsif ( x66 and x65 and x61 and not x60 and not x62 and not x15 and not x16 and not x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x66 and x65 and not x61 and x60 and x15 and x12 and x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x66 and x65 and not x61 and x60 and x15 and x12 and not x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s250;

      elsif ( x66 and x65 and not x61 and x60 and x15 and not x12 and x7 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x66 and x65 and not x61 and x60 and x15 and not x12 and not x7 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s262;

      elsif ( x66 and x65 and not x61 and x60 and not x15 and x16 and x7 and x12 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s251;

      elsif ( x66 and x65 and not x61 and x60 and not x15 and x16 and x7 and not x12 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s252;

      elsif ( x66 and x65 and not x61 and x60 and not x15 and x16 and not x7 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s252;

      elsif ( x66 and x65 and not x61 and x60 and not x15 and not x16 and x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s253;

      elsif ( x66 and x65 and not x61 and x60 and not x15 and not x16 and not x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x66 and x65 and not x61 and not x60 and x62 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( x66 and x65 and not x61 and not x60 and not x62 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and not x65 and x67 and x62 and x61 and x13 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x66 and not x65 and x67 and x62 and x61 and not x13 and x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x66 and not x65 and x67 and x62 and x61 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and x67 and x62 and not x61 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and x67 and not x62 and x63 and x17 and x13 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and not x65 and x67 and not x62 and x63 and x17 and x13 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( x66 and not x65 and x67 and not x62 and x63 and x17 and not x13 and x12 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and not x65 and x67 and not x62 and x63 and x17 and not x13 and x12 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( x66 and not x65 and x67 and not x62 and x63 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and x67 and not x62 and x63 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and x67 and not x62 and not x63 and x19 and x13 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x66 and not x65 and x67 and not x62 and not x63 and x19 and x13 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x66 and not x65 and x67 and not x62 and not x63 and x19 and not x13 and x12 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x66 and not x65 and x67 and not x62 and not x63 and x19 and not x13 and x12 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x66 and not x65 and x67 and not x62 and not x63 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and x67 and not x62 and not x63 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and x21 and x68 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x66 and not x65 and not x67 and x21 and x68 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x66 and not x65 and not x67 and x21 and x68 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and x21 and x68 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and x21 and not x68 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x66 and not x65 and not x67 and x21 and not x68 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x66 and not x65 and not x67 and x21 and not x68 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and x21 and not x68 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and x22 and x68 and x7 and x8 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( x66 and not x65 and not x67 and not x21 and x22 and x68 and x7 and not x8 and x9 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( x66 and not x65 and not x67 and not x21 and x22 and x68 and x7 and not x8 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and x22 and x68 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and x22 and not x68 and x23 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( x66 and not x65 and not x67 and not x21 and x22 and not x68 and x23 and x17 and not x14 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( x66 and not x65 and not x67 and not x21 and x22 and not x68 and x23 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and x22 and not x68 and x23 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and x22 and not x68 and not x23 and x18 and x14 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and not x65 and not x67 and not x21 and x22 and not x68 and not x23 and x18 and not x14 and x13 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and not x65 and not x67 and not x21 and x22 and not x68 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and x22 and not x68 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and not x22 and x68 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x65 and not x67 and not x21 and not x22 and x68 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x66 and not x65 and not x67 and not x21 and not x22 and x68 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and not x22 and x68 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and not x22 and not x68 and x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x66 and not x65 and not x67 and not x21 and not x22 and not x68 and not x23 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x66 and x65 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and x24 and x26 and x18 and x15 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x66 and not x65 and x67 and x24 and x26 and x18 and not x15 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x66 and not x65 and x67 and x24 and x26 and x18 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and x24 and x26 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and x24 and not x26 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x66 and not x65 and x67 and x24 and not x26 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x66 and not x65 and x67 and x24 and not x26 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and x24 and not x26 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and not x24 and x25 and x26 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x66 and not x65 and x67 and not x24 and x25 and x26 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x66 and not x65 and x67 and not x24 and x25 and x26 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s89;

      elsif ( not x66 and not x65 and x67 and not x24 and x25 and x26 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and not x24 and x25 and not x26 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and x26 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and x26 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and x26 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and x26 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and not x26 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and not x26 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and not x26 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and not x26 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x67 and x21 and x19 and x17 and x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s272;

      elsif ( not x66 and not x65 and not x67 and x21 and x19 and x17 and not x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s272;

      elsif ( not x66 and not x65 and not x67 and x21 and x19 and not x17 and x12 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and not x65 and not x67 and x21 and x19 and not x17 and not x12 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s273;

      elsif ( not x66 and not x65 and not x67 and x21 and not x19 and x20 and x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s272;

      elsif ( not x66 and not x65 and not x67 and x21 and not x19 and x20 and not x12 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s105;

      elsif ( not x66 and not x65 and not x67 and x21 and not x19 and not x20 and x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s270;

      elsif ( not x66 and not x65 and not x67 and x21 and not x19 and not x20 and not x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s109;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and x12 and x4 and x18 and x17 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s203;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and x12 and x4 and x18 and not x17 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s275;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and x12 and x4 and not x18 and x19 and x17 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s272;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and x12 and x4 and not x18 and x19 and not x17 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s275;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and x12 and x4 and not x18 and not x19 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s272;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and x12 and not x4 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s275;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and x18 and x4 and x17 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s234;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and x18 and x4 and not x17 ) = '1' then
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s273;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and x18 and not x4 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s275;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and not x18 and x19 and x17 and x14 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s275;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and not x18 and x19 and x17 and not x14 and x16 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s275;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and not x18 and x19 and x17 and not x14 and not x16 and x6 and x7 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and not x18 and x19 and x17 and not x14 and not x16 and x6 and not x7 and x8 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and not x18 and x19 and x17 and not x14 and not x16 and x6 and not x7 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and not x18 and x19 and x17 and not x14 and not x16 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and not x18 and x19 and not x17 and x16 and x15 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s275;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and not x18 and x19 and not x17 and x16 and not x15 and x6 and x7 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and not x18 and x19 and not x17 and x16 and not x15 and x6 and not x7 and x8 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and not x18 and x19 and not x17 and x16 and not x15 and x6 and not x7 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and not x18 and x19 and not x17 and x16 and not x15 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and not x18 and x19 and not x17 and not x16 and x13 and x6 and x7 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and not x18 and x19 and not x17 and not x16 and x13 and x6 and not x7 and x8 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and not x18 and x19 and not x17 and not x16 and x13 and x6 and not x7 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and not x18 and x19 and not x17 and not x16 and x13 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and not x18 and x19 and not x17 and not x16 and not x13 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s275;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and not x18 and not x19 and x4 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x66 and not x65 and not x67 and not x21 and x22 and not x12 and not x18 and not x19 and not x4 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s275;

      elsif ( not x66 and not x65 and not x67 and not x21 and not x22 and x15 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x66 and not x65 and not x67 and not x21 and not x22 and not x15 and x19 and x18 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x66 and not x65 and not x67 and not x21 and not x22 and not x15 and x19 and not x18 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s342;

      else
         y5 <= '1' ;
         current_group15m <= s101;

      end if;

   when s90 =>
         y2 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s364;

   when s91 =>
      if ( x65 and x21 and x18 and x20 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( x65 and x21 and x18 and not x20 ) = '1' then
         current_group15m <= s91;

      elsif ( x65 and x21 and not x18 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x21 and x22 and x15 and x9 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x65 and not x21 and x22 and x15 and not x9 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x65 and not x21 and x22 and not x15 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s205;

      elsif ( x65 and not x21 and not x22 and x23 and x20 and x14 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x21 and not x22 and x23 and x20 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x21 and not x22 and x23 and x20 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x22 and x23 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and x14 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x21 and not x22 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x22 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and x68 and x21 and x19 and x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and x67 and x66 and x68 and x21 and x19 and not x15 and x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and x67 and x66 and x68 and x21 and x19 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and x68 and x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and x68 and not x21 and x20 and x15 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( not x65 and x67 and x66 and x68 and not x21 and x20 and not x15 and x14 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( not x65 and x67 and x66 and x68 and not x21 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and x68 and not x21 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and x15 and x14 and x8 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and x15 and x14 and not x8 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and x15 and not x14 and x7 and x8 ) = '1' then
         y24 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s157;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and x15 and not x14 and x7 and not x8 ) = '1' then
         y26 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s158;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and x15 and not x14 and not x7 and x8 and x12 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s65;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and x15 and not x14 and not x7 and x8 and not x12 and x17 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and x15 and not x14 and not x7 and x8 and not x12 and x17 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and x15 and not x14 and not x7 and x8 and not x12 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and x15 and not x14 and not x7 and not x8 and x13 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s65;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and x15 and not x14 and not x7 and not x8 and not x13 and x17 and x12 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and x15 and not x14 and not x7 and not x8 and not x13 and x17 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and x15 and not x14 and not x7 and not x8 and not x13 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and x2 and x8 and x7 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and x2 and x8 and not x7 and x9 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and x2 and x8 and not x7 and not x9 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and x2 and not x8 and x7 and x11 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and x2 and not x8 and x7 and not x11 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and x2 and not x8 and not x7 and x10 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and x2 and not x8 and not x7 and not x10 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and not x2 and x7 and x8 and x1 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and not x2 and x7 and x8 and not x1 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and not x2 and x7 and not x8 and x11 and x1 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and not x2 and x7 and not x8 and x11 and not x1 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and not x2 and x7 and not x8 and not x11 and x17 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and not x2 and x7 and not x8 and not x11 and x17 and not x13 and x12 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and not x2 and x7 and not x8 and not x11 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and not x2 and x7 and not x8 and not x11 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and not x2 and not x7 and x8 and x9 and x1 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and not x2 and not x7 and x8 and x9 and not x1 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and not x2 and not x7 and x8 and not x9 and x17 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and not x2 and not x7 and x8 and not x9 and x17 and not x13 and x12 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and not x2 and not x7 and x8 and not x9 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and not x2 and not x7 and x8 and not x9 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and not x2 and not x7 and not x8 and x10 and x1 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and not x2 and not x7 and not x8 and x10 and not x1 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and not x2 and not x7 and not x8 and not x10 and x17 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and not x2 and not x7 and not x8 and not x10 and x17 and not x13 and x12 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and not x2 and not x7 and not x8 and not x10 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and x16 and not x15 and not x2 and not x7 and not x8 and not x10 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and not x16 and x15 and x7 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s159;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and not x16 and x15 and not x7 and x2 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and not x16 and x15 and not x7 and not x2 and x1 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and not x16 and x15 and not x7 and not x2 and not x1 and x8 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and not x16 and x15 and not x7 and not x2 and not x1 and not x8 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s203;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and not x16 and not x15 and x2 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and not x16 and not x15 and not x2 and x1 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and x64 and not x16 and not x15 and not x2 and not x1 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s135;

      elsif ( not x65 and x67 and x66 and not x68 and x63 and not x64 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and x16 and x8 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and x16 and not x8 and x6 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and x16 and not x8 and not x6 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and not x16 and x4 and x8 and x7 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and not x16 and x4 and x8 and not x7 and x9 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and not x16 and x4 and x8 and not x7 and not x9 and x19 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and not x16 and x4 and x8 and not x7 and not x9 and x19 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and not x16 and x4 and x8 and not x7 and not x9 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and not x16 and x4 and x8 and not x7 and not x9 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and not x16 and x4 and not x8 and x7 and x11 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and not x16 and x4 and not x8 and x7 and not x11 and x19 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and not x16 and x4 and not x8 and x7 and not x11 and x19 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and not x16 and x4 and not x8 and x7 and not x11 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and not x16 and x4 and not x8 and x7 and not x11 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and not x16 and x4 and not x8 and not x7 and x10 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and not x16 and x4 and not x8 and not x7 and not x10 and x19 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and not x16 and x4 and not x8 and not x7 and not x10 and x19 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and not x16 and x4 and not x8 and not x7 and not x10 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and not x16 and x4 and not x8 and not x7 and not x10 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and not x16 and not x4 and x6 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s135;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and x64 and not x16 and not x4 and not x6 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and not x64 and x19 and x13 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and not x64 and x19 and not x13 and x12 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and not x64 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x66 and not x68 and not x63 and not x64 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and not x66 and x24 and x26 and x16 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x67 and not x66 and x24 and x26 and not x16 and x17 and x13 and x11 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x67 and not x66 and x24 and x26 and not x16 and x17 and x13 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s282;

      elsif ( not x65 and x67 and not x66 and x24 and x26 and not x16 and x17 and x13 and not x11 and not x12 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x67 and not x66 and x24 and x26 and not x16 and x17 and not x13 and x11 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s17;

      elsif ( not x65 and x67 and not x66 and x24 and x26 and not x16 and x17 and not x13 and not x11 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x67 and not x66 and x24 and x26 and not x16 and not x17 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s51;

      elsif ( not x65 and x67 and not x66 and x24 and not x26 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x65 and x67 and not x66 and not x24 and x25 and x26 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and x67 and not x66 and not x24 and x25 and x26 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and x67 and not x66 and not x24 and x25 and x26 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s91;

      elsif ( not x65 and x67 and not x66 and not x24 and x25 and x26 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and not x66 and not x24 and x25 and not x26 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and x67 and not x66 and not x24 and not x25 and x26 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      elsif ( not x65 and x67 and not x66 and not x24 and not x25 and not x26 and x15 and x12 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and x67 and not x66 and not x24 and not x25 and not x26 and x15 and not x12 and x11 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and x67 and not x66 and not x24 and not x25 and not x26 and x15 and not x12 and not x11 and x10 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and x67 and not x66 and not x24 and not x25 and not x26 and x15 and not x12 and not x11 and not x10 ) = '1' then
         y12 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s49;

      elsif ( not x65 and x67 and not x66 and not x24 and not x25 and not x26 and not x15 and x16 and x10 and x12 ) = '1' then
         y15 <= '1' ;
         y112 <= '1' ;
         current_group15m <= s46;

      elsif ( not x65 and x67 and not x66 and not x24 and not x25 and not x26 and not x15 and x16 and x10 and not x12 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and x67 and not x66 and not x24 and not x25 and not x26 and not x15 and x16 and not x10 ) = '1' then
         y15 <= '1' ;
         y112 <= '1' ;
         current_group15m <= s46;

      elsif ( not x65 and x67 and not x66 and not x24 and not x25 and not x26 and not x15 and not x16 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x67 and x66 and x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and x66 and not x21 and x22 and x7 and x8 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and not x67 and x66 and not x21 and x22 and x7 and not x8 and x9 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and not x67 and x66 and not x21 and x22 and x7 and not x8 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and x66 and not x21 and x22 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and x66 and not x21 and not x22 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and not x67 and x66 and not x21 and not x22 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and not x67 and x66 and not x21 and not x22 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x66 and x3 and x4 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( not x65 and not x67 and not x66 and x3 and not x4 and x5 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( not x65 and not x67 and not x66 and x3 and not x4 and not x5 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s92 =>
      if ( x65 and x67 and x21 ) = '1' then
         y8 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s365;

      elsif ( x65 and x67 and not x21 and x23 and x22 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x21 and x23 and x22 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x21 and x23 and x22 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x21 and x23 and x22 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x21 and x23 and not x22 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x21 and x23 and not x22 and x9 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x21 and x23 and not x22 and x9 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x21 and x23 and not x22 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x21 and not x23 and x8 and x22 and x9 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x21 and not x23 and x8 and x22 and not x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x21 and not x23 and x8 and x22 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x21 and not x23 and x8 and not x22 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x21 and not x23 and x8 and not x22 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and not x21 and not x23 and x8 and not x22 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x21 and not x23 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x68 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x67 and x68 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x67 and x68 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x68 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x68 and x21 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and x23 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and x23 and not x19 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and x23 and not x19 and x17 and not x14 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and x23 and not x19 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and x23 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and x15 and x16 and x7 and x9 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and x15 and x16 and x7 and not x9 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and x15 and x16 and not x7 and x8 and x9 ) = '1' then
         y24 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s157;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and x15 and x16 and not x7 and x8 and not x9 ) = '1' then
         y26 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s158;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and x15 and x16 and not x7 and not x8 and x9 and x13 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s191;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and x15 and x16 and not x7 and not x8 and x9 and not x13 and x18 and x14 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and x15 and x16 and not x7 and not x8 and x9 and not x13 and x18 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and x15 and x16 and not x7 and not x8 and x9 and not x13 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and x15 and x16 and not x7 and not x8 and not x9 and x14 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s191;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and x15 and x16 and not x7 and not x8 and not x9 and not x14 and x18 and x13 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and x15 and x16 and not x7 and not x8 and not x9 and not x14 and x18 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and x15 and x16 and not x7 and not x8 and not x9 and not x14 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and x15 and not x16 and x7 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and x15 and not x16 and not x7 and x8 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and x15 and not x16 and not x7 and not x8 and x1 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s22;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and x15 and not x16 and not x7 and not x8 and not x1 and x5 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and x15 and not x16 and not x7 and not x8 and not x1 and not x5 and x9 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and x15 and not x16 and not x7 and not x8 and not x1 and not x5 and not x9 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and not x15 and x1 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s22;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and not x15 and not x1 and x16 and x9 and x10 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and not x15 and not x1 and x16 and x9 and not x10 and x8 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and not x15 and not x1 and x16 and x9 and not x10 and not x8 and x18 and x14 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and not x15 and not x1 and x16 and x9 and not x10 and not x8 and x18 and not x14 and x13 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and not x15 and not x1 and x16 and x9 and not x10 and not x8 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and not x15 and not x1 and x16 and x9 and not x10 and not x8 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and not x15 and not x1 and x16 and not x9 and x8 and x12 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and not x15 and not x1 and x16 and not x9 and x8 and not x12 and x18 and x14 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and not x15 and not x1 and x16 and not x9 and x8 and not x12 and x18 and not x14 and x13 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and not x15 and not x1 and x16 and not x9 and x8 and not x12 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and not x15 and not x1 and x16 and not x9 and x8 and not x12 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and not x15 and not x1 and x16 and not x9 and not x8 and x11 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and not x15 and not x1 and x16 and not x9 and not x8 and not x11 and x18 and x14 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and not x15 and not x1 and x16 and not x9 and not x8 and not x11 and x18 and not x14 and x13 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and not x15 and not x1 and x16 and not x9 and not x8 and not x11 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and not x15 and not x1 and x16 and not x9 and not x8 and not x11 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and not x15 and not x1 and not x16 and x5 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x67 and not x68 and not x21 and x22 and not x23 and not x15 and not x1 and not x16 and not x5 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s205;

      elsif ( x65 and not x67 and not x68 and not x21 and not x22 and x4 and x18 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x67 and not x68 and not x21 and not x22 and x4 and not x18 and x19 ) = '1' then
         current_group15m <= s92;

      elsif ( x65 and not x67 and not x68 and not x21 and not x22 and x4 and not x18 and not x19 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s97;

      elsif ( x65 and not x67 and not x68 and not x21 and not x22 and not x4 and x3 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and not x67 and not x68 and not x21 and not x22 and not x4 and not x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      elsif ( not x65 and x66 and x68 and x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x68 and not x21 and x16 and x10 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s67;

      elsif ( not x65 and x66 and x68 and not x21 and x16 and not x10 ) = '1' then
         y5 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s113;

      elsif ( not x65 and x66 and x68 and not x21 and not x16 ) = '1' then
         y5 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s115;

      elsif ( not x65 and x66 and not x68 and x63 and x64 and x6 and x15 and x8 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s298;

      elsif ( not x65 and x66 and not x68 and x63 and x64 and x6 and x15 and not x8 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x65 and x66 and not x68 and x63 and x64 and x6 and not x15 and x16 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s298;

      elsif ( not x65 and x66 and not x68 and x63 and x64 and x6 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s204;

      elsif ( not x65 and x66 and not x68 and x63 and x64 and not x6 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s298;

      elsif ( not x65 and x66 and not x68 and x63 and not x64 and x5 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s20;

      elsif ( not x65 and x66 and not x68 and x63 and not x64 and not x5 and x18 and x15 and x8 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and x66 and not x68 and x63 and not x64 and not x5 and x18 and x15 and not x8 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x65 and x66 and not x68 and x63 and not x64 and not x5 and x18 and not x15 and x16 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( not x65 and x66 and not x68 and x63 and not x64 and not x5 and x18 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s135;

      elsif ( not x65 and x66 and not x68 and x63 and not x64 and not x5 and not x18 ) = '1' then
         y31 <= '1' ;
         current_group15m <= s96;

      elsif ( not x65 and x66 and not x68 and not x63 and x64 and x19 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x66 and not x68 and not x63 and x64 and x19 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x66 and not x68 and not x63 and x64 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x68 and not x63 and x64 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x68 and not x63 and not x64 and x4 ) = '1' then
         y31 <= '1' ;
         current_group15m <= s96;

      elsif ( not x65 and x66 and not x68 and not x63 and not x64 and not x4 and x17 and x15 and x8 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x65 and x66 and not x68 and not x63 and not x64 and not x4 and x17 and x15 and not x8 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x65 and x66 and not x68 and not x63 and not x64 and not x4 and x17 and not x15 and x16 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s151;

      elsif ( not x65 and x66 and not x68 and not x63 and not x64 and not x4 and x17 and not x15 and not x16 and x14 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s135;

      elsif ( not x65 and x66 and not x68 and not x63 and not x64 and not x4 and x17 and not x15 and not x16 and not x14 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s152;

      elsif ( not x65 and x66 and not x68 and not x63 and not x64 and not x4 and not x17 ) = '1' then
         y14 <= '1' ;
         y28 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_group15m <= s18;

      elsif ( not x65 and not x66 and x67 and x68 and x20 and x18 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x66 and x67 and x68 and x20 and x18 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x66 and x67 and x68 and x20 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x68 and x20 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x68 and not x20 and x21 and x3 ) = '1' then
         y2 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s366;

      elsif ( not x65 and not x66 and x67 and x68 and not x20 and x21 and not x3 and x17 and x15 and x8 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s254;

      elsif ( not x65 and not x66 and x67 and x68 and not x20 and x21 and not x3 and x17 and x15 and not x8 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s198;

      elsif ( not x65 and not x66 and x67 and x68 and not x20 and x21 and not x3 and x17 and not x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x65 and not x66 and x67 and x68 and not x20 and x21 and not x3 and x17 and not x15 and not x16 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s209;

      elsif ( not x65 and not x66 and x67 and x68 and not x20 and x21 and not x3 and not x17 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x66 and x67 and x68 and not x20 and not x21 and x15 and x8 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x66 and x67 and x68 and not x20 and not x21 and x15 and not x8 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s198;

      elsif ( not x65 and not x66 and x67 and x68 and not x20 and not x21 and not x15 and x16 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s59;

      elsif ( not x65 and not x66 and x67 and x68 and not x20 and not x21 and not x15 and not x16 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s209;

      elsif ( not x65 and not x66 and x67 and not x68 and x24 and x26 and x16 and x18 and x15 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and not x66 and x67 and not x68 and x24 and x26 and x16 and x18 and not x15 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and not x66 and x67 and not x68 and x24 and x26 and x16 and x18 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and not x68 and x24 and x26 and x16 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and not x68 and x24 and x26 and not x16 ) = '1' then
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s165;

      elsif ( not x65 and not x66 and x67 and not x68 and x24 and not x26 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and not x66 and x67 and not x68 and x24 and not x26 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x65 and not x66 and x67 and not x68 and x24 and not x26 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and not x68 and x24 and not x26 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and not x68 and not x24 and x25 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and x67 and not x68 and not x24 and x25 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and x67 and not x68 and not x24 and x25 and x19 and not x14 and not x13 and x26 ) = '1' then
         current_group15m <= s92;

      elsif ( not x65 and not x66 and x67 and not x68 and not x24 and x25 and x19 and not x14 and not x13 and not x26 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and not x68 and not x24 and x25 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and not x68 and not x24 and not x25 and x26 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s17;

      elsif ( not x65 and not x66 and x67 and not x68 and not x24 and not x25 and not x26 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x65 and not x66 and x67 and not x68 and not x24 and not x25 and not x26 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x65 and not x66 and x67 and not x68 and not x24 and not x25 and not x26 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and not x68 and not x24 and not x25 and not x26 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and x68 and x3 and x4 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( not x65 and not x66 and not x67 and x68 and x3 and not x4 and x5 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( not x65 and not x66 and not x67 and x68 and x3 and not x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and x68 and not x3 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and not x68 and x21 and x9 and x3 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x66 and not x67 and not x68 and x21 and x9 and not x3 and x4 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x66 and not x67 and not x68 and x21 and x9 and not x3 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and not x68 and x21 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x5 and not x4 and x22 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x5 and not x4 and x22 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and x5 and not x4 and not x22 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and not x5 and x22 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and not x5 and not x22 and x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x67 and not x68 and not x21 and not x5 and not x22 and x4 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s93 =>
      if ( x22 and x20 and x19 ) = '1' then
         y1 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s93;

      elsif ( x22 and x20 and not x19 and x23 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x22 and x20 and not x19 and not x23 ) = '1' then
         current_group15m <= s93;

      elsif ( x22 and not x20 and x23 and x19 ) = '1' then
         current_group15m <= s93;

      elsif ( x22 and not x20 and x23 and not x19 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x22 and not x20 and not x23 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      else
         y25 <= '1' ;
         current_group15m <= s78;

      end if;

   when s94 =>
      if ( x22 and x4 and x19 ) = '1' then
         y1 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s93;

      elsif ( x22 and x4 and not x19 and x20 ) = '1' then
         current_group15m <= s94;

      elsif ( x22 and x4 and not x19 and not x20 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x22 and not x4 and x3 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x22 and not x4 and not x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s24;

      else
         y8 <= '1' ;
         y16 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s1;

      end if;

   when s95 =>
      if ( x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and x18 and x15 and x9 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x21 and x22 and x23 and x18 and x15 and not x9 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x21 and x22 and x23 and x18 and not x15 and x16 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x21 and x22 and x23 and x18 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s205;

      elsif ( not x21 and x22 and x23 and not x18 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s97;

      elsif ( not x21 and x22 and not x23 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s97;

      elsif ( not x21 and not x22 and x23 and x15 and x9 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x21 and not x22 and x23 and x15 and not x9 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x21 and not x22 and x23 and not x15 and x16 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and x23 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s205;

      else
         current_group15m <= s1;

      end if;

   when s96 =>
      if ( x65 and x21 and x17 and x15 and x9 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( x65 and x21 and x17 and x15 and not x9 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( x65 and x21 and x17 and not x15 and x16 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x65 and x21 and x17 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s212;

      elsif ( x65 and x21 and not x17 ) = '1' then
         y15 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_group15m <= s294;

      elsif ( x65 and not x21 and x23 ) = '1' then
         y15 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_group15m <= s294;

      elsif ( x65 and not x21 and not x23 and x22 and x5 ) = '1' then
         y15 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_group15m <= s294;

      elsif ( x65 and not x21 and not x23 and x22 and not x5 and x17 and x15 and x9 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x21 and not x23 and x22 and not x5 and x17 and x15 and not x9 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x65 and not x21 and not x23 and x22 and not x5 and x17 and not x15 and x16 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and not x23 and x22 and not x5 and x17 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s205;

      elsif ( x65 and not x21 and not x23 and x22 and not x5 and not x17 ) = '1' then
         y35 <= '1' ;
         current_group15m <= s26;

      elsif ( x65 and not x21 and not x23 and not x22 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s147;

      elsif ( not x65 and x63 ) = '1' then
         y14 <= '1' ;
         y28 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_group15m <= s18;

      elsif ( not x65 and not x63 and x64 and x18 and x16 and x8 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and not x63 and x64 and x18 and x16 and not x8 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x65 and not x63 and x64 and x18 and not x16 and x4 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( not x65 and not x63 and x64 and x18 and not x16 and not x4 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s135;

      elsif ( not x65 and not x63 and x64 and not x18 ) = '1' then
         y14 <= '1' ;
         y28 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_group15m <= s18;

      elsif ( not x65 and not x63 and not x64 and x17 and x15 and x8 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x65 and not x63 and not x64 and x17 and x15 and not x8 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x65 and not x63 and not x64 and x17 and not x15 and x16 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s151;

      elsif ( not x65 and not x63 and not x64 and x17 and not x15 and not x16 and x14 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s135;

      elsif ( not x65 and not x63 and not x64 and x17 and not x15 and not x16 and not x14 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s152;

      else
         y14 <= '1' ;
         y28 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_group15m <= s18;

      end if;

   when s97 =>
      if ( x23 and x22 ) = '1' then
         y2 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s98;

      elsif ( x23 and not x22 ) = '1' then
         current_group15m <= s1;

      elsif ( not x23 and x22 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s298;

      elsif ( not x23 and not x22 and x4 and x20 ) = '1' then
         y2 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s98;

      elsif ( not x23 and not x22 and x4 and not x20 and x19 ) = '1' then
         current_group15m <= s97;

      elsif ( not x23 and not x22 and x4 and not x20 and not x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( not x23 and not x22 and not x4 and x3 ) = '1' then
         y1 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s93;

      else
         y1 <= '1' ;
         current_group15m <= s24;

      end if;

   when s98 =>
      if ( x22 and x15 and x9 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x22 and x15 and not x9 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x22 and not x15 and x16 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x22 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s205;

      elsif ( not x22 and x19 and x20 ) = '1' then
         y2 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s98;

      elsif ( not x22 and x19 and not x20 ) = '1' then
         current_group15m <= s98;

      else
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      end if;

   when s99 =>
      if ( x23 and x22 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x23 and x22 and x17 and not x14 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x23 and x22 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x23 and x22 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x23 and not x22 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s100 =>
      if ( x65 and x66 and x67 and x23 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and x66 and x67 and x23 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and x66 and x67 and x23 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x67 and x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x67 and not x23 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x65 and x66 and not x67 and x61 and x60 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x66 and not x67 and x61 and x60 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x66 and not x67 and x61 and x60 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x66 and not x67 and x61 and x60 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x66 and not x67 and x61 and not x60 and x62 and x2 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( x65 and x66 and not x67 and x61 and not x60 and x62 and not x2 and x20 ) = '1' then
         y2 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s367;

      elsif ( x65 and x66 and not x67 and x61 and not x60 and x62 and not x2 and not x20 and x16 and x11 and x12 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s153;

      elsif ( x65 and x66 and not x67 and x61 and not x60 and x62 and not x2 and not x20 and x16 and x11 and not x12 and x13 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s153;

      elsif ( x65 and x66 and not x67 and x61 and not x60 and x62 and not x2 and not x20 and x16 and x11 and not x12 and not x13 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s154;

      elsif ( x65 and x66 and not x67 and x61 and not x60 and x62 and not x2 and not x20 and x16 and not x11 and x13 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s63;

      elsif ( x65 and x66 and not x67 and x61 and not x60 and x62 and not x2 and not x20 and x16 and not x11 and not x13 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( x65 and x66 and not x67 and x61 and not x60 and x62 and not x2 and not x20 and not x16 and x17 and x11 and x13 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x65 and x66 and not x67 and x61 and not x60 and x62 and not x2 and not x20 and not x16 and x17 and x11 and not x13 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( x65 and x66 and not x67 and x61 and not x60 and x62 and not x2 and not x20 and not x16 and x17 and not x11 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x65 and x66 and not x67 and x61 and not x60 and x62 and not x2 and not x20 and not x16 and not x17 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( x65 and x66 and not x67 and x61 and not x60 and not x62 and x7 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x65 and x66 and not x67 and x61 and not x60 and not x62 and not x7 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x66 and not x67 and not x61 and x60 and x7 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x65 and x66 and not x67 and not x61 and x60 and not x7 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x66 and not x67 and not x61 and not x60 and x62 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( x65 and x66 and not x67 and not x61 and not x60 and not x62 ) = '1' then
         current_group15m <= s316;

      elsif ( x65 and not x66 and x21 and x18 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x65 and not x66 and x21 and not x18 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x21 and not x18 and x19 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and x21 and not x18 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x21 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and x15 and x9 ) = '1' then
         y31 <= '1' ;
         current_group15m <= s96;

      elsif ( x65 and not x66 and not x21 and x22 and x15 and not x9 and x6 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( x65 and not x66 and not x21 and x22 and x15 and not x9 and not x6 ) = '1' then
         y31 <= '1' ;
         current_group15m <= s96;

      elsif ( x65 and not x66 and not x21 and x22 and not x15 and x16 and x9 and x8 ) = '1' then
         y31 <= '1' ;
         current_group15m <= s96;

      elsif ( x65 and not x66 and not x21 and x22 and not x15 and x16 and x9 and not x8 and x10 ) = '1' then
         y31 <= '1' ;
         current_group15m <= s96;

      elsif ( x65 and not x66 and not x21 and x22 and not x15 and x16 and x9 and not x8 and not x10 and x18 and x14 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x21 and x22 and not x15 and x16 and x9 and not x8 and not x10 and x18 and not x14 and x13 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x21 and x22 and not x15 and x16 and x9 and not x8 and not x10 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x15 and x16 and x9 and not x8 and not x10 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x15 and x16 and not x9 and x8 and x12 ) = '1' then
         y31 <= '1' ;
         current_group15m <= s96;

      elsif ( x65 and not x66 and not x21 and x22 and not x15 and x16 and not x9 and x8 and not x12 and x18 and x14 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x21 and x22 and not x15 and x16 and not x9 and x8 and not x12 and x18 and not x14 and x13 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x21 and x22 and not x15 and x16 and not x9 and x8 and not x12 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x15 and x16 and not x9 and x8 and not x12 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x15 and x16 and not x9 and not x8 and x11 ) = '1' then
         y31 <= '1' ;
         current_group15m <= s96;

      elsif ( x65 and not x66 and not x21 and x22 and not x15 and x16 and not x9 and not x8 and not x11 and x18 and x14 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x21 and x22 and not x15 and x16 and not x9 and not x8 and not x11 and x18 and not x14 and x13 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x21 and x22 and not x15 and x16 and not x9 and not x8 and not x11 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x15 and x16 and not x9 and not x8 and not x11 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x15 and not x16 and x6 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s212;

      elsif ( x65 and not x66 and not x21 and x22 and not x15 and not x16 and not x6 ) = '1' then
         y31 <= '1' ;
         current_group15m <= s96;

      elsif ( x65 and not x66 and not x21 and not x22 ) = '1' then
         y31 <= '1' ;
         current_group15m <= s96;

      elsif ( not x65 and x66 and x21 and x68 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x21 and not x68 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x65 and x66 and x21 and not x68 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x65 and x66 and x21 and not x68 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x21 and not x68 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x21 and x22 and x68 and x17 and x10 and x15 and x6 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s283;

      elsif ( not x65 and x66 and not x21 and x22 and x68 and x17 and x10 and x15 and not x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and x66 and not x21 and x22 and x68 and x17 and x10 and not x15 and x16 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( not x65 and x66 and not x21 and x22 and x68 and x17 and x10 and not x15 and not x16 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and x66 and not x21 and x22 and x68 and x17 and not x10 and x6 ) = '1' then
         y13 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s284;

      elsif ( not x65 and x66 and not x21 and x22 and x68 and x17 and not x10 and not x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and x66 and not x21 and x22 and x68 and not x17 and x18 and x6 and x10 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s219;

      elsif ( not x65 and x66 and not x21 and x22 and x68 and not x17 and x18 and x6 and not x10 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( not x65 and x66 and not x21 and x22 and x68 and not x17 and x18 and not x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and x66 and not x21 and x22 and x68 and not x17 and not x18 and x6 and x10 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s219;

      elsif ( not x65 and x66 and not x21 and x22 and x68 and not x17 and not x18 and x6 and not x10 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s28;

      elsif ( not x65 and x66 and not x21 and x22 and x68 and not x17 and not x18 and not x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x66 and not x21 and x22 and not x68 and x23 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x65 and x66 and not x21 and x22 and not x68 and not x23 and x18 and x14 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and x66 and not x21 and x22 and not x68 and not x23 and x18 and not x14 and x13 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and x66 and not x21 and x22 and not x68 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x21 and x22 and not x68 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x21 and not x22 and x68 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x66 and not x21 and not x22 and x68 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x66 and not x21 and not x22 and x68 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x21 and not x22 and x68 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x21 and not x22 and not x68 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x20 and x18 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x66 and x67 and x20 and x18 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x66 and x67 and x20 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x20 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and not x20 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x65 and not x66 and not x67 and x21 and x9 and x3 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x66 and not x67 and x21 and x9 and not x3 and x4 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x66 and not x67 and x21 and x9 and not x3 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and x21 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x5 and not x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x5 and not x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and not x5 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s101 =>
      if ( x65 and x66 and x22 and x20 and x15 and x8 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x66 and x22 and x20 and x15 and not x8 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x65 and x66 and x22 and x20 and not x15 and x16 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s302;

      elsif ( x65 and x66 and x22 and x20 and not x15 and not x16 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s122;

      elsif ( x65 and x66 and x22 and not x20 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s368;

      elsif ( x65 and x66 and not x22 and x23 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x22 and not x23 and x3 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s368;

      elsif ( x65 and x66 and not x22 and not x23 and not x3 and x19 and x15 and x8 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s8;

      elsif ( x65 and x66 and not x22 and not x23 and not x3 and x19 and x15 and not x8 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s111;

      elsif ( x65 and x66 and not x22 and not x23 and not x3 and x19 and not x15 and x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s50;

      elsif ( x65 and x66 and not x22 and not x23 and not x3 and x19 and not x15 and not x16 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( x65 and x66 and not x22 and not x23 and not x3 and not x19 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s314;

      elsif ( x65 and not x66 and x68 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x68 and x21 and x5 ) = '1' then
         y31 <= '1' ;
         current_group15m <= s96;

      elsif ( x65 and not x66 and not x68 and x21 and not x5 and x17 and x15 and x9 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( x65 and not x66 and not x68 and x21 and not x5 and x17 and x15 and not x9 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( x65 and not x66 and not x68 and x21 and not x5 and x17 and not x15 and x16 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x65 and not x66 and not x68 and x21 and not x5 and x17 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s212;

      elsif ( x65 and not x66 and not x68 and x21 and not x5 and not x17 ) = '1' then
         y15 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         y34 <= '1' ;
         current_group15m <= s294;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and x15 and x9 and x23 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and x15 and x9 and not x23 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and x15 and not x9 and x23 and x6 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and x15 and not x9 and x23 and not x6 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and x15 and not x9 and not x23 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and x16 and x9 and x8 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and x16 and x9 and not x8 and x10 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and x16 and x9 and not x8 and not x10 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and x16 and x9 and not x8 and not x10 and not x19 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and x16 and x9 and not x8 and not x10 and not x19 and x17 and not x14 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and x16 and x9 and not x8 and not x10 and not x19 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and x16 and x9 and not x8 and not x10 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and x16 and not x9 and x8 and x12 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and x16 and not x9 and x8 and not x12 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and x16 and not x9 and x8 and not x12 and not x19 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and x16 and not x9 and x8 and not x12 and not x19 and x17 and not x14 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and x16 and not x9 and x8 and not x12 and not x19 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and x16 and not x9 and x8 and not x12 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and x16 and not x9 and not x8 and x11 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and x16 and not x9 and not x8 and not x11 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and x16 and not x9 and not x8 and not x11 and not x19 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and x16 and not x9 and not x8 and not x11 and not x19 and x17 and not x14 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and x16 and not x9 and not x8 and not x11 and not x19 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and x16 and not x9 and not x8 and not x11 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and not x16 and x6 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s205;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and x23 and not x16 and not x6 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x66 and not x68 and not x21 and x22 and not x15 and not x23 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s205;

      elsif ( x65 and not x66 and not x68 and not x21 and not x22 and x23 and x20 and x14 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x66 and not x68 and not x21 and not x22 and x23 and x20 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x66 and not x68 and not x21 and not x22 and x23 and x20 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x68 and not x21 and not x22 and x23 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x68 and not x21 and not x22 and not x23 and x18 and x14 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x66 and not x68 and not x21 and not x22 and not x23 and x18 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x66 and not x68 and not x21 and not x22 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x68 and not x21 and not x22 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and x62 and x6 and x15 and x8 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s369;

      elsif ( not x65 and x66 and x67 and x62 and x6 and x15 and not x8 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s203;

      elsif ( not x65 and x66 and x67 and x62 and x6 and not x15 and x16 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s369;

      elsif ( not x65 and x66 and x67 and x62 and x6 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s135;

      elsif ( not x65 and x66 and x67 and x62 and not x6 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s369;

      elsif ( not x65 and x66 and x67 and not x62 and x63 and x17 and x13 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and x66 and x67 and not x62 and x63 and x17 and not x13 and x12 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and x66 and x67 and not x62 and x63 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x62 and x63 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and x16 and x4 and x14 and x8 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and x16 and x4 and x14 and not x8 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and x16 and x4 and not x14 and x7 and x8 ) = '1' then
         y24 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s157;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and x16 and x4 and not x14 and x7 and not x8 ) = '1' then
         y26 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s158;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and x16 and x4 and not x14 and not x7 and x8 and x12 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s65;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and x16 and x4 and not x14 and not x7 and x8 and not x12 and x19 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and x16 and x4 and not x14 and not x7 and x8 and not x12 and x19 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and x16 and x4 and not x14 and not x7 and x8 and not x12 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and x16 and x4 and not x14 and not x7 and not x8 and x13 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s65;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and x16 and x4 and not x14 and not x7 and not x8 and not x13 and x19 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and x16 and x4 and not x14 and not x7 and not x8 and not x13 and x19 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and x16 and x4 and not x14 and not x7 and not x8 and not x13 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and x16 and not x4 and x7 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s159;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and x16 and not x4 and not x7 and x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s190;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and x16 and not x4 and not x7 and not x3 and x8 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and x16 and not x4 and not x7 and not x3 and not x8 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s203;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and not x16 and x3 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s190;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and not x16 and not x3 and x4 and x7 and x11 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and not x16 and not x3 and x4 and x7 and not x11 and x8 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and not x16 and not x3 and x4 and x7 and not x11 and not x8 and x19 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and not x16 and not x3 and x4 and x7 and not x11 and not x8 and x19 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and not x16 and not x3 and x4 and x7 and not x11 and not x8 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and not x16 and not x3 and x4 and x7 and not x11 and not x8 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and not x16 and not x3 and x4 and not x7 and x8 and x9 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and not x16 and not x3 and x4 and not x7 and x8 and not x9 and x19 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and not x16 and not x3 and x4 and not x7 and x8 and not x9 and x19 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and not x16 and not x3 and x4 and not x7 and x8 and not x9 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and not x16 and not x3 and x4 and not x7 and x8 and not x9 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and not x16 and not x3 and x4 and not x7 and not x8 and x10 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and not x16 and not x3 and x4 and not x7 and not x8 and not x10 and x19 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and not x16 and not x3 and x4 and not x7 and not x8 and not x10 and x19 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and not x16 and not x3 and x4 and not x7 and not x8 and not x10 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and not x16 and not x3 and x4 and not x7 and not x8 and not x10 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and not x16 and not x3 and not x4 and x15 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and x64 and not x16 and not x3 and not x4 and not x15 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s204;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and not x64 and x15 and x8 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and not x64 and x15 and not x8 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and not x64 and not x15 and x16 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and not x64 and not x15 and not x16 and x14 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s135;

      elsif ( not x65 and x66 and x67 and not x62 and not x63 and not x64 and not x15 and not x16 and not x14 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s152;

      elsif ( not x65 and x66 and not x67 and x21 and x68 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x66 and not x67 and x21 and x68 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x66 and not x67 and x21 and x68 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and x21 and x68 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and x21 and not x68 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x65 and x66 and not x67 and x21 and not x68 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x65 and x66 and not x67 and x21 and not x68 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and x21 and not x68 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and x68 and x17 and x10 and x15 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s283;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and x68 and x17 and x10 and not x15 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and x68 and x17 and not x10 ) = '1' then
         y13 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s284;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and x68 and not x17 and x10 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s219;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and x68 and not x17 and not x10 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and not x68 and x23 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and not x68 and x23 and x17 and not x14 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and not x68 and x23 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and not x68 and x23 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and not x68 and not x23 and x10 and x12 and x18 and x14 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and not x68 and not x23 and x10 and x12 and x18 and not x14 and x13 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and not x68 and not x23 and x10 and x12 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and not x68 and not x23 and x10 and x12 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and not x68 and not x23 and x10 and not x12 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and not x68 and not x23 and not x10 and x18 and x14 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and not x68 and not x23 and not x10 and x18 and not x14 and x13 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and not x68 and not x23 and not x10 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and not x21 and x22 and not x68 and not x23 and not x10 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and not x21 and not x22 and x68 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x67 and not x21 and not x22 and not x68 and x23 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s180;

      elsif ( not x65 and x66 and not x67 and not x21 and not x22 and not x68 and not x23 and x15 and x9 ) = '1' then
         y4 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s370;

      elsif ( not x65 and x66 and not x67 and not x21 and not x22 and not x68 and not x23 and x15 and not x9 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and x66 and not x67 and not x21 and not x22 and not x68 and not x23 and not x15 and x16 and x7 and x9 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s330;

      elsif ( not x65 and x66 and not x67 and not x21 and not x22 and not x68 and not x23 and not x15 and x16 and x7 and not x9 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s333;

      elsif ( not x65 and x66 and not x67 and not x21 and not x22 and not x68 and not x23 and not x15 and x16 and not x7 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s330;

      elsif ( not x65 and x66 and not x67 and not x21 and not x22 and not x68 and not x23 and not x15 and not x16 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s285;

      elsif ( not x65 and not x66 and x21 and x68 ) = '1' then
         y1 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s142;

      elsif ( not x65 and not x66 and x21 and not x68 and x19 and x13 and x20 and x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and not x66 and x21 and not x68 and x19 and x13 and x20 and not x15 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and not x66 and x21 and not x68 and x19 and x13 and not x20 ) = '1' then
         y2 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s371;

      elsif ( not x65 and not x66 and x21 and not x68 and x19 and not x13 and x20 and x14 and x15 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x65 and not x66 and x21 and not x68 and x19 and not x13 and x20 and x14 and not x15 ) = '1' then
         y22 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s123;

      elsif ( not x65 and not x66 and x21 and not x68 and x19 and not x13 and x20 and not x14 and x15 and x4 ) = '1' then
         y2 <= '1' ;
         y11 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s372;

      elsif ( not x65 and not x66 and x21 and not x68 and x19 and not x13 and x20 and not x14 and x15 and not x4 and x9 and x3 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x66 and x21 and not x68 and x19 and not x13 and x20 and not x14 and x15 and not x4 and x9 and not x3 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x21 and not x68 and x19 and not x13 and x20 and not x14 and x15 and not x4 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x21 and not x68 and x19 and not x13 and x20 and not x14 and not x15 and x3 ) = '1' then
         y2 <= '1' ;
         y11 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s372;

      elsif ( not x65 and not x66 and x21 and not x68 and x19 and not x13 and x20 and not x14 and not x15 and not x3 and x9 and x4 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x66 and x21 and not x68 and x19 and not x13 and x20 and not x14 and not x15 and not x3 and x9 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x21 and not x68 and x19 and not x13 and x20 and not x14 and not x15 and not x3 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x21 and not x68 and x19 and not x13 and not x20 and x14 ) = '1' then
         y2 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s371;

      elsif ( not x65 and not x66 and x21 and not x68 and x19 and not x13 and not x20 and not x14 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s328;

      elsif ( not x65 and not x66 and x21 and not x68 and x19 and not x13 and not x20 and not x14 and not x5 and x6 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s107;

      elsif ( not x65 and not x66 and x21 and not x68 and x19 and not x13 and not x20 and not x14 and not x5 and not x6 and x15 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x66 and x21 and not x68 and x19 and not x13 and not x20 and not x14 and not x5 and not x6 and not x15 ) = '1' then
         y2 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      elsif ( not x65 and not x66 and x21 and not x68 and not x19 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s328;

      elsif ( not x65 and not x66 and x21 and not x68 and not x19 and not x5 and x20 and x14 and x18 ) = '1' then
         y2 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      elsif ( not x65 and not x66 and x21 and not x68 and not x19 and not x5 and x20 and x14 and not x18 and x15 ) = '1' then
         y2 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      elsif ( not x65 and not x66 and x21 and not x68 and not x19 and not x5 and x20 and x14 and not x18 and not x15 and x9 and x3 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x66 and x21 and not x68 and not x19 and not x5 and x20 and x14 and not x18 and not x15 and x9 and not x3 and x4 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x66 and x21 and not x68 and not x19 and not x5 and x20 and x14 and not x18 and not x15 and x9 and not x3 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x21 and not x68 and not x19 and not x5 and x20 and x14 and not x18 and not x15 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x21 and not x68 and not x19 and not x5 and x20 and not x14 and x15 and x16 ) = '1' then
         y2 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      elsif ( not x65 and not x66 and x21 and not x68 and not x19 and not x5 and x20 and not x14 and x15 and not x16 and x9 and x3 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x66 and x21 and not x68 and not x19 and not x5 and x20 and not x14 and x15 and not x16 and x9 and not x3 and x4 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x66 and x21 and not x68 and not x19 and not x5 and x20 and not x14 and x15 and not x16 and x9 and not x3 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x21 and not x68 and not x19 and not x5 and x20 and not x14 and x15 and not x16 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x21 and not x68 and not x19 and not x5 and x20 and not x14 and not x15 and x17 ) = '1' then
         y2 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      elsif ( not x65 and not x66 and x21 and not x68 and not x19 and not x5 and x20 and not x14 and not x15 and not x17 and x9 and x3 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x66 and x21 and not x68 and not x19 and not x5 and x20 and not x14 and not x15 and not x17 and x9 and not x3 and x4 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x66 and x21 and not x68 and not x19 and not x5 and x20 and not x14 and not x15 and not x17 and x9 and not x3 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x21 and not x68 and not x19 and not x5 and x20 and not x14 and not x15 and not x17 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x21 and not x68 and not x19 and not x5 and not x20 and x6 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s107;

      elsif ( not x65 and not x66 and x21 and not x68 and not x19 and not x5 and not x20 and not x6 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s373;

      elsif ( not x65 and not x66 and not x21 and x68 and x22 and x6 and x7 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x65 and not x66 and not x21 and x68 and x22 and x6 and not x7 and x8 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x65 and not x66 and not x21 and x68 and x22 and x6 and not x7 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x21 and x68 and x22 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x21 and x68 and not x22 and x15 ) = '1' then
         y1 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s142;

      elsif ( not x65 and not x66 and not x21 and x68 and not x22 and not x15 and x19 and x18 ) = '1' then
         y1 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s142;

      elsif ( not x65 and not x66 and not x21 and x68 and not x22 and not x15 and x19 and not x18 and x8 and x9 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x65 and not x66 and not x21 and x68 and not x22 and not x15 and x19 and not x18 and x8 and not x9 and x10 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x65 and not x66 and not x21 and x68 and not x22 and not x15 and x19 and not x18 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x21 and x68 and not x22 and not x15 and x19 and not x18 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x21 and x68 and not x22 and not x15 and not x19 ) = '1' then
         y1 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s142;

      elsif ( not x65 and not x66 and not x21 and not x68 and x22 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s108;

      elsif ( not x65 and not x66 and not x21 and not x68 and not x22 and x9 and x11 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x66 and not x21 and not x68 and not x22 and x9 and not x11 and x2 ) = '1' then
         current_group15m <= s101;

      elsif ( not x65 and not x66 and not x21 and not x68 and not x22 and x9 and not x11 and not x2 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( not x65 and not x66 and not x21 and not x68 and not x22 and not x9 and x8 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s108;

      else
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      end if;

   when s102 =>
      if ( x65 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and x16 and x12 and x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and x16 and x12 and not x19 and x18 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x65 and not x21 and x22 and x16 and x12 and not x19 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and x16 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and not x16 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and not x22 and x18 and x15 ) = '1' then
         y8 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s82;

      elsif ( not x65 and not x21 and not x22 and x18 and not x15 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s374;

      elsif ( not x65 and not x21 and not x22 and not x18 and x19 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s320;

      elsif ( not x65 and not x21 and not x22 and not x18 and x19 and not x15 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      else
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      end if;

   when s103 =>
      if ( x21 and x12 and x11 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( x21 and x12 and not x11 and x10 ) = '1' then
         current_group15m <= s103;

      elsif ( x21 and x12 and not x11 and not x10 ) = '1' then
         y10 <= '1' ;
         y17 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s104;

      elsif ( x21 and not x12 and x2 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( x21 and not x12 and not x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( not x21 and x22 and x19 and x15 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s177;

      elsif ( not x21 and x22 and x19 and not x15 ) = '1' then
         y2 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      elsif ( not x21 and x22 and not x19 and x20 and x14 and x18 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s178;

      elsif ( not x21 and x22 and not x19 and x20 and x14 and not x18 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and not x19 and x20 and x14 and not x18 and x5 and not x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and not x19 and x20 and x14 and not x18 and x5 and not x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x19 and x20 and x14 and not x18 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x19 and x20 and not x14 and x15 and x16 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s178;

      elsif ( not x21 and x22 and not x19 and x20 and not x14 and x15 and not x16 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and not x19 and x20 and not x14 and x15 and not x16 and x5 and not x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and not x19 and x20 and not x14 and x15 and not x16 and x5 and not x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x19 and x20 and not x14 and x15 and not x16 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x19 and x20 and not x14 and not x15 and x17 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s178;

      elsif ( not x21 and x22 and not x19 and x20 and not x14 and not x15 and not x17 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and not x19 and x20 and not x14 and not x15 and not x17 and x5 and not x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and not x19 and x20 and not x14 and not x15 and not x17 and x5 and not x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x19 and x20 and not x14 and not x15 and not x17 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x19 and not x20 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s151;

      elsif ( not x21 and not x22 and x7 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( not x21 and not x22 and not x7 and x10 and x19 and x15 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x21 and not x22 and not x7 and x10 and x19 and not x15 ) = '1' then
         y2 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      elsif ( not x21 and not x22 and not x7 and x10 and not x19 and x20 ) = '1' then
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s179;

      elsif ( not x21 and not x22 and not x7 and x10 and not x19 and not x20 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s151;

      else
         y10 <= '1' ;
         y17 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s104;

      end if;

   when s104 =>
      if ( x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x19 and x15 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s177;

      elsif ( not x21 and x22 and x19 and not x15 ) = '1' then
         y2 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      elsif ( not x21 and x22 and not x19 and x20 and x15 and x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s178;

      elsif ( not x21 and x22 and not x19 and x20 and x15 and not x14 and x16 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s178;

      elsif ( not x21 and x22 and not x19 and x20 and x15 and not x14 and not x16 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and not x19 and x20 and x15 and not x14 and not x16 and x5 and not x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and not x19 and x20 and x15 and not x14 and not x16 and x5 and not x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x19 and x20 and x15 and not x14 and not x16 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x19 and x20 and not x15 and x14 and x18 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s178;

      elsif ( not x21 and x22 and not x19 and x20 and not x15 and x14 and not x18 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and not x19 and x20 and not x15 and x14 and not x18 and x5 and not x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and not x19 and x20 and not x15 and x14 and not x18 and x5 and not x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x19 and x20 and not x15 and x14 and not x18 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x19 and x20 and not x15 and not x14 and x17 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s178;

      elsif ( not x21 and x22 and not x19 and x20 and not x15 and not x14 and not x17 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and not x19 and x20 and not x15 and not x14 and not x17 and x5 and not x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and not x19 and x20 and not x15 and not x14 and not x17 and x5 and not x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x19 and x20 and not x15 and not x14 and not x17 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x19 and not x20 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s151;

      else
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s176;

      end if;

   when s105 =>
      if ( x21 and x3 and x4 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( x21 and x3 and not x4 and x5 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( x21 and x3 and not x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x3 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 ) = '1' then
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s375;

      elsif ( not x21 and not x22 and x18 and x15 ) = '1' then
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s375;

      elsif ( not x21 and not x22 and x18 and not x15 and x4 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s273;

      elsif ( not x21 and not x22 and x18 and not x15 and not x4 ) = '1' then
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s375;

      elsif ( not x21 and not x22 and not x18 and x19 and x15 ) = '1' then
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s375;

      elsif ( not x21 and not x22 and not x18 and x19 and not x15 and x17 and x13 ) = '1' then
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s375;

      elsif ( not x21 and not x22 and not x18 and x19 and not x15 and x17 and not x13 and x16 ) = '1' then
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s375;

      elsif ( not x21 and not x22 and not x18 and x19 and not x15 and x17 and not x13 and not x16 and x8 and x9 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x21 and not x22 and not x18 and x19 and not x15 and x17 and not x13 and not x16 and x8 and not x9 and x10 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x21 and not x22 and not x18 and x19 and not x15 and x17 and not x13 and not x16 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x18 and x19 and not x15 and x17 and not x13 and not x16 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x18 and x19 and not x15 and not x17 and x16 and x14 ) = '1' then
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s375;

      elsif ( not x21 and not x22 and not x18 and x19 and not x15 and not x17 and x16 and not x14 and x8 and x9 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x21 and not x22 and not x18 and x19 and not x15 and not x17 and x16 and not x14 and x8 and not x9 and x10 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x21 and not x22 and not x18 and x19 and not x15 and not x17 and x16 and not x14 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x18 and x19 and not x15 and not x17 and x16 and not x14 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x18 and x19 and not x15 and not x17 and not x16 and x12 ) = '1' then
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s375;

      elsif ( not x21 and not x22 and not x18 and x19 and not x15 and not x17 and not x16 and not x12 and x8 and x9 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x21 and not x22 and not x18 and x19 and not x15 and not x17 and not x16 and not x12 and x8 and not x9 and x10 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x21 and not x22 and not x18 and x19 and not x15 and not x17 and not x16 and not x12 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x18 and x19 and not x15 and not x17 and not x16 and not x12 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x18 and not x19 and x4 ) = '1' then
         y14 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s376;

      else
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s375;

      end if;

   when s106 =>
      if ( x21 and x8 and x19 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( x21 and x8 and not x19 and x20 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s176;

      elsif ( x21 and x8 and not x19 and not x20 ) = '1' then
         y17 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s377;

      elsif ( x21 and not x8 ) = '1' then
         y8 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s378;

      elsif ( not x21 and x22 and x11 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s107;

      elsif ( not x21 and x22 and x11 and not x2 ) = '1' then
         current_group15m <= s40;

      elsif ( not x21 and x22 and not x11 and x9 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( not x21 and x22 and not x11 and not x9 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      else
         current_group15m <= s1;

      end if;

   when s107 =>
      if ( x21 and x19 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( x21 and not x19 ) = '1' then
         y17 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s377;

      elsif ( not x21 and x22 and x3 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s107;

      elsif ( not x21 and x22 and x3 and not x2 ) = '1' then
         current_group15m <= s40;

      elsif ( not x21 and x22 and not x3 ) = '1' then
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s179;

      else
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s379;

      end if;

   when s108 =>
      if ( x21 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s380;

      elsif ( not x21 and x22 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      else
         y1 <= '1' ;
         y2 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s107;

      end if;

   when s109 =>
      if ( x21 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s203;

      elsif ( not x21 and x22 and x6 and x7 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x21 and x22 and x6 and not x7 and x8 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x21 and x22 and x6 and not x7 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s110 =>
      if ( x66 and x21 and x5 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( x66 and x21 and not x5 and x19 and x15 and x10 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s330;

      elsif ( x66 and x21 and not x5 and x19 and x15 and not x10 and x12 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( x66 and x21 and not x5 and x19 and x15 and not x10 and not x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s48;

      elsif ( x66 and x21 and not x5 and x19 and not x15 and x16 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x66 and x21 and not x5 and x19 and not x15 and not x16 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s340;

      elsif ( x66 and x21 and not x5 and not x19 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s84;

      elsif ( x66 and not x21 and x22 and x23 and x3 and x15 and x10 ) = '1' then
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s339;

      elsif ( x66 and not x21 and x22 and x23 and x3 and x15 and not x10 and x12 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s126;

      elsif ( x66 and not x21 and x22 and x23 and x3 and x15 and not x10 and not x12 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      elsif ( x66 and not x21 and x22 and x23 and x3 and not x15 and x16 and x10 and x12 ) = '1' then
         y4 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s370;

      elsif ( x66 and not x21 and x22 and x23 and x3 and not x15 and x16 and x10 and not x12 ) = '1' then
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s381;

      elsif ( x66 and not x21 and x22 and x23 and x3 and not x15 and x16 and not x10 ) = '1' then
         y4 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s370;

      elsif ( x66 and not x21 and x22 and x23 and x3 and not x15 and not x16 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s180;

      elsif ( x66 and not x21 and x22 and x23 and not x3 ) = '1' then
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s339;

      elsif ( x66 and not x21 and x22 and not x23 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x66 and not x21 and not x22 and x15 and x4 and x7 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and not x21 and not x22 and x15 and x4 and not x7 and x23 and x9 ) = '1' then
         y4 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s370;

      elsif ( x66 and not x21 and not x22 and x15 and x4 and not x7 and x23 and not x9 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( x66 and not x21 and not x22 and x15 and x4 and not x7 and not x23 and x9 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s341;

      elsif ( x66 and not x21 and not x22 and x15 and x4 and not x7 and not x23 and not x9 ) = '1' then
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s339;

      elsif ( x66 and not x21 and not x22 and x15 and not x4 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x66 and not x21 and not x22 and not x15 and x16 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x66 and not x21 and not x22 and not x15 and not x16 and x23 and x4 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s285;

      elsif ( x66 and not x21 and not x22 and not x15 and not x16 and x23 and not x4 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s48;

      elsif ( x66 and not x21 and not x22 and not x15 and not x16 and not x23 and x4 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s336;

      elsif ( x66 and not x21 and not x22 and not x15 and not x16 and not x23 and not x4 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      elsif ( not x66 and x67 and x24 and x26 and x20 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x66 and x67 and x24 and x26 and not x20 and x21 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x66 and x67 and x24 and x26 and not x20 and not x21 and x22 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x66 and x67 and x24 and x26 and not x20 and not x21 and not x22 and x23 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x66 and x67 and x24 and x26 and not x20 and not x21 and not x22 and not x23 and x16 and x11 ) = '1' then
         y12 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s49;

      elsif ( not x66 and x67 and x24 and x26 and not x20 and not x21 and not x22 and not x23 and x16 and not x11 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x66 and x67 and x24 and x26 and not x20 and not x21 and not x22 and not x23 and not x16 and x17 and x13 and x11 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x66 and x67 and x24 and x26 and not x20 and not x21 and not x22 and not x23 and not x16 and x17 and x13 and not x11 and x12 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( not x66 and x67 and x24 and x26 and not x20 and not x21 and not x22 and not x23 and not x16 and x17 and x13 and not x11 and not x12 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x66 and x67 and x24 and x26 and not x20 and not x21 and not x22 and not x23 and not x16 and x17 and not x13 and x11 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x66 and x67 and x24 and x26 and not x20 and not x21 and not x22 and not x23 and not x16 and x17 and not x13 and not x11 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x66 and x67 and x24 and x26 and not x20 and not x21 and not x22 and not x23 and not x16 and not x17 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s51;

      elsif ( not x66 and x67 and x24 and not x26 and x16 and x11 and x12 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s188;

      elsif ( not x66 and x67 and x24 and not x26 and x16 and x11 and not x12 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s172;

      elsif ( not x66 and x67 and x24 and not x26 and x16 and not x11 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s160;

      elsif ( not x66 and x67 and x24 and not x26 and not x16 and x17 and x11 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x66 and x67 and x24 and not x26 and not x16 and x17 and x11 and not x13 ) = '1' then
         y15 <= '1' ;
         y112 <= '1' ;
         current_group15m <= s46;

      elsif ( not x66 and x67 and x24 and not x26 and not x16 and x17 and not x11 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x66 and x67 and x24 and not x26 and not x16 and not x17 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and x67 and not x24 and x25 and x26 and x4 and x15 and x10 and x11 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x66 and x67 and not x24 and x25 and x26 and x4 and x15 and x10 and not x11 and x12 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s65;

      elsif ( not x66 and x67 and not x24 and x25 and x26 and x4 and x15 and x10 and not x11 and not x12 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s161;

      elsif ( not x66 and x67 and not x24 and x25 and x26 and x4 and x15 and not x10 and x12 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s186;

      elsif ( not x66 and x67 and not x24 and x25 and x26 and x4 and x15 and not x10 and not x12 ) = '1' then
         y12 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s49;

      elsif ( not x66 and x67 and not x24 and x25 and x26 and x4 and not x15 and x16 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x66 and x67 and not x24 and x25 and x26 and x4 and not x15 and not x16 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and x67 and not x24 and x25 and x26 and not x4 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x66 and x67 and not x24 and x25 and not x26 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x66 and x67 and not x24 and x25 and not x26 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x66 and x67 and not x24 and x25 and not x26 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and x25 and not x26 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and x17 and x10 and x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and x17 and x10 and not x12 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s160;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and x17 and not x10 and x11 and x12 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s171;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and x17 and not x10 and x11 and not x12 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s160;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and x17 and not x10 and not x11 and x12 and x13 ) = '1' then
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s239;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and x17 and not x10 and not x11 and x12 and not x13 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and x17 and not x10 and not x11 and x12 and not x13 and x18 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and x17 and not x10 and not x11 and x12 and not x13 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and x17 and not x10 and not x11 and not x12 and x14 ) = '1' then
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s239;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and x17 and not x10 and not x11 and not x12 and not x14 and x18 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and x17 and not x10 and not x11 and not x12 and not x14 and x18 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and x17 and not x10 and not x11 and not x12 and not x14 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and not x17 and x12 and x10 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and not x17 and x12 and x10 and not x2 and x4 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and not x17 and x12 and x10 and not x2 and not x4 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s382;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and not x17 and x12 and not x10 and x11 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and not x17 and x12 and not x10 and not x11 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and not x17 and x12 and not x10 and not x11 and not x2 and x4 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and not x17 and x12 and not x10 and not x11 and not x2 and not x4 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s382;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and not x17 and not x12 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and not x17 and not x12 and not x2 and x11 and x4 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and not x17 and not x12 and not x2 and x11 and not x4 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s382;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and not x17 and not x12 and not x2 and not x11 and x10 and x4 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and not x17 and not x12 and not x2 and not x11 and x10 and not x4 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s48;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and not x17 and not x12 and not x2 and not x11 and not x10 and x4 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and x26 and not x17 and not x12 and not x2 and not x11 and not x10 and not x4 ) = '1' then
         y8 <= '1' ;
         y17 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s164;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and x15 and x10 and x12 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and x15 and x10 and not x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and x15 and not x10 and x11 and x12 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s160;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and x15 and not x10 and x11 and not x12 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s171;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and x15 and not x10 and not x11 and x12 and x13 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s181;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and x15 and not x10 and not x11 and x12 and not x13 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and x15 and not x10 and not x11 and x12 and not x13 and x17 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and x15 and not x10 and not x11 and x12 and not x13 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and x15 and not x10 and not x11 and not x12 and x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s181;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and x15 and not x10 and not x11 and not x12 and not x14 and x17 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and x15 and not x10 and not x11 and not x12 and not x14 and x17 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and x15 and not x10 and not x11 and not x12 and not x14 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and x12 and x10 and x8 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and x12 and x10 and x8 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and x12 and x10 and x8 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and x12 and x10 and x8 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and x12 and x10 and not x8 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and x12 and x10 and not x8 and not x3 and x5 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and x12 and x10 and not x8 and not x3 and not x5 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and x12 and not x10 and x7 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and x12 and not x10 and x7 and not x3 and x5 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and x12 and not x10 and x7 and not x3 and not x5 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and x12 and not x10 and not x7 and x11 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and x12 and not x10 and not x7 and x11 and not x3 and x5 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and x12 and not x10 and not x7 and x11 and not x3 and not x5 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and x12 and not x10 and not x7 and not x11 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and x12 and not x10 and not x7 and not x11 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and x12 and not x10 and not x7 and not x11 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and x12 and not x10 and not x7 and not x11 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and not x12 and x10 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and not x12 and x10 and not x3 and x5 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s172;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and not x12 and x10 and not x3 and not x5 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and not x12 and not x10 and x11 and x9 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and not x12 and not x10 and x11 and x9 and not x3 and x5 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and not x12 and not x10 and x11 and x9 and not x3 and not x5 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and not x12 and not x10 and x11 and not x9 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and not x12 and not x10 and x11 and not x9 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and not x12 and not x10 and x11 and not x9 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and not x12 and not x10 and x11 and not x9 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and not x12 and not x10 and not x11 and x8 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and not x12 and not x10 and not x11 and x8 and not x3 and x5 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and not x12 and not x10 and not x11 and x8 and not x3 and not x5 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and not x12 and not x10 and not x11 and not x8 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and not x12 and not x10 and not x11 and not x8 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and not x12 and not x10 and not x11 and not x8 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and x16 and not x26 and not x15 and not x12 and not x10 and not x11 and not x8 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and x12 and x10 and x8 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and x12 and x10 and x8 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and x12 and x10 and x8 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and x12 and x10 and x8 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and x12 and x10 and not x8 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and x12 and x10 and not x8 and not x2 and x4 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and x12 and x10 and not x8 and not x2 and not x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and x12 and not x10 and x7 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and x12 and not x10 and x7 and not x2 and x4 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and x12 and not x10 and x7 and not x2 and not x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and x12 and not x10 and not x7 and x11 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and x12 and not x10 and not x7 and x11 and not x2 and x4 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and x12 and not x10 and not x7 and x11 and not x2 and not x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and x12 and not x10 and not x7 and not x11 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and x12 and not x10 and not x7 and not x11 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and x12 and not x10 and not x7 and not x11 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and x12 and not x10 and not x7 and not x11 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and not x12 and x10 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and not x12 and x10 and not x2 and x4 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s297;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and not x12 and x10 and not x2 and not x4 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and not x12 and not x10 and x11 and x9 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and not x12 and not x10 and x11 and x9 and not x2 and x4 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and not x12 and not x10 and x11 and x9 and not x2 and not x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and not x12 and not x10 and x11 and not x9 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and not x12 and not x10 and x11 and not x9 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and not x12 and not x10 and x11 and not x9 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and not x12 and not x10 and x11 and not x9 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and not x12 and not x10 and not x11 and x8 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and not x12 and not x10 and not x11 and x8 and not x2 and x4 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and not x12 and not x10 and not x11 and x8 and not x2 and not x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and not x12 and not x10 and not x11 and not x8 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and not x12 and not x10 and not x11 and not x8 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and not x12 and not x10 and not x11 and not x8 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and x17 and not x12 and not x10 and not x11 and not x8 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and not x17 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and not x17 and not x2 and x4 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and x26 and not x17 and not x2 and not x4 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s382;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and not x26 and x12 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and not x26 and x12 and not x3 and x5 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and not x26 and x12 and not x3 and not x5 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and not x26 and not x12 and x15 and x11 and x10 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and not x26 and not x12 and x15 and x11 and x10 and not x3 and x5 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and not x26 and not x12 and x15 and x11 and x10 and not x3 and not x5 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and not x26 and not x12 and x15 and x11 and not x10 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and not x26 and not x12 and x15 and not x11 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and not x26 and not x12 and x15 and not x11 and not x3 and x5 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and not x26 and not x12 and x15 and not x11 and not x3 and not x5 and x10 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s160;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and not x26 and not x12 and x15 and not x11 and not x3 and not x5 and not x10 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s48;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and not x26 and not x12 and not x15 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s242;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and not x26 and not x12 and not x15 and not x3 and x5 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and x67 and not x24 and not x25 and not x16 and not x26 and not x12 and not x15 and not x3 and not x5 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x66 and not x67 and x21 and x68 and x12 and x7 and x19 and x17 ) = '1' then
         y14 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s383;

      elsif ( not x66 and not x67 and x21 and x68 and x12 and x7 and x19 and not x17 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s385;

      elsif ( not x66 and not x67 and x21 and x68 and x12 and x7 and not x19 and x20 ) = '1' then
         y14 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s383;

      elsif ( not x66 and not x67 and x21 and x68 and x12 and x7 and not x19 and not x20 ) = '1' then
         y14 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s384;

      elsif ( not x66 and not x67 and x21 and x68 and x12 and not x7 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s385;

      elsif ( not x66 and not x67 and x21 and x68 and not x12 and x19 and x7 and x17 ) = '1' then
         y14 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s383;

      elsif ( not x66 and not x67 and x21 and x68 and not x12 and x19 and x7 and not x17 ) = '1' then
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s273;

      elsif ( not x66 and not x67 and x21 and x68 and not x12 and x19 and not x7 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s385;

      elsif ( not x66 and not x67 and x21 and x68 and not x12 and not x19 and x20 and x17 and x14 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s385;

      elsif ( not x66 and not x67 and x21 and x68 and not x12 and not x19 and x20 and x17 and not x14 and x16 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s385;

      elsif ( not x66 and not x67 and x21 and x68 and not x12 and not x19 and x20 and x17 and not x14 and not x16 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x67 and x21 and x68 and not x12 and not x19 and x20 and not x17 and x16 and x15 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s385;

      elsif ( not x66 and not x67 and x21 and x68 and not x12 and not x19 and x20 and not x17 and x16 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x67 and x21 and x68 and not x12 and not x19 and x20 and not x17 and not x16 and x13 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s385;

      elsif ( not x66 and not x67 and x21 and x68 and not x12 and not x19 and x20 and not x17 and not x16 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x67 and x21 and x68 and not x12 and not x19 and not x20 and x7 ) = '1' then
         y14 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s376;

      elsif ( not x66 and not x67 and x21 and x68 and not x12 and not x19 and not x20 and not x7 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s385;

      elsif ( not x66 and not x67 and x21 and not x68 and x19 and x7 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s177;

      elsif ( not x66 and not x67 and x21 and not x68 and x19 and not x7 ) = '1' then
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s179;

      elsif ( not x66 and not x67 and x21 and not x68 and not x19 and x20 and x15 and x14 ) = '1' then
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s179;

      elsif ( not x66 and not x67 and x21 and not x68 and not x19 and x20 and x15 and not x14 and x16 ) = '1' then
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s179;

      elsif ( not x66 and not x67 and x21 and not x68 and not x19 and x20 and x15 and not x14 and not x16 and x9 and x3 ) = '1' then
         current_group15m <= s40;

      elsif ( not x66 and not x67 and x21 and not x68 and not x19 and x20 and x15 and not x14 and not x16 and x9 and not x3 and x4 ) = '1' then
         current_group15m <= s40;

      elsif ( not x66 and not x67 and x21 and not x68 and not x19 and x20 and x15 and not x14 and not x16 and x9 and not x3 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x67 and x21 and not x68 and not x19 and x20 and x15 and not x14 and not x16 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x67 and x21 and not x68 and not x19 and x20 and not x15 and x14 and x18 ) = '1' then
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s179;

      elsif ( not x66 and not x67 and x21 and not x68 and not x19 and x20 and not x15 and x14 and not x18 and x9 and x3 ) = '1' then
         current_group15m <= s40;

      elsif ( not x66 and not x67 and x21 and not x68 and not x19 and x20 and not x15 and x14 and not x18 and x9 and not x3 and x4 ) = '1' then
         current_group15m <= s40;

      elsif ( not x66 and not x67 and x21 and not x68 and not x19 and x20 and not x15 and x14 and not x18 and x9 and not x3 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x67 and x21 and not x68 and not x19 and x20 and not x15 and x14 and not x18 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x67 and x21 and not x68 and not x19 and x20 and not x15 and not x14 and x17 ) = '1' then
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s179;

      elsif ( not x66 and not x67 and x21 and not x68 and not x19 and x20 and not x15 and not x14 and not x17 and x9 and x3 ) = '1' then
         current_group15m <= s40;

      elsif ( not x66 and not x67 and x21 and not x68 and not x19 and x20 and not x15 and not x14 and not x17 and x9 and not x3 and x4 ) = '1' then
         current_group15m <= s40;

      elsif ( not x66 and not x67 and x21 and not x68 and not x19 and x20 and not x15 and not x14 and not x17 and x9 and not x3 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x67 and x21 and not x68 and not x19 and x20 and not x15 and not x14 and not x17 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x67 and x21 and not x68 and not x19 and not x20 and x7 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s151;

      elsif ( not x66 and not x67 and x21 and not x68 and not x19 and not x20 and not x7 ) = '1' then
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s179;

      elsif ( not x66 and not x67 and not x21 and x22 and x68 and x12 and x18 and x17 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s271;

      elsif ( not x66 and not x67 and not x21 and x22 and x68 and x12 and x18 and not x17 ) = '1' then
         y6 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s386;

      elsif ( not x66 and not x67 and not x21 and x22 and x68 and x12 and not x18 and x19 and x17 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s271;

      elsif ( not x66 and not x67 and not x21 and x22 and x68 and x12 and not x18 and x19 and not x17 and x3 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s387;

      elsif ( not x66 and not x67 and not x21 and x22 and x68 and x12 and not x18 and x19 and not x17 and not x3 ) = '1' then
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s388;

      elsif ( not x66 and not x67 and not x21 and x22 and x68 and x12 and not x18 and not x19 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s271;

      elsif ( not x66 and not x67 and not x21 and x22 and x68 and not x12 and x18 and x17 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s271;

      elsif ( not x66 and not x67 and not x21 and x22 and x68 and not x12 and x18 and not x17 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s374;

      elsif ( not x66 and not x67 and not x21 and x22 and x68 and not x12 and not x18 and x19 ) = '1' then
         y4 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s273;

      elsif ( not x66 and not x67 and not x21 and x22 and x68 and not x12 and not x18 and not x19 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x66 and not x67 and not x21 and x22 and not x68 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x67 and not x21 and not x22 and x68 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and x19 and x13 and x20 and x15 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and x19 and x13 and x20 and not x15 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and x19 and x13 and not x20 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and x19 and not x13 and x14 and x20 and x15 ) = '1' then
         y22 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s123;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and x19 and not x13 and x14 and x20 and not x15 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s373;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and x19 and not x13 and x14 and not x20 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and x19 and not x13 and not x14 and x20 and x15 and x6 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s181;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and x19 and not x13 and not x14 and x20 and x15 and not x6 and x4 and x5 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and x19 and not x13 and not x14 and x20 and x15 and not x6 and x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and x19 and not x13 and not x14 and x20 and x15 and not x6 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and x19 and not x13 and not x14 and x20 and not x15 and x5 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s181;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and x19 and not x13 and not x14 and x20 and not x15 and not x5 and x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and x19 and not x13 and not x14 and x20 and not x15 and not x5 and x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and x19 and not x13 and not x14 and x20 and not x15 and not x5 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and x19 and not x13 and not x14 and not x20 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s328;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and x19 and not x13 and not x14 and not x20 and not x3 and x7 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s177;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and x19 and not x13 and not x14 and not x20 and not x3 and not x7 and x15 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s126;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and x19 and not x13 and not x14 and not x20 and not x3 and not x7 and not x15 ) = '1' then
         y2 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s371;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and not x19 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s328;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and not x19 and not x3 and x20 and x14 and x18 ) = '1' then
         y2 <= '1' ;
         y11 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s123;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and not x19 and not x3 and x20 and x14 and not x18 and x15 ) = '1' then
         y2 <= '1' ;
         y11 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s123;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and not x19 and not x3 and x20 and x14 and not x18 and not x15 and x4 and x5 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and not x19 and not x3 and x20 and x14 and not x18 and not x15 and x4 and not x5 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and not x19 and not x3 and x20 and x14 and not x18 and not x15 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and not x19 and not x3 and x20 and x14 and not x18 and not x15 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and not x19 and not x3 and x20 and not x14 and x15 and x16 ) = '1' then
         y2 <= '1' ;
         y11 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s123;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and not x19 and not x3 and x20 and not x14 and x15 and not x16 and x4 and x5 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and not x19 and not x3 and x20 and not x14 and x15 and not x16 and x4 and not x5 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and not x19 and not x3 and x20 and not x14 and x15 and not x16 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and not x19 and not x3 and x20 and not x14 and x15 and not x16 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and not x19 and not x3 and x20 and not x14 and not x15 and x17 ) = '1' then
         y2 <= '1' ;
         y11 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s123;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and not x19 and not x3 and x20 and not x14 and not x15 and not x17 and x4 and x5 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and not x19 and not x3 and x20 and not x14 and not x15 and not x17 and x4 and not x5 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and not x19 and not x3 and x20 and not x14 and not x15 and not x17 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and not x19 and not x3 and x20 and not x14 and not x15 and not x17 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x67 and not x21 and not x22 and not x68 and not x19 and not x3 and not x20 and x7 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s177;

      else
         y17 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s377;

      end if;

   when s111 =>
      if ( x22 and x17 and x18 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x22 and x17 and not x18 and x19 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x22 and x17 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x22 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x22 and x18 and x13 and x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( not x22 and x18 and x13 and not x23 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( not x22 and x18 and not x13 and x12 and x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( not x22 and x18 and not x13 and x12 and not x23 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( not x22 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s112 =>
      if ( x65 and x66 and x22 ) = '1' then
         y9 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s111;

      elsif ( x65 and x66 and not x22 and x23 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and x66 and not x22 and not x23 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x65 and not x66 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x21 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x65 and x66 and x21 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x65 and x66 and x21 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x21 and x22 and x23 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s286;

      elsif ( not x65 and x66 and not x21 and x22 and not x23 and x18 and x14 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and x66 and not x21 and x22 and not x23 and x18 and not x14 and x13 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and x66 and not x21 and x22 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x21 and x22 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x21 and not x22 and x23 and x19 and x14 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x65 and x66 and not x21 and not x22 and x23 and x19 and not x14 and x13 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x65 and x66 and not x21 and not x22 and x23 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x21 and not x22 and x23 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x21 and not x22 and not x23 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and not x66 and x20 and x15 and x16 and x8 and x14 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x65 and not x66 and x20 and x15 and x16 and x8 and not x14 and x7 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s126;

      elsif ( not x65 and not x66 and x20 and x15 and x16 and x8 and not x14 and not x7 and x12 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s191;

      elsif ( not x65 and not x66 and x20 and x15 and x16 and x8 and not x14 and not x7 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x20 and x15 and x16 and not x8 and x14 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x65 and not x66 and x20 and x15 and x16 and not x8 and not x14 and x7 ) = '1' then
         y1 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y13 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s207;

      elsif ( not x65 and not x66 and x20 and x15 and x16 and not x8 and not x14 and not x7 and x13 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s191;

      elsif ( not x65 and not x66 and x20 and x15 and x16 and not x8 and not x14 and not x7 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x20 and x15 and not x16 and x7 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s191;

      elsif ( not x65 and not x66 and x20 and x15 and not x16 and not x7 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s44;

      elsif ( not x65 and not x66 and x20 and x15 and not x16 and not x7 and not x5 and x8 and x1 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s254;

      elsif ( not x65 and not x66 and x20 and x15 and not x16 and not x7 and not x5 and x8 and not x1 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( not x65 and not x66 and x20 and x15 and not x16 and not x7 and not x5 and not x8 and x1 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x65 and not x66 and x20 and x15 and not x16 and not x7 and not x5 and not x8 and not x1 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x65 and not x66 and x20 and not x15 and x16 and x7 and x8 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s44;

      elsif ( not x65 and not x66 and x20 and not x15 and x16 and x7 and x8 and not x5 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x65 and not x66 and x20 and not x15 and x16 and x7 and not x8 and x11 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s44;

      elsif ( not x65 and not x66 and x20 and not x15 and x16 and x7 and not x8 and x11 and not x5 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x65 and not x66 and x20 and not x15 and x16 and x7 and not x8 and not x11 and x18 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x66 and x20 and not x15 and x16 and x7 and not x8 and not x11 and x18 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x66 and x20 and not x15 and x16 and x7 and not x8 and not x11 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x20 and not x15 and x16 and x7 and not x8 and not x11 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x20 and not x15 and x16 and not x7 and x8 and x9 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s44;

      elsif ( not x65 and not x66 and x20 and not x15 and x16 and not x7 and x8 and x9 and not x5 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x65 and not x66 and x20 and not x15 and x16 and not x7 and x8 and not x9 and x18 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x66 and x20 and not x15 and x16 and not x7 and x8 and not x9 and x18 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x66 and x20 and not x15 and x16 and not x7 and x8 and not x9 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x20 and not x15 and x16 and not x7 and x8 and not x9 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x20 and not x15 and x16 and not x7 and not x8 and x10 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s44;

      elsif ( not x65 and not x66 and x20 and not x15 and x16 and not x7 and not x8 and x10 and not x5 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x65 and not x66 and x20 and not x15 and x16 and not x7 and not x8 and not x10 and x18 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x66 and x20 and not x15 and x16 and not x7 and not x8 and not x10 and x18 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x66 and x20 and not x15 and x16 and not x7 and not x8 and not x10 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x20 and not x15 and x16 and not x7 and not x8 and not x10 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x20 and not x15 and not x16 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s44;

      elsif ( not x65 and not x66 and x20 and not x15 and not x16 and not x5 and x1 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x65 and not x66 and x20 and not x15 and not x16 and not x5 and not x1 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s210;

      else
         current_group15m <= s1;

      end if;

   when s113 =>
      if ( x21 and x19 and x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x21 and x19 and not x15 and x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x21 and x19 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x20 and x15 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( not x21 and x20 and not x15 and x14 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( not x21 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s114 =>
      if ( x67 and x65 and x21 and x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x67 and x65 and x21 and x8 and not x9 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x67 and x65 and x21 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x65 and x21 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x65 and not x21 and x23 and x22 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x67 and x65 and not x21 and x23 and x22 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x67 and x65 and not x21 and x23 and x22 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x65 and not x21 and x23 and x22 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x65 and not x21 and x23 and not x22 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x67 and x65 and not x21 and x23 and not x22 and x9 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x67 and x65 and not x21 and x23 and not x22 and x9 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x65 and not x21 and x23 and not x22 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x65 and not x21 and not x23 and x8 and x22 and x9 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x67 and x65 and not x21 and not x23 and x8 and x22 and not x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x67 and x65 and not x21 and not x23 and x8 and x22 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x65 and not x21 and not x23 and x8 and not x22 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x67 and x65 and not x21 and not x23 and x8 and not x22 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x67 and x65 and not x21 and not x23 and x8 and not x22 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x65 and not x21 and not x23 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x65 and x66 and x68 and x21 and x19 and x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x67 and not x65 and x66 and x68 and x21 and x19 and not x15 and x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x67 and not x65 and x66 and x68 and x21 and x19 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x65 and x66 and x68 and x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x65 and x66 and x68 and not x21 and x20 and x15 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x67 and not x65 and x66 and x68 and not x21 and x20 and not x15 and x14 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x67 and not x65 and x66 and x68 and not x21 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x65 and x66 and x68 and not x21 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x65 and x66 and not x68 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x65 and not x66 and x24 and x26 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s183;

      elsif ( x67 and not x65 and not x66 and x24 and not x26 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( x67 and not x65 and not x66 and x24 and not x26 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( x67 and not x65 and not x66 and x24 and not x26 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x65 and not x66 and x24 and not x26 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x65 and not x66 and not x24 and x25 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( x67 and not x65 and not x66 and not x24 and x25 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( x67 and not x65 and not x66 and not x24 and x25 and x19 and not x14 and not x13 and x26 ) = '1' then
         current_group15m <= s114;

      elsif ( x67 and not x65 and not x66 and not x24 and x25 and x19 and not x14 and not x13 and not x26 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x65 and not x66 and not x24 and x25 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x65 and not x66 and not x24 and not x25 and x26 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( x67 and not x65 and not x66 and not x24 and not x25 and x26 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( x67 and not x65 and not x66 and not x24 and not x25 and x26 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x65 and not x66 and not x24 and not x25 and x26 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x65 and not x66 and not x24 and not x25 and not x26 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( x67 and not x65 and not x66 and not x24 and not x25 and not x26 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( x67 and not x65 and not x66 and not x24 and not x25 and not x26 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x65 and not x66 and not x24 and not x25 and not x26 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x65 and x21 and x18 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x67 and x65 and x21 and not x18 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x67 and x65 and x21 and not x18 and x19 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x67 and x65 and x21 and not x18 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x65 and x21 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x65 and not x21 and x23 and x22 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( not x67 and x65 and not x21 and x23 and x22 and not x19 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( not x67 and x65 and not x21 and x23 and x22 and not x19 and x17 and not x14 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( not x67 and x65 and not x21 and x23 and x22 and not x19 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x65 and not x21 and x23 and x22 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x65 and not x21 and x23 and not x22 and x20 and x14 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( not x67 and x65 and not x21 and x23 and not x22 and x20 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( not x67 and x65 and not x21 and x23 and not x22 and x20 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x65 and not x21 and x23 and not x22 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x65 and not x21 and not x23 and x18 and x14 and x22 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( not x67 and x65 and not x21 and not x23 and x18 and x14 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x67 and x65 and not x21 and not x23 and x18 and not x14 and x13 and x22 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( not x67 and x65 and not x21 and not x23 and x18 and not x14 and x13 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x67 and x65 and not x21 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x65 and not x21 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x65 and x21 and x66 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x67 and not x65 and x21 and x66 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x67 and not x65 and x21 and x66 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x65 and x21 and x66 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x65 and x21 and not x66 and x3 and x4 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( not x67 and not x65 and x21 and not x66 and x3 and not x4 and x5 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( not x67 and not x65 and x21 and not x66 and x3 and not x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x65 and x21 and not x66 and not x3 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x65 and not x21 and x22 and x66 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x67 and not x65 and not x21 and x22 and not x66 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x67 and not x65 and not x21 and not x22 and x66 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x67 and not x65 and not x21 and not x22 and x66 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x67 and not x65 and not x21 and not x22 and x66 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x65 and not x21 and not x22 and x66 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x65 and not x21 and not x22 and not x66 and x8 and x9 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x67 and not x65 and not x21 and not x22 and not x66 and x8 and not x9 and x10 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x67 and not x65 and not x21 and not x22 and not x66 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s115 =>
      if ( x21 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s344;

      end if;

   when s116 =>
      if ( x21 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( not x21 and x22 and x8 and x9 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x8 and not x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x12 and x23 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s247;

      elsif ( not x21 and not x22 and x12 and not x23 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x21 and not x22 and not x12 and x23 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and not x12 and x23 and x9 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and not x12 and x23 and x9 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x12 and x23 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x12 and not x23 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and not x12 and not x23 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and not x12 and not x23 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s117 =>
      if ( x21 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( not x21 and x22 and x23 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x21 and x22 and x23 and not x12 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x23 and not x12 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x23 and not x12 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and not x12 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 and x18 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and not x23 and not x18 and x8 and x9 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and not x23 and not x18 and x8 and not x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and not x23 and not x18 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 and not x18 and not x8 ) = '1' then
         current_group15m <= s1;

      else
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s243;

      end if;

   when s118 =>
      if ( x60 and x61 and x18 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s38;

      elsif ( x60 and x61 and not x18 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( x60 and not x61 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s356;

      elsif ( not x60 and x61 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s356;

      elsif ( not x60 and not x61 and x62 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s154;

      else
         y7 <= '1' ;
         current_group15m <= s338;

      end if;

   when s119 =>
      if ( x21 and x15 and x16 and x9 and x7 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and x15 and x16 and x9 and not x7 and x8 ) = '1' then
         y24 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s157;

      elsif ( x21 and x15 and x16 and x9 and not x7 and not x8 and x13 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s191;

      elsif ( x21 and x15 and x16 and x9 and not x7 and not x8 and not x13 and x18 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x21 and x15 and x16 and x9 and not x7 and not x8 and not x13 and not x18 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x21 and x15 and x16 and x9 and not x7 and not x8 and not x13 and not x18 and x19 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x15 and x16 and x9 and not x7 and not x8 and not x13 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x15 and x16 and not x9 and x7 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x21 and x15 and x16 and not x9 and not x7 and x8 ) = '1' then
         y26 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s158;

      elsif ( x21 and x15 and x16 and not x9 and not x7 and not x8 and x14 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s191;

      elsif ( x21 and x15 and x16 and not x9 and not x7 and not x8 and not x14 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( x21 and x15 and not x16 and x7 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s147;

      elsif ( x21 and x15 and not x16 and not x7 and x8 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s147;

      elsif ( x21 and x15 and not x16 and not x7 and not x8 and x2 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s22;

      elsif ( x21 and x15 and not x16 and not x7 and not x8 and not x2 and x5 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x21 and x15 and not x16 and not x7 and not x8 and not x2 and not x5 and x9 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x21 and x15 and not x16 and not x7 and not x8 and not x2 and not x5 and not x9 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( x21 and not x15 and x2 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s22;

      elsif ( x21 and not x15 and not x2 and x16 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and not x15 and not x2 and x16 and x9 and not x10 and x8 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and not x15 and not x2 and x16 and x9 and not x10 and not x8 and x18 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x21 and not x15 and not x2 and x16 and x9 and not x10 and not x8 and not x18 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x21 and not x15 and not x2 and x16 and x9 and not x10 and not x8 and not x18 and x19 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x21 and not x15 and not x2 and x16 and x9 and not x10 and not x8 and not x18 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x15 and not x2 and x16 and x9 and not x10 and not x8 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x15 and not x2 and x16 and not x9 and x8 and x12 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and not x15 and not x2 and x16 and not x9 and x8 and not x12 and x18 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x21 and not x15 and not x2 and x16 and not x9 and x8 and not x12 and not x18 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x21 and not x15 and not x2 and x16 and not x9 and x8 and not x12 and not x18 and x19 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x21 and not x15 and not x2 and x16 and not x9 and x8 and not x12 and not x18 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x15 and not x2 and x16 and not x9 and x8 and not x12 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x15 and not x2 and x16 and not x9 and not x8 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and not x15 and not x2 and x16 and not x9 and not x8 and not x11 and x18 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x21 and not x15 and not x2 and x16 and not x9 and not x8 and not x11 and not x18 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x21 and not x15 and not x2 and x16 and not x9 and not x8 and not x11 and not x18 and x19 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x21 and not x15 and not x2 and x16 and not x9 and not x8 and not x11 and not x18 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x15 and not x2 and x16 and not x9 and not x8 and not x11 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x15 and not x2 and not x16 and x5 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x21 and not x15 and not x2 and not x16 and not x5 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s205;

      elsif ( not x21 and x22 and x18 and x14 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( not x21 and x22 and x18 and not x14 and x13 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( not x21 and x22 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x18 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s120 =>
      if ( x21 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s363;

      elsif ( not x21 and x23 and x22 and x5 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x21 and x23 and x22 and not x5 and x18 and x15 and x9 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x21 and x23 and x22 and not x5 and x18 and x15 and not x9 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x21 and x23 and x22 and not x5 and x18 and not x15 and x16 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x21 and x23 and x22 and not x5 and x18 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s205;

      elsif ( not x21 and x23 and x22 and not x5 and not x18 ) = '1' then
         y1 <= '1' ;
         y5 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s97;

      elsif ( not x21 and x23 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x21 and not x23 and x22 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x23 and not x22 and x15 and x9 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x21 and not x23 and not x22 and x15 and not x9 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( not x21 and not x23 and not x22 and not x15 and x16 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      else
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s205;

      end if;

   when s121 =>
      if ( x67 and x22 and x3 and x15 and x8 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x67 and x22 and x3 and x15 and not x8 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s154;

      elsif ( x67 and x22 and x3 and not x15 and x16 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s255;

      elsif ( x67 and x22 and x3 and not x15 and not x16 ) = '1' then
         y3 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s6;

      elsif ( x67 and x22 and not x3 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s255;

      elsif ( x67 and not x22 and x23 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x67 and not x22 and x23 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x67 and not x22 and x23 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x22 and x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x22 and not x23 and x16 and x15 and x14 and x8 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( x67 and not x22 and not x23 and x16 and x15 and x14 and not x8 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x67 and not x22 and not x23 and x16 and x15 and not x14 and x7 and x8 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( x67 and not x22 and not x23 and x16 and x15 and not x14 and x7 and not x8 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s126;

      elsif ( x67 and not x22 and not x23 and x16 and x15 and not x14 and not x7 and x8 and x12 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s125;

      elsif ( x67 and not x22 and not x23 and x16 and x15 and not x14 and not x7 and x8 and not x12 and x18 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x67 and not x22 and not x23 and x16 and x15 and not x14 and not x7 and x8 and not x12 and x18 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x22 and not x23 and x16 and x15 and not x14 and not x7 and x8 and not x12 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x22 and not x23 and x16 and x15 and not x14 and not x7 and not x8 and x13 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s125;

      elsif ( x67 and not x22 and not x23 and x16 and x15 and not x14 and not x7 and not x8 and not x13 and x18 and x12 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x67 and not x22 and not x23 and x16 and x15 and not x14 and not x7 and not x8 and not x13 and x18 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x22 and not x23 and x16 and x15 and not x14 and not x7 and not x8 and not x13 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and x8 and x9 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and x8 and x9 and not x2 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and x8 and x9 and not x2 and not x3 ) = '1' then
         y4 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s111;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and x8 and not x9 and x7 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and x8 and not x9 and x7 and not x2 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and x8 and not x9 and x7 and not x2 and not x3 ) = '1' then
         y4 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s111;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and x8 and not x9 and not x7 and x18 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and x8 and not x9 and not x7 and x18 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and x8 and not x9 and not x7 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and x8 and not x9 and not x7 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and not x8 and x7 and x11 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and not x8 and x7 and x11 and not x2 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and not x8 and x7 and x11 and not x2 and not x3 ) = '1' then
         y4 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s111;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and not x8 and x7 and not x11 and x18 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and not x8 and x7 and not x11 and x18 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and not x8 and x7 and not x11 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and not x8 and x7 and not x11 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and not x8 and not x7 and x10 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and not x8 and not x7 and x10 and not x2 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and not x8 and not x7 and x10 and not x2 and not x3 ) = '1' then
         y4 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s111;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and not x8 and not x7 and not x10 and x18 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and not x8 and not x7 and not x10 and x18 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and not x8 and not x7 and not x10 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x22 and not x23 and x16 and not x15 and not x8 and not x7 and not x10 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x22 and not x23 and not x16 and x15 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x67 and not x22 and not x23 and not x16 and x15 and not x7 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( x67 and not x22 and not x23 and not x16 and x15 and not x7 and not x2 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x67 and not x22 and not x23 and not x16 and x15 and not x7 and not x2 and not x3 and x8 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s129;

      elsif ( x67 and not x22 and not x23 and not x16 and x15 and not x7 and not x2 and not x3 and not x8 ) = '1' then
         y9 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s111;

      elsif ( x67 and not x22 and not x23 and not x16 and not x15 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

      elsif ( x67 and not x22 and not x23 and not x16 and not x15 and not x2 and x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x67 and not x22 and not x23 and not x16 and not x15 and not x2 and not x3 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         y12 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s127;

      elsif ( not x67 and x21 and x20 and x15 and x10 and x11 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s192;

      elsif ( not x67 and x21 and x20 and x15 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s193;

      elsif ( not x67 and x21 and x20 and x15 and x10 and not x11 and not x12 ) = '1' then
         y1 <= '1' ;
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s194;

      elsif ( not x67 and x21 and x20 and x15 and not x10 and x12 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s300;

      elsif ( not x67 and x21 and x20 and x15 and not x10 and not x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s192;

      elsif ( not x67 and x21 and x20 and not x15 and x16 and x10 and x12 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s259;

      elsif ( not x67 and x21 and x20 and not x15 and x16 and x10 and not x12 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( not x67 and x21 and x20 and not x15 and x16 and not x10 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s259;

      elsif ( not x67 and x21 and x20 and not x15 and not x16 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( not x67 and x21 and not x20 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s57;

      elsif ( not x67 and not x21 and x4 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s306;

      elsif ( not x67 and not x21 and not x4 and x18 and x15 and x10 and x11 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x67 and not x21 and not x4 and x18 and x15 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s301;

      elsif ( not x67 and not x21 and not x4 and x18 and x15 and x10 and not x11 and not x12 ) = '1' then
         y8 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s195;

      elsif ( not x67 and not x21 and not x4 and x18 and x15 and not x10 and x12 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      elsif ( not x67 and not x21 and not x4 and x18 and x15 and not x10 and not x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s192;

      elsif ( not x67 and not x21 and not x4 and x18 and not x15 and x16 and x10 and x12 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s259;

      elsif ( not x67 and not x21 and not x4 and x18 and not x15 and x16 and x10 and not x12 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s302;

      elsif ( not x67 and not x21 and not x4 and x18 and not x15 and x16 and not x10 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s259;

      elsif ( not x67 and not x21 and not x4 and x18 and not x15 and not x16 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s303;

      else
         y5 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s57;

      end if;

   when s122 =>
      if ( x65 and x22 ) = '1' then
         y9 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s111;

      elsif ( x65 and not x22 and x23 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x65 and not x22 and not x23 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x68 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x68 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x68 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x68 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x68 and x23 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      else
         y11 <= '1' ;
         current_group15m <= s53;

      end if;

   when s123 =>
      if ( x21 and x9 and x3 ) = '1' then
         current_group15m <= s40;

      elsif ( x21 and x9 and not x3 and x4 ) = '1' then
         current_group15m <= s40;

      elsif ( x21 and x9 and not x3 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x5 and not x4 and x22 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x5 and not x4 and x22 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x5 and not x4 and not x22 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x5 and x22 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x5 and not x22 and x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and not x5 and not x22 and x4 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s124 =>
      if ( x65 and x22 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x22 and x23 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s255;

      elsif ( x65 and not x22 and not x23 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s389;

      elsif ( not x65 and x21 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x21 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x21 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and x7 and x8 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and not x21 and x22 and x7 and not x8 and x9 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and not x21 and x22 and x7 and not x8 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and not x22 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and not x21 and not x22 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and not x21 and not x22 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s125 =>
      if ( x67 and x22 ) = '1' then
         y2 <= '1' ;
         y16 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s124;

      elsif ( x67 and not x22 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s302;

      else
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s302;

      end if;

   when s126 =>
      if ( x65 and x67 and x22 and x17 and x18 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and x22 and x17 and not x18 and x19 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and x22 and x17 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and x22 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x22 and x18 and x13 and x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and x67 and not x22 and x18 and x13 and not x23 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x67 and not x22 and x18 and not x13 and x12 and x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and x67 and not x22 and x18 and not x13 and x12 and not x23 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x67 and not x22 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x22 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x21 and x20 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x67 and x21 and x20 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x67 and x21 and x20 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x21 and x20 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x21 and not x20 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and not x67 and x21 and not x20 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and not x67 and x21 and not x20 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x21 and not x20 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x21 and x19 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x67 and not x21 and x19 and not x14 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x67 and not x21 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x21 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s143;

      elsif ( not x65 and x66 and not x21 and x23 and x22 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x65 and x66 and not x21 and x23 and not x22 and x19 and x14 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x65 and x66 and not x21 and x23 and not x22 and x19 and not x14 and x13 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x65 and x66 and not x21 and x23 and not x22 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x21 and x23 and not x22 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x21 and not x23 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and not x66 and x67 and x20 and x18 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x66 and x67 and x20 and x18 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x66 and x67 and x20 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and x20 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and not x20 and x21 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x66 and x67 and not x20 and x21 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x66 and x67 and not x20 and x21 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and not x20 and x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and not x20 and not x21 and x17 and x13 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x65 and not x66 and x67 and not x20 and not x21 and x17 and not x13 and x12 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x65 and not x66 and x67 and not x20 and not x21 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x67 and not x20 and not x21 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and x21 and x19 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x67 and x21 and not x19 and x20 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s176;

      elsif ( not x65 and not x66 and not x67 and x21 and not x19 and not x20 ) = '1' then
         y17 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s377;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x19 and x13 and x20 and x15 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x19 and x13 and x20 and not x15 ) = '1' then
         y22 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s123;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x19 and x13 and not x20 ) = '1' then
         y2 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s371;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x19 and not x13 and x20 and x14 and x15 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s373;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x19 and not x13 and x20 and x14 and not x15 ) = '1' then
         y17 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s377;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x19 and not x13 and x20 and not x14 and x15 and x6 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s293;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x19 and not x13 and x20 and not x14 and x15 and not x6 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x19 and not x13 and x20 and not x14 and x15 and not x6 and x5 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x19 and not x13 and x20 and not x14 and x15 and not x6 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x19 and not x13 and x20 and not x14 and not x15 and x4 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s293;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x19 and not x13 and x20 and not x14 and not x15 and not x4 and x5 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x19 and not x13 and x20 and not x14 and not x15 and not x4 and x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x19 and not x13 and x20 and not x14 and not x15 and not x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x19 and not x13 and not x20 and x14 ) = '1' then
         y2 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s371;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x19 and not x13 and not x20 and not x14 and x7 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s329;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x19 and not x13 and not x20 and not x14 and not x7 and x8 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s103;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x19 and not x13 and not x20 and not x14 and not x7 and not x8 and x15 ) = '1' then
         y8 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s378;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and x19 and not x13 and not x20 and not x14 and not x7 and not x8 and not x15 ) = '1' then
         y2 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and not x19 and x7 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s329;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and not x19 and not x7 and x20 and x15 and x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and not x19 and not x7 and x20 and x15 and not x14 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s103;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and not x19 and not x7 and x20 and not x15 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s103;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and not x19 and not x7 and not x20 and x8 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s103;

      elsif ( not x65 and not x66 and not x67 and not x21 and x22 and not x19 and not x7 and not x20 and not x8 ) = '1' then
         y21 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s225;

      elsif ( not x65 and not x66 and not x67 and not x21 and not x22 and x4 and x5 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x67 and not x21 and not x22 and x4 and not x5 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x66 and not x67 and not x21 and not x22 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s127 =>
      if ( x22 and x17 and x18 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x22 and x17 and not x18 and x19 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x22 and x17 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x22 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x22 and x23 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      else
         y11 <= '1' ;
         current_group15m <= s53;

      end if;

   when s128 =>
      if ( x65 and x67 and x22 and x15 and x8 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x67 and x22 and x15 and not x8 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x65 and x67 and x22 and not x15 and x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s50;

      elsif ( x65 and x67 and x22 and not x15 and not x16 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s122;

      elsif ( x65 and x67 and not x22 and x15 and x8 and x23 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x67 and not x22 and x15 and x8 and not x23 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s8;

      elsif ( x65 and x67 and not x22 and x15 and not x8 and x23 and x6 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s111;

      elsif ( x65 and x67 and not x22 and x15 and not x8 and x23 and not x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x67 and not x22 and x15 and not x8 and not x23 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s111;

      elsif ( x65 and x67 and not x22 and not x15 and x16 and x23 and x8 and x7 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x67 and not x22 and not x15 and x16 and x23 and x8 and not x7 and x9 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x67 and not x22 and not x15 and x16 and x23 and x8 and not x7 and not x9 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and x67 and not x22 and not x15 and x16 and x23 and x8 and not x7 and not x9 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and x67 and not x22 and not x15 and x16 and x23 and x8 and not x7 and not x9 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x22 and not x15 and x16 and x23 and x8 and not x7 and not x9 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x22 and not x15 and x16 and x23 and not x8 and x7 and x11 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x67 and not x22 and not x15 and x16 and x23 and not x8 and x7 and not x11 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and x67 and not x22 and not x15 and x16 and x23 and not x8 and x7 and not x11 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and x67 and not x22 and not x15 and x16 and x23 and not x8 and x7 and not x11 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x22 and not x15 and x16 and x23 and not x8 and x7 and not x11 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x22 and not x15 and x16 and x23 and not x8 and not x7 and x10 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x67 and not x22 and not x15 and x16 and x23 and not x8 and not x7 and not x10 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and x67 and not x22 and not x15 and x16 and x23 and not x8 and not x7 and not x10 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and x67 and not x22 and not x15 and x16 and x23 and not x8 and not x7 and not x10 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x22 and not x15 and x16 and x23 and not x8 and not x7 and not x10 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x22 and not x15 and x16 and not x23 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s154;

      elsif ( x65 and x67 and not x22 and not x15 and not x16 and x23 and x6 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( x65 and x67 and not x22 and not x15 and not x16 and x23 and not x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x67 and not x22 and not x15 and not x16 and not x23 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( x65 and not x67 and x61 and x60 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s67;

      elsif ( x65 and not x67 and x61 and not x60 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      elsif ( x65 and not x67 and not x61 and x60 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      elsif ( x65 and not x67 and not x61 and not x60 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and x22 ) = '1' then
         y2 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s79;

      else
         y9 <= '1' ;
         current_group15m <= s27;

      end if;

   when s129 =>
      if ( x22 and x17 and x18 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x22 and x17 and not x18 and x19 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x22 and x17 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x22 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x22 and x23 and x15 and x8 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( not x22 and x23 and x15 and not x8 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x22 and x23 and not x15 and x16 ) = '1' then
         y4 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s111;

      elsif ( not x22 and x23 and not x15 and not x16 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s122;

      elsif ( not x22 and not x23 and x18 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( not x22 and not x23 and x18 and not x13 and x12 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( not x22 and not x23 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s130 =>
      if ( x65 and x22 ) = '1' then
         y2 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s121;

      elsif ( x65 and not x22 and x23 and x15 and x16 and x14 and x8 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( x65 and not x22 and x23 and x15 and x16 and x14 and not x8 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x65 and not x22 and x23 and x15 and x16 and not x14 and x7 and x8 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( x65 and not x22 and x23 and x15 and x16 and not x14 and x7 and not x8 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s126;

      elsif ( x65 and not x22 and x23 and x15 and x16 and not x14 and not x7 and x8 and x12 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s302;

      elsif ( x65 and not x22 and x23 and x15 and x16 and not x14 and not x7 and x8 and not x12 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and not x22 and x23 and x15 and x16 and not x14 and not x7 and x8 and not x12 and x18 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x22 and x23 and x15 and x16 and not x14 and not x7 and x8 and not x12 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x22 and x23 and x15 and x16 and not x14 and not x7 and not x8 and x13 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s302;

      elsif ( x65 and not x22 and x23 and x15 and x16 and not x14 and not x7 and not x8 and not x13 and x18 and x12 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and not x22 and x23 and x15 and x16 and not x14 and not x7 and not x8 and not x13 and x18 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x22 and x23 and x15 and x16 and not x14 and not x7 and not x8 and not x13 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x22 and x23 and x15 and not x16 and x7 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x65 and not x22 and x23 and x15 and not x16 and not x7 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s44;

      elsif ( x65 and not x22 and x23 and x15 and not x16 and not x7 and not x2 and x3 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s129;

      elsif ( x65 and not x22 and x23 and x15 and not x16 and not x7 and not x2 and not x3 and x8 ) = '1' then
         y2 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s121;

      elsif ( x65 and not x22 and x23 and x15 and not x16 and not x7 and not x2 and not x3 and not x8 ) = '1' then
         y9 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s111;

      elsif ( x65 and not x22 and x23 and not x15 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s44;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and x16 and x7 and x11 and x3 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s129;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and x16 and x7 and x11 and not x3 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s154;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and x16 and x7 and not x11 and x8 and x3 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s129;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and x16 and x7 and not x11 and x8 and not x3 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s154;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and x16 and x7 and not x11 and not x8 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and x16 and x7 and not x11 and not x8 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and x16 and x7 and not x11 and not x8 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and x16 and x7 and not x11 and not x8 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and x16 and not x7 and x8 and x9 and x3 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s129;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and x16 and not x7 and x8 and x9 and not x3 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s154;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and x16 and not x7 and x8 and not x9 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and x16 and not x7 and x8 and not x9 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and x16 and not x7 and x8 and not x9 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and x16 and not x7 and x8 and not x9 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and x16 and not x7 and not x8 and x10 and x3 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s129;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and x16 and not x7 and not x8 and x10 and not x3 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s154;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and x16 and not x7 and not x8 and not x10 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and x16 and not x7 and not x8 and not x10 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and x16 and not x7 and not x8 and not x10 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and x16 and not x7 and not x8 and not x10 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and not x16 and x3 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s129;

      elsif ( x65 and not x22 and x23 and not x15 and not x2 and not x16 and not x3 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         y12 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s127;

      elsif ( x65 and not x22 and not x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( not x65 and x67 and x15 and x8 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x65 and x67 and x15 and not x8 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x65 and x67 and not x15 and x16 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s151;

      elsif ( not x65 and x67 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s135;

      else
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      end if;

   when s131 =>
      if ( x68 and x6 and x15 and x10 and x11 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s301;

      elsif ( x68 and x6 and x15 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s192;

      elsif ( x68 and x6 and x15 and x10 and not x11 and not x12 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s60;

      elsif ( x68 and x6 and x15 and not x10 and x12 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s196;

      elsif ( x68 and x6 and x15 and not x10 and not x12 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s61;

      elsif ( x68 and x6 and not x15 and x16 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s60;

      elsif ( x68 and x6 and not x15 and not x16 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s303;

      elsif ( x68 and not x6 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s60;

      elsif ( not x68 and x60 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s68;

      else
         y11 <= '1' ;
         current_group15m <= s53;

      end if;

   when s132 =>
      if ( x21 and x15 and x20 and x10 and x11 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s192;

      elsif ( x21 and x15 and x20 and x10 and not x11 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s193;

      elsif ( x21 and x15 and x20 and not x10 and x12 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s300;

      elsif ( x21 and x15 and x20 and not x10 and not x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s192;

      elsif ( x21 and x15 and not x20 and x5 and x10 and x11 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s301;

      elsif ( x21 and x15 and not x20 and x5 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s192;

      elsif ( x21 and x15 and not x20 and x5 and x10 and not x11 and not x12 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( x21 and x15 and not x20 and x5 and not x10 and x12 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s196;

      elsif ( x21 and x15 and not x20 and x5 and not x10 and not x12 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s61;

      elsif ( x21 and x15 and not x20 and not x5 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( x21 and not x15 and x16 and x10 and x12 and x20 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s192;

      elsif ( x21 and not x15 and x16 and x10 and x12 and not x20 and x8 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( x21 and not x15 and x16 and x10 and x12 and not x20 and not x8 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x15 and x16 and x10 and x12 and not x20 and not x8 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x15 and x16 and x10 and x12 and not x20 and not x8 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x15 and x16 and x10 and x12 and not x20 and not x8 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x15 and x16 and x10 and not x12 and x20 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( x21 and not x15 and x16 and x10 and not x12 and not x20 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( x21 and not x15 and x16 and not x10 and x20 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s192;

      elsif ( x21 and not x15 and x16 and not x10 and not x20 and x12 and x7 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( x21 and not x15 and x16 and not x10 and not x20 and x12 and not x7 and x11 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( x21 and not x15 and x16 and not x10 and not x20 and x12 and not x7 and not x11 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x15 and x16 and not x10 and not x20 and x12 and not x7 and not x11 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x15 and x16 and not x10 and not x20 and x12 and not x7 and not x11 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x15 and x16 and not x10 and not x20 and x12 and not x7 and not x11 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x15 and x16 and not x10 and not x20 and not x12 and x11 and x9 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( x21 and not x15 and x16 and not x10 and not x20 and not x12 and x11 and not x9 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x15 and x16 and not x10 and not x20 and not x12 and x11 and not x9 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x15 and x16 and not x10 and not x20 and not x12 and x11 and not x9 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x15 and x16 and not x10 and not x20 and not x12 and x11 and not x9 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x15 and x16 and not x10 and not x20 and not x12 and not x11 and x8 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x15 and x16 and not x10 and not x20 and not x12 and not x11 and x8 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x15 and x16 and not x10 and not x20 and not x12 and not x11 and x8 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x15 and x16 and not x10 and not x20 and not x12 and not x11 and x8 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x15 and x16 and not x10 and not x20 and not x12 and not x11 and not x8 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( x21 and not x15 and not x16 and x20 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x21 and not x15 and not x16 and not x20 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x21 and not x15 and not x16 and not x20 and not x5 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x21 and x3 and x15 and x10 and x11 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s192;

      elsif ( not x21 and x3 and x15 and x10 and not x11 and x12 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s193;

      elsif ( not x21 and x3 and x15 and x10 and not x11 and not x12 ) = '1' then
         y1 <= '1' ;
         y8 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s192;

      elsif ( not x21 and x3 and x15 and not x10 and x12 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s300;

      elsif ( not x21 and x3 and x15 and not x10 and not x12 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s198;

      elsif ( not x21 and x3 and not x15 and x16 ) = '1' then
         y2 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s121;

      elsif ( not x21 and x3 and not x15 and not x16 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s390;

      else
         y2 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s121;

      end if;

   when s133 =>
      if ( x65 and x66 and x20 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and x20 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x66 and x20 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and x20 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x66 and not x20 and x15 and x10 and x11 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s192;

      elsif ( x65 and x66 and not x20 and x15 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s193;

      elsif ( x65 and x66 and not x20 and x15 and x10 and not x11 and not x12 ) = '1' then
         y1 <= '1' ;
         y8 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s192;

      elsif ( x65 and x66 and not x20 and x15 and not x10 and x12 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s300;

      elsif ( x65 and x66 and not x20 and x15 and not x10 and not x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s192;

      elsif ( x65 and x66 and not x20 and not x15 and x16 and x10 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s306;

      elsif ( x65 and x66 and not x20 and not x15 and x16 and not x10 and x12 and x11 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s259;

      elsif ( x65 and x66 and not x20 and not x15 and x16 and not x10 and x12 and not x11 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s306;

      elsif ( x65 and x66 and not x20 and not x15 and x16 and not x10 and not x12 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s306;

      elsif ( x65 and x66 and not x20 and not x15 and not x16 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s201;

      elsif ( x65 and not x66 and x21 and x68 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x65 and not x66 and x21 and not x68 and x7 and x16 and x13 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and x21 and not x68 and x7 and x16 and not x13 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and x21 and not x68 and x7 and not x16 and x17 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and x21 and not x68 and x7 and not x16 and not x17 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and x21 and not x68 and not x7 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and x22 and x68 and x8 and x23 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x66 and not x21 and x22 and x68 and x8 and x23 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x66 and not x21 and x22 and x68 and x8 and x23 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and x68 and x8 and not x23 and x9 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x66 and not x21 and x22 and x68 and x8 and not x23 and not x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x66 and not x21 and x22 and x68 and x8 and not x23 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and x68 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and x16 and x18 and x19 and x10 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and x16 and x18 and x19 and not x10 and x7 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and x16 and x18 and x19 and not x10 and not x7 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and x16 and x18 and not x19 and x7 and x13 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and x16 and x18 and not x19 and x7 and not x13 ) = '1' then
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and x16 and x18 and not x19 and not x7 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and x16 and not x18 and x13 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and x16 and not x18 and not x13 and x7 and x19 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s362;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and x16 and not x18 and not x13 and x7 and not x19 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and x16 and not x18 and not x13 and not x7 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and x18 and x19 and x10 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and x18 and x19 and not x10 and x15 and x12 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and x18 and x19 and not x10 and x15 and not x12 and x14 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and x18 and x19 and not x10 and x15 and not x12 and not x14 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and x18 and x19 and not x10 and x15 and not x12 and not x14 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and x18 and x19 and not x10 and x15 and not x12 and not x14 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and x18 and x19 and not x10 and x15 and not x12 and not x14 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and x18 and x19 and not x10 and not x15 and x14 and x13 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and x18 and x19 and not x10 and not x15 and x14 and not x13 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and x18 and x19 and not x10 and not x15 and x14 and not x13 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and x18 and x19 and not x10 and not x15 and x14 and not x13 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and x18 and x19 and not x10 and not x15 and x14 and not x13 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and x18 and x19 and not x10 and not x15 and not x14 and x11 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and x18 and x19 and not x10 and not x15 and not x14 and not x11 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and x18 and x19 and not x10 and not x15 and not x14 and not x11 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and x18 and x19 and not x10 and not x15 and not x14 and not x11 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and x18 and x19 and not x10 and not x15 and not x14 and not x11 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and x18 and not x19 and x7 and x13 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and x18 and not x19 and x7 and not x13 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and x18 and not x19 and not x7 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and x13 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and x15 and x11 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and x15 and not x11 and x14 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and x15 and not x11 and not x14 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and x15 and not x11 and not x14 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and x15 and not x11 and not x14 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and x15 and not x11 and not x14 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and not x15 and x14 and x12 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and not x15 and x14 and not x12 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and not x15 and x14 and not x12 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and not x15 and x14 and not x12 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and not x15 and x14 and not x12 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and not x15 and not x14 and x10 and x19 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and not x15 and not x14 and x10 and not x19 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and not x15 and not x14 and x10 and not x19 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and not x15 and not x14 and x10 and not x19 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and not x15 and not x14 and x10 and not x19 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and not x15 and not x14 and not x10 and x19 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and not x15 and not x14 and not x10 and x19 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and not x15 and not x14 and not x10 and x19 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and not x15 and not x14 and not x10 and x19 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and x17 and not x18 and not x13 and not x15 and not x14 and not x10 and not x19 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and not x17 and x7 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and x22 and not x68 and not x16 and not x17 and not x7 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and not x22 and x68 and x23 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x66 and not x21 and not x22 and x68 and x23 and x9 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x66 and not x21 and not x22 and x68 and x23 and x9 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x22 and x68 and x23 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x22 and x68 and not x23 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x66 and not x21 and not x22 and x68 and not x23 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x66 and not x21 and not x22 and x68 and not x23 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x22 and x68 and not x23 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and x17 and x13 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and x17 and not x13 and x7 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s362;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and x17 and not x13 and not x7 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and not x17 and x18 and x13 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and not x17 and x18 and not x13 and x15 and x11 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and not x17 and x18 and not x13 and x15 and not x11 and x14 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and not x17 and x18 and not x13 and x15 and not x11 and not x14 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and not x17 and x18 and not x13 and x15 and not x11 and not x14 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and not x17 and x18 and not x13 and x15 and not x11 and not x14 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and not x17 and x18 and not x13 and x15 and not x11 and not x14 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and not x17 and x18 and not x13 and not x15 and x14 and x12 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and not x17 and x18 and not x13 and not x15 and x14 and not x12 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and not x17 and x18 and not x13 and not x15 and x14 and not x12 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and not x17 and x18 and not x13 and not x15 and x14 and not x12 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and not x17 and x18 and not x13 and not x15 and x14 and not x12 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and not x17 and x18 and not x13 and not x15 and not x14 and x10 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and not x17 and x18 and not x13 and not x15 and not x14 and not x10 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and not x17 and x18 and not x13 and not x15 and not x14 and not x10 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and not x17 and x18 and not x13 and not x15 and not x14 and not x10 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and not x17 and x18 and not x13 and not x15 and not x14 and not x10 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and not x17 and not x18 and x7 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and x19 and not x17 and not x18 and not x7 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and not x19 and x16 and x13 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and not x19 and x16 and not x13 and x7 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and not x19 and x16 and not x13 and not x7 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and not x19 and not x16 and x17 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and not x19 and not x16 and not x17 and x7 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s146;

      elsif ( x65 and not x66 and not x21 and not x22 and not x68 and not x19 and not x16 and not x17 and not x7 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s391;

      elsif ( not x65 and x20 and x18 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x20 and x18 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x20 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x20 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x20 and x21 and x15 and x16 and x14 and x8 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s126;

      elsif ( not x65 and not x20 and x21 and x15 and x16 and x14 and not x8 ) = '1' then
         y1 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y13 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s207;

      elsif ( not x65 and not x20 and x21 and x15 and x16 and not x14 and x7 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s210;

      elsif ( not x65 and not x20 and x21 and x15 and x16 and not x14 and x7 and not x8 ) = '1' then
         y7 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s211;

      elsif ( not x65 and not x20 and x21 and x15 and x16 and not x14 and not x7 and x8 and x12 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s279;

      elsif ( not x65 and not x20 and x21 and x15 and x16 and not x14 and not x7 and x8 and not x12 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x20 and x21 and x15 and x16 and not x14 and not x7 and x8 and not x12 and x18 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x20 and x21 and x15 and x16 and not x14 and not x7 and x8 and not x12 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x20 and x21 and x15 and x16 and not x14 and not x7 and not x8 and x13 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s279;

      elsif ( not x65 and not x20 and x21 and x15 and x16 and not x14 and not x7 and not x8 and not x13 and x18 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x20 and x21 and x15 and x16 and not x14 and not x7 and not x8 and not x13 and x18 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x20 and x21 and x15 and x16 and not x14 and not x7 and not x8 and not x13 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x20 and x21 and x15 and not x16 and x7 and x8 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x65 and not x20 and x21 and x15 and not x16 and x7 and not x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and not x20 and x21 and x15 and not x16 and not x7 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s392;

      elsif ( not x65 and not x20 and x21 and x15 and not x16 and not x7 and not x2 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s41;

      elsif ( not x65 and not x20 and x21 and x15 and not x16 and not x7 and not x2 and not x3 and x8 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x20 and x21 and x15 and not x16 and not x7 and not x2 and not x3 and not x8 ) = '1' then
         y2 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s206;

      elsif ( not x65 and not x20 and x21 and not x15 and x2 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s392;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and x16 and x7 and x11 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s41;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and x16 and x7 and x11 and not x3 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and x16 and x7 and not x11 and x8 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s41;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and x16 and x7 and not x11 and x8 and not x3 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and x16 and x7 and not x11 and not x8 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and x16 and x7 and not x11 and not x8 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and x16 and x7 and not x11 and not x8 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and x16 and x7 and not x11 and not x8 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and x16 and not x7 and x8 and x9 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s41;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and x16 and not x7 and x8 and x9 and not x3 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and x16 and not x7 and x8 and not x9 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and x16 and not x7 and x8 and not x9 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and x16 and not x7 and x8 and not x9 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and x16 and not x7 and x8 and not x9 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and x16 and not x7 and not x8 and x10 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s41;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and x16 and not x7 and not x8 and x10 and not x3 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and x16 and not x7 and not x8 and not x10 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and x16 and not x7 and not x8 and not x10 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and x16 and not x7 and not x8 and not x10 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and x16 and not x7 and not x8 and not x10 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and not x16 and x3 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s41;

      elsif ( not x65 and not x20 and x21 and not x15 and not x2 and not x16 and not x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s393;

      elsif ( not x65 and not x20 and not x21 and x6 and x15 and x8 ) = '1' then
         y2 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s366;

      elsif ( not x65 and not x20 and not x21 and x6 and x15 and not x8 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s207;

      elsif ( not x65 and not x20 and not x21 and x6 and not x15 and x16 ) = '1' then
         y2 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s366;

      elsif ( not x65 and not x20 and not x21 and x6 and not x15 and not x16 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s393;

      else
         y2 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s366;

      end if;

   when s134 =>
      if ( x21 and x20 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x20 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x20 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x20 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x20 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x20 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x20 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x20 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x15 and x10 and x11 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x21 and x15 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s301;

      elsif ( not x21 and x15 and x10 and not x11 and not x12 ) = '1' then
         y8 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s195;

      elsif ( not x21 and x15 and not x10 and x12 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      elsif ( not x21 and x15 and not x10 and not x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s192;

      elsif ( not x21 and not x15 and x16 and x10 and x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s192;

      elsif ( not x21 and not x15 and x16 and x10 and not x12 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s302;

      elsif ( not x21 and not x15 and x16 and not x10 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s192;

      else
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s303;

      end if;

   when s135 =>
      if ( x62 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s159;

      else
         y15 <= '1' ;
         current_group15m <= s149;

      end if;

   when s136 =>
      if ( x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x23 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x23 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 and x18 and x19 and x15 and x17 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( not x21 and x22 and not x23 and x18 and x19 and x15 and not x17 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x21 and x22 and not x23 and x18 and x19 and not x15 and x16 and x17 ) = '1' then
         y24 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s157;

      elsif ( not x21 and x22 and not x23 and x18 and x19 and not x15 and x16 and not x17 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         y20 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s227;

      elsif ( not x21 and x22 and not x23 and x18 and x19 and not x15 and not x16 and x8 and x9 and x17 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and not x23 and x18 and x19 and not x15 and not x16 and x8 and x9 and not x17 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s117;

      elsif ( not x21 and x22 and not x23 and x18 and x19 and not x15 and not x16 and x8 and not x9 and x10 and x17 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s117;

      elsif ( not x21 and x22 and not x23 and x18 and x19 and not x15 and not x16 and x8 and not x9 and x10 and not x17 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and not x23 and x18 and x19 and not x15 and not x16 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 and x18 and x19 and not x15 and not x16 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 and x18 and not x19 and x16 and x15 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s203;

      elsif ( not x21 and x22 and not x23 and x18 and not x19 and x16 and not x15 and x17 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x21 and x22 and not x23 and x18 and not x19 and x16 and not x15 and not x17 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s233;

      elsif ( not x21 and x22 and not x23 and x18 and not x19 and not x16 and x17 and x15 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s234;

      elsif ( not x21 and x22 and not x23 and x18 and not x19 and not x16 and x17 and not x15 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s235;

      elsif ( not x21 and x22 and not x23 and x18 and not x19 and not x16 and not x17 and x5 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s31;

      elsif ( not x21 and x22 and not x23 and x18 and not x19 and not x16 and not x17 and not x5 and x3 ) = '1' then
         y15 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s36;

      elsif ( not x21 and x22 and not x23 and x18 and not x19 and not x16 and not x17 and not x5 and not x3 and x15 ) = '1' then
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s227;

      elsif ( not x21 and x22 and not x23 and x18 and not x19 and not x16 and not x17 and not x5 and not x3 and not x15 ) = '1' then
         y16 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s227;

      elsif ( not x21 and x22 and not x23 and not x18 and x19 and x15 and x5 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s31;

      elsif ( not x21 and x22 and not x23 and not x18 and x19 and x15 and not x5 and x3 ) = '1' then
         y15 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s36;

      elsif ( not x21 and x22 and not x23 and not x18 and x19 and x15 and not x5 and not x3 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s228;

      elsif ( not x21 and x22 and not x23 and not x18 and x19 and not x15 and x16 and x14 and x5 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s31;

      elsif ( not x21 and x22 and not x23 and not x18 and x19 and not x15 and x16 and x14 and not x5 and x3 ) = '1' then
         y15 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s36;

      elsif ( not x21 and x22 and not x23 and not x18 and x19 and not x15 and x16 and x14 and not x5 and not x3 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x21 and x22 and not x23 and not x18 and x19 and not x15 and x16 and not x14 and x17 and x5 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s31;

      elsif ( not x21 and x22 and not x23 and not x18 and x19 and not x15 and x16 and not x14 and x17 and not x5 and x3 ) = '1' then
         y15 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s36;

      elsif ( not x21 and x22 and not x23 and not x18 and x19 and not x15 and x16 and not x14 and x17 and not x5 and not x3 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x21 and x22 and not x23 and not x18 and x19 and not x15 and x16 and not x14 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 and not x18 and x19 and not x15 and not x16 and x17 and x13 and x5 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s31;

      elsif ( not x21 and x22 and not x23 and not x18 and x19 and not x15 and not x16 and x17 and x13 and not x5 and x3 ) = '1' then
         y15 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s36;

      elsif ( not x21 and x22 and not x23 and not x18 and x19 and not x15 and not x16 and x17 and x13 and not x5 and not x3 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x21 and x22 and not x23 and not x18 and x19 and not x15 and not x16 and x17 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 and not x18 and x19 and not x15 and not x16 and not x17 and x12 and x5 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s31;

      elsif ( not x21 and x22 and not x23 and not x18 and x19 and not x15 and not x16 and not x17 and x12 and not x5 and x3 ) = '1' then
         y15 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s36;

      elsif ( not x21 and x22 and not x23 and not x18 and x19 and not x15 and not x16 and not x17 and x12 and not x5 and not x3 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x21 and x22 and not x23 and not x18 and x19 and not x15 and not x16 and not x17 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 and not x18 and not x19 and x5 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s31;

      elsif ( not x21 and x22 and not x23 and not x18 and not x19 and not x5 and x3 ) = '1' then
         y15 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s36;

      elsif ( not x21 and x22 and not x23 and not x18 and not x19 and not x5 and not x3 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      else
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s161;

      end if;

   when s137 =>
      if ( x21 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x21 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x21 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 ) = '1' then
         current_group15m <= s1;

      else
         y17 <= '1' ;
         current_group15m <= s77;

      end if;

   when s138 =>
      if ( x21 and x19 and x20 and x17 and x5 ) = '1' then
         y23 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s269;

      elsif ( x21 and x19 and x20 and x17 and not x5 and x3 and x4 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( x21 and x19 and x20 and x17 and not x5 and x3 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x19 and x20 and x17 and not x5 and not x3 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x19 and x20 and not x17 and x4 ) = '1' then
         y4 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s273;

      elsif ( x21 and x19 and x20 and not x17 and not x4 and x3 and x5 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( x21 and x19 and x20 and not x17 and not x4 and x3 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x19 and x20 and not x17 and not x4 and not x3 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x19 and not x20 and x12 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( x21 and x19 and not x20 and x12 and not x2 and x17 and x8 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( x21 and x19 and not x20 and x12 and not x2 and x17 and not x8 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s272;

      elsif ( x21 and x19 and not x20 and x12 and not x2 and not x17 and x8 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( x21 and x19 and not x20 and x12 and not x2 and not x17 and not x8 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s172;

      elsif ( x21 and x19 and not x20 and not x12 and x16 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x21 and x19 and not x20 and not x12 and not x16 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s62;

      elsif ( x21 and x19 and not x20 and not x12 and not x16 and not x2 and x8 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( x21 and x19 and not x20 and not x12 and not x16 and not x2 and not x8 and x17 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s234;

      elsif ( x21 and x19 and not x20 and not x12 and not x16 and not x2 and not x8 and not x17 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s374;

      elsif ( x21 and not x19 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s328;

      elsif ( x21 and not x19 and not x2 and x20 and x12 and x8 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( x21 and not x19 and not x2 and x20 and x12 and not x8 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s272;

      elsif ( x21 and not x19 and not x2 and x20 and not x12 and x17 and x16 and x8 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( x21 and not x19 and not x2 and x20 and not x12 and x17 and x16 and not x8 ) = '1' then
         y10 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s273;

      elsif ( x21 and not x19 and not x2 and x20 and not x12 and x17 and not x16 and x14 and x8 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( x21 and not x19 and not x2 and x20 and not x12 and x17 and not x16 and x14 and not x8 ) = '1' then
         y10 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s273;

      elsif ( x21 and not x19 and not x2 and x20 and not x12 and x17 and not x16 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x19 and not x2 and x20 and not x12 and not x17 and x16 and x15 and x8 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( x21 and not x19 and not x2 and x20 and not x12 and not x17 and x16 and x15 and not x8 ) = '1' then
         y10 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s273;

      elsif ( x21 and not x19 and not x2 and x20 and not x12 and not x17 and x16 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x19 and not x2 and x20 and not x12 and not x17 and not x16 and x13 and x8 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( x21 and not x19 and not x2 and x20 and not x12 and not x17 and not x16 and x13 and not x8 ) = '1' then
         y10 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s273;

      elsif ( x21 and not x19 and not x2 and x20 and not x12 and not x17 and not x16 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x19 and not x2 and not x20 and x8 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( x21 and not x19 and not x2 and not x20 and not x8 and x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s394;

      elsif ( x21 and not x19 and not x2 and not x20 and not x8 and not x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s203;

      elsif ( not x21 and x22 ) = '1' then
         current_group15m <= s1;

      else
         y18 <= '1' ;
         current_group15m <= s114;

      end if;

   when s139 =>
         y7 <= '1' ;
         current_group15m <= s30;

   when s140 =>
      if ( x65 and x66 and x68 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x65 and x66 and not x68 and x60 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and x62 and x20 ) = '1' then
         y2 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s367;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and x62 and not x20 and x16 and x11 and x12 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s153;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and x62 and not x20 and x16 and x11 and not x12 and x13 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s153;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and x62 and not x20 and x16 and x11 and not x12 and not x13 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s154;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and x62 and not x20 and x16 and not x11 and x13 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s63;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and x62 and not x20 and x16 and not x11 and not x13 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and x62 and not x20 and not x16 and x17 and x11 and x13 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and x62 and not x20 and not x16 and x17 and x11 and not x13 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and x62 and not x20 and not x16 and x17 and not x11 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and x62 and not x20 and not x16 and not x17 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( x65 and x66 and not x68 and not x60 and x61 and not x62 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x65 and x66 and not x68 and not x60 and not x61 ) = '1' then
         y2 <= '1' ;
         y19 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s321;

      elsif ( x65 and not x66 and x67 and x21 and x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x65 and not x66 and x67 and x21 and x8 and not x9 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x65 and not x66 and x67 and x21 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and x21 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and not x21 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s32;

      elsif ( x65 and not x66 and not x67 and x20 and x19 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x20 and x19 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x20 and x19 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x20 and x19 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x20 and not x19 ) = '1' then
         y6 <= '1' ;
         y8 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and not x20 ) = '1' then
         y6 <= '1' ;
         y8 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s1;

      elsif ( not x65 and x67 and x68 and x21 and x19 and x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and x67 and x68 and x21 and x19 and not x15 and x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and x67 and x68 and x21 and x19 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x68 and x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x68 and not x21 and x20 and x15 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( not x65 and x67 and x68 and not x21 and x20 and not x15 and x14 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( not x65 and x67 and x68 and not x21 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x68 and not x21 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and not x68 and x62 and x61 and x13 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and x67 and not x68 and x62 and x61 and not x13 and x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and x67 and not x68 and x62 and x61 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and not x68 and x62 and not x61 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and not x68 and not x62 and x63 and x17 and x13 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and x67 and not x68 and not x62 and x63 and x17 and not x13 and x12 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and x67 and not x68 and not x62 and x63 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and not x68 and not x62 and x63 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and not x68 and not x62 and not x63 and x64 and x4 ) = '1' then
         y31 <= '1' ;
         current_group15m <= s96;

      elsif ( not x65 and x67 and not x68 and not x62 and not x63 and x64 and not x4 and x18 and x16 and x8 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and x67 and not x68 and not x62 and not x63 and x64 and not x4 and x18 and x16 and not x8 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x65 and x67 and not x68 and not x62 and not x63 and x64 and not x4 and x18 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s135;

      elsif ( not x65 and x67 and not x68 and not x62 and not x63 and x64 and not x4 and not x18 ) = '1' then
         y14 <= '1' ;
         y28 <= '1' ;
         y32 <= '1' ;
         y33 <= '1' ;
         current_group15m <= s18;

      elsif ( not x65 and x67 and not x68 and not x62 and not x63 and not x64 and x19 and x13 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x67 and not x68 and not x62 and not x63 and not x64 and x19 and not x13 and x12 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x67 and not x68 and not x62 and not x63 and not x64 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and not x68 and not x62 and not x63 and not x64 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and x21 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s143;

      elsif ( not x65 and not x67 and not x21 and x23 and x22 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x65 and not x67 and not x21 and x23 and not x22 and x19 and x14 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x65 and not x67 and not x21 and x23 and not x22 and x19 and not x14 and x13 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x65 and not x67 and not x21 and x23 and not x22 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and x23 and not x22 and not x19 ) = '1' then
         current_group15m <= s1;

      else
         y12 <= '1' ;
         current_group15m <= s100;

      end if;

   when s141 =>
      if ( x21 and x20 and x16 and x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s113;

      elsif ( x21 and x20 and x16 and not x10 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x21 and x20 and not x16 and x17 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( x21 and x20 and not x16 and not x17 ) = '1' then
         y5 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s115;

      elsif ( x21 and not x20 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s317;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s317;

      end if;

   when s142 =>
      if ( x66 and x16 and x17 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and x16 and x17 and x8 and not x10 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x66 and x16 and x17 and not x8 and x9 and x10 ) = '1' then
         y23 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s269;

      elsif ( x66 and x16 and x17 and not x8 and x9 and not x10 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s113;

      elsif ( x66 and x16 and x17 and not x8 and not x9 and x21 and x10 and x14 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s188;

      elsif ( x66 and x16 and x17 and not x8 and not x9 and x21 and x10 and not x14 and x19 and x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and x16 and x17 and not x8 and not x9 and x21 and x10 and not x14 and x19 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x16 and x17 and not x8 and not x9 and x21 and x10 and not x14 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x16 and x17 and not x8 and not x9 and x21 and not x10 and x15 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s188;

      elsif ( x66 and x16 and x17 and not x8 and not x9 and x21 and not x10 and not x15 and x19 and x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and x16 and x17 and not x8 and not x9 and x21 and not x10 and not x15 and x19 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x16 and x17 and not x8 and not x9 and x21 and not x10 and not x15 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x16 and x17 and not x8 and not x9 and not x21 and x10 and x14 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s188;

      elsif ( x66 and x16 and x17 and not x8 and not x9 and not x21 and x10 and not x14 and x20 and x15 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x66 and x16 and x17 and not x8 and not x9 and not x21 and x10 and not x14 and x20 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x16 and x17 and not x8 and not x9 and not x21 and x10 and not x14 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x16 and x17 and not x8 and not x9 and not x21 and not x10 and x15 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s188;

      elsif ( x66 and x16 and x17 and not x8 and not x9 and not x21 and not x10 and not x15 and x20 and x14 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x66 and x16 and x17 and not x8 and not x9 and not x21 and not x10 and not x15 and x20 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x16 and x17 and not x8 and not x9 and not x21 and not x10 and not x15 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x16 and not x17 and x9 and x21 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s344;

      elsif ( x66 and x16 and not x17 and x9 and not x21 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( x66 and x16 and not x17 and not x9 and x8 and x21 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s344;

      elsif ( x66 and x16 and not x17 and not x9 and x8 and not x21 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( x66 and x16 and not x17 and not x9 and not x8 and x2 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( x66 and x16 and not x17 and not x9 and not x8 and not x2 and x21 and x3 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x66 and x16 and not x17 and not x9 and not x8 and not x2 and x21 and not x3 and x10 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x66 and x16 and not x17 and not x9 and not x8 and not x2 and x21 and not x3 and not x10 ) = '1' then
         y4 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s395;

      elsif ( x66 and x16 and not x17 and not x9 and not x8 and not x2 and not x21 and x3 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and x16 and not x17 and not x9 and not x8 and not x2 and not x21 and not x3 and x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s113;

      elsif ( x66 and x16 and not x17 and not x9 and not x8 and not x2 and not x21 and not x3 and not x10 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x66 and not x16 and x2 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( x66 and not x16 and not x2 and x17 and x10 and x11 ) = '1' then
         y7 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s211;

      elsif ( x66 and not x16 and not x2 and x17 and x10 and not x11 and x9 ) = '1' then
         y7 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s211;

      elsif ( x66 and not x16 and not x2 and x17 and x10 and not x11 and not x9 and x21 and x19 and x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and not x16 and not x2 and x17 and x10 and not x11 and not x9 and x21 and x19 and not x15 and x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and not x16 and not x2 and x17 and x10 and not x11 and not x9 and x21 and x19 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and not x2 and x17 and x10 and not x11 and not x9 and x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and not x2 and x17 and x10 and not x11 and not x9 and not x21 and x20 and x15 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x66 and not x16 and not x2 and x17 and x10 and not x11 and not x9 and not x21 and x20 and not x15 and x14 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x66 and not x16 and not x2 and x17 and x10 and not x11 and not x9 and not x21 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and not x2 and x17 and x10 and not x11 and not x9 and not x21 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and not x2 and x17 and not x10 and x9 and x13 ) = '1' then
         y7 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s211;

      elsif ( x66 and not x16 and not x2 and x17 and not x10 and x9 and not x13 and x21 and x19 and x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and not x16 and not x2 and x17 and not x10 and x9 and not x13 and x21 and x19 and not x15 and x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and not x16 and not x2 and x17 and not x10 and x9 and not x13 and x21 and x19 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and not x2 and x17 and not x10 and x9 and not x13 and x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and not x2 and x17 and not x10 and x9 and not x13 and not x21 and x20 and x15 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x66 and not x16 and not x2 and x17 and not x10 and x9 and not x13 and not x21 and x20 and not x15 and x14 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x66 and not x16 and not x2 and x17 and not x10 and x9 and not x13 and not x21 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and not x2 and x17 and not x10 and x9 and not x13 and not x21 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and not x2 and x17 and not x10 and not x9 and x12 ) = '1' then
         y7 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s211;

      elsif ( x66 and not x16 and not x2 and x17 and not x10 and not x9 and not x12 and x21 and x19 and x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and not x16 and not x2 and x17 and not x10 and not x9 and not x12 and x21 and x19 and not x15 and x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and not x16 and not x2 and x17 and not x10 and not x9 and not x12 and x21 and x19 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and not x2 and x17 and not x10 and not x9 and not x12 and x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and not x2 and x17 and not x10 and not x9 and not x12 and not x21 and x20 and x15 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x66 and not x16 and not x2 and x17 and not x10 and not x9 and not x12 and not x21 and x20 and not x15 and x14 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x66 and not x16 and not x2 and x17 and not x10 and not x9 and not x12 and not x21 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and not x2 and x17 and not x10 and not x9 and not x12 and not x21 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and not x2 and not x17 and x3 and x21 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x66 and not x16 and not x2 and not x17 and x3 and not x21 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and not x16 and not x2 and not x17 and not x3 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s279;

      elsif ( not x66 and x21 and x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s328;

      elsif ( not x66 and x21 and not x19 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s396;

      elsif ( not x66 and not x21 and x22 and x18 and x17 and x12 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s271;

      elsif ( not x66 and not x21 and x22 and x18 and x17 and not x12 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s271;

      elsif ( not x66 and not x21 and x22 and x18 and not x17 and x12 ) = '1' then
         y6 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s386;

      elsif ( not x66 and not x21 and x22 and x18 and not x17 and not x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s374;

      elsif ( not x66 and not x21 and x22 and not x18 and x19 and x12 and x17 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s271;

      elsif ( not x66 and not x21 and x22 and not x18 and x19 and x12 and not x17 ) = '1' then
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s388;

      elsif ( not x66 and not x21 and x22 and not x18 and x19 and not x12 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( not x66 and not x21 and x22 and not x18 and not x19 and x12 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s271;

      elsif ( not x66 and not x21 and x22 and not x18 and not x19 and not x12 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      else
         current_group15m <= s1;

      end if;

   when s143 =>
      if ( x21 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x23 and x15 and x10 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( not x21 and x23 and x15 and not x10 and x12 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x21 and x23 and x15 and not x10 and not x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s285;

      elsif ( not x21 and x23 and not x15 and x16 and x10 and x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s286;

      elsif ( not x21 and x23 and not x15 and x16 and x10 and not x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x21 and x23 and not x15 and x16 and not x10 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s286;

      elsif ( not x21 and x23 and not x15 and not x16 ) = '1' then
         current_group15m <= s40;

      elsif ( not x21 and not x23 and x15 and x10 and x11 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s334;

      elsif ( not x21 and not x23 and x15 and x10 and not x11 and x12 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s334;

      elsif ( not x21 and not x23 and x15 and x10 and not x11 and not x12 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x21 and not x23 and x15 and not x10 and x12 and x11 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      elsif ( not x21 and not x23 and x15 and not x10 and x12 and not x11 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x21 and not x23 and x15 and not x10 and not x12 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      elsif ( not x21 and not x23 and not x15 and x16 and x10 and x12 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x21 and not x23 and not x15 and x16 and x10 and not x12 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s341;

      elsif ( not x21 and not x23 and not x15 and x16 and not x10 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      else
         y3 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s81;

      end if;

   when s144 =>
      if ( x65 and x21 and x20 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x21 and x20 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x21 and x20 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x21 and x20 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x21 and not x20 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x21 and not x20 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x21 and not x20 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x21 and not x20 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x19 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x21 and x19 and not x14 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x21 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x21 and x22 and x23 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and x66 and not x21 and x22 and x23 and x17 and not x14 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and x66 and not x21 and x22 and x23 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x21 and x22 and x23 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x21 and x22 and not x23 and x19 ) = '1' then
         y4 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s304;

      elsif ( not x65 and x66 and not x21 and x22 and not x23 and not x19 and x20 and x15 and x10 and x11 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s334;

      elsif ( not x65 and x66 and not x21 and x22 and not x23 and not x19 and x20 and x15 and x10 and not x11 and x12 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s334;

      elsif ( not x65 and x66 and not x21 and x22 and not x23 and not x19 and x20 and x15 and x10 and not x11 and not x12 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and x66 and not x21 and x22 and not x23 and not x19 and x20 and x15 and not x10 and x12 and x11 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      elsif ( not x65 and x66 and not x21 and x22 and not x23 and not x19 and x20 and x15 and not x10 and x12 and not x11 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x65 and x66 and not x21 and x22 and not x23 and not x19 and x20 and x15 and not x10 and not x12 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      elsif ( not x65 and x66 and not x21 and x22 and not x23 and not x19 and x20 and not x15 and x16 and x10 and x12 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and x66 and not x21 and x22 and not x23 and not x19 and x20 and not x15 and x16 and x10 and not x12 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s341;

      elsif ( not x65 and x66 and not x21 and x22 and not x23 and not x19 and x20 and not x15 and x16 and not x10 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and x66 and not x21 and x22 and not x23 and not x19 and x20 and not x15 and not x16 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s81;

      elsif ( not x65 and x66 and not x21 and x22 and not x23 and not x19 and not x20 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x65 and x66 and not x21 and not x22 and x23 and x3 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s320;

      elsif ( not x65 and x66 and not x21 and not x22 and x23 and not x3 and x18 and x15 and x7 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s81;

      elsif ( not x65 and x66 and not x21 and not x22 and x23 and not x3 and x18 and x15 and not x7 and x9 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and x66 and not x21 and not x22 and x23 and not x3 and x18 and x15 and not x7 and not x9 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x66 and not x21 and not x22 and x23 and not x3 and x18 and not x15 and x7 and x9 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s330;

      elsif ( not x65 and x66 and not x21 and not x22 and x23 and not x3 and x18 and not x15 and x7 and not x9 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( not x65 and x66 and not x21 and not x22 and x23 and not x3 and x18 and not x15 and not x7 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s330;

      elsif ( not x65 and x66 and not x21 and not x22 and x23 and not x3 and not x18 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s84;

      elsif ( not x65 and x66 and not x21 and not x22 and not x23 and x15 and x7 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s81;

      elsif ( not x65 and x66 and not x21 and not x22 and not x23 and x15 and not x7 and x9 ) = '1' then
         y4 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s370;

      elsif ( not x65 and x66 and not x21 and not x22 and not x23 and x15 and not x7 and not x9 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and x66 and not x21 and not x22 and not x23 and not x15 and x7 and x9 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s320;

      elsif ( not x65 and x66 and not x21 and not x22 and not x23 and not x15 and x7 and not x9 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s333;

      elsif ( not x65 and x66 and not x21 and not x22 and not x23 and not x15 and not x7 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s320;

      elsif ( not x65 and not x66 and x24 and x26 and x18 and x15 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and not x66 and x24 and x26 and x18 and not x15 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and not x66 and x24 and x26 and x18 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x24 and x26 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x24 and not x26 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x65 and not x66 and not x24 and x25 and x26 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and not x24 and x25 and x26 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x66 and not x24 and x25 and x26 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s144;

      elsif ( not x65 and not x66 and not x24 and x25 and x26 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x24 and x25 and not x26 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x65 and not x66 and not x24 and not x25 and x26 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and not x66 and not x24 and not x25 and not x26 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x65 and not x66 and not x24 and not x25 and not x26 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x65 and not x66 and not x24 and not x25 and not x26 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s145 =>
      if ( x21 and x15 and x10 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s330;

      elsif ( x21 and x15 and not x10 and x12 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( x21 and x15 and not x10 and not x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s48;

      elsif ( x21 and not x15 and x16 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x21 and not x15 and not x16 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s340;

      elsif ( not x21 and x22 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s143;

      else
         current_group15m <= s1;

      end if;

   when s146 =>
      if ( x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s147 =>
      if ( x21 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x21 and x23 and x22 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x21 and x23 and not x22 and x20 and x14 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( not x21 and x23 and not x22 and x20 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( not x21 and x23 and not x22 and x20 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x23 and not x22 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x23 and x18 and x14 and x22 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( not x21 and not x23 and x18 and x14 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x21 and not x23 and x18 and not x14 and x13 and x22 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( not x21 and not x23 and x18 and not x14 and x13 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x21 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s148 =>
      if ( x20 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s302;

      elsif ( not x20 and x21 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      else
         current_group15m <= s1;

      end if;

   when s149 =>
      if ( x66 and x65 and x61 and x60 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and x65 and x61 and x60 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x66 and x65 and x61 and x60 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x66 and x65 and x61 and x60 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x66 and x65 and x61 and not x60 and x62 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x66 and x65 and x61 and not x60 and x62 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x66 and x65 and x61 and not x60 and x62 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and x61 and not x60 and x62 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x65 and x61 and not x60 and not x62 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and x65 and x61 and not x60 and not x62 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and x65 and x61 and not x60 and not x62 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x66 and x65 and x61 and not x60 and not x62 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x66 and x65 and not x61 and x60 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and x65 and not x61 and x60 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and x65 and not x61 and x60 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x66 and x65 and not x61 and x60 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x66 and x65 and not x61 and not x60 and x62 and x11 and x10 and x15 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and x65 and not x61 and not x60 and x62 and x11 and x10 and not x15 and x7 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and x65 and not x61 and not x60 and x62 and x11 and x10 and not x15 and not x7 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( x66 and x65 and not x61 and not x60 and x62 and x11 and not x10 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and x65 and not x61 and not x60 and x62 and not x11 and x12 and x9 and x15 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and x65 and not x61 and not x60 and x62 and not x11 and x12 and x9 and not x15 and x7 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and x65 and not x61 and not x60 and x62 and not x11 and x12 and x9 and not x15 and not x7 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( x66 and x65 and not x61 and not x60 and x62 and not x11 and x12 and not x9 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and x65 and not x61 and not x60 and x62 and not x11 and not x12 and x8 and x15 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and x65 and not x61 and not x60 and x62 and not x11 and not x12 and x8 and not x15 and x7 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and x65 and not x61 and not x60 and x62 and not x11 and not x12 and x8 and not x15 and not x7 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( x66 and x65 and not x61 and not x60 and x62 and not x11 and not x12 and not x8 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and x65 and not x61 and not x60 and not x62 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and not x65 and x67 and x62 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s159;

      elsif ( x66 and not x65 and x67 and not x62 and x63 and x17 and x13 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and not x65 and x67 and not x62 and x63 and x17 and x13 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( x66 and not x65 and x67 and not x62 and x63 and x17 and not x13 and x12 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and not x65 and x67 and not x62 and x63 and x17 and not x13 and x12 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( x66 and not x65 and x67 and not x62 and x63 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and x67 and not x62 and x63 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and x67 and not x62 and not x63 and x19 and x13 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x66 and not x65 and x67 and not x62 and not x63 and x19 and x13 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x66 and not x65 and x67 and not x62 and not x63 and x19 and not x13 and x12 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x66 and not x65 and x67 and not x62 and not x63 and x19 and not x13 and x12 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x66 and not x65 and x67 and not x62 and not x63 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and x67 and not x62 and not x63 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and x21 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x66 and not x65 and not x67 and x21 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x66 and not x65 and not x67 and x21 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and x23 and x22 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( x66 and not x65 and not x67 and not x21 and x23 and x22 and x17 and not x14 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( x66 and not x65 and not x67 and not x21 and x23 and x22 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and x23 and x22 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and x23 and not x22 and x19 and x14 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( x66 and not x65 and not x67 and not x21 and x23 and not x22 and x19 and not x14 and x13 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( x66 and not x65 and not x67 and not x21 and x23 and not x22 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and x23 and not x22 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and not x23 and x22 and x18 and x14 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and not x65 and not x67 and not x21 and not x23 and x22 and x18 and not x14 and x13 ) = '1' then
         current_group15m <= s40;

      elsif ( x66 and not x65 and not x67 and not x21 and not x23 and x22 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and not x23 and x22 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x65 and not x67 and not x21 and not x23 and not x22 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x66 and x65 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x66 and x65 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x65 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and x24 and x26 and x11 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s160;

      elsif ( not x66 and not x65 and x67 and x24 and x26 and not x11 and x18 and x15 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x66 and not x65 and x67 and x24 and x26 and not x11 and x18 and not x15 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x66 and not x65 and x67 and x24 and x26 and not x11 and x18 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and x24 and x26 and not x11 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and x24 and not x26 and x19 and x16 and x11 and x12 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s188;

      elsif ( not x66 and not x65 and x67 and x24 and not x26 and x19 and x16 and x11 and not x12 and x13 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s172;

      elsif ( not x66 and not x65 and x67 and x24 and not x26 and x19 and x16 and x11 and not x12 and not x13 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x66 and not x65 and x67 and x24 and not x26 and x19 and x16 and not x11 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s160;

      elsif ( not x66 and not x65 and x67 and x24 and not x26 and x19 and not x16 and x17 and x11 and x13 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      elsif ( not x66 and not x65 and x67 and x24 and not x26 and x19 and not x16 and x17 and x11 and not x13 ) = '1' then
         y15 <= '1' ;
         y112 <= '1' ;
         current_group15m <= s46;

      elsif ( not x66 and not x65 and x67 and x24 and not x26 and x19 and not x16 and x17 and not x11 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      elsif ( not x66 and not x65 and x67 and x24 and not x26 and x19 and not x16 and not x17 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and not x65 and x67 and x24 and not x26 and not x19 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x66 and not x65 and x67 and not x24 and x25 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x66 and not x65 and x67 and not x24 and x25 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x66 and not x65 and x67 and not x24 and x25 and x19 and not x14 and not x13 and x26 ) = '1' then
         current_group15m <= s149;

      elsif ( not x66 and not x65 and x67 and not x24 and x25 and x19 and not x14 and not x13 and not x26 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and not x24 and x25 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and x26 and x10 and x12 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and x26 and x10 and x12 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and x26 and x10 and x12 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and x26 and x10 and x12 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and x26 and x10 and not x12 ) = '1' then
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s165;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and x26 and not x10 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and x26 and not x10 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and x26 and not x10 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and x26 and not x10 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and not x26 and x10 and x12 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and not x26 and x10 and x12 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and not x26 and x10 and x12 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and not x26 and x10 and x12 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and not x26 and x10 and not x12 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and not x26 and not x10 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and not x26 and not x10 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and not x26 and not x10 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and x67 and not x24 and not x25 and not x26 and not x10 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x67 and x21 and x9 and x3 ) = '1' then
         current_group15m <= s40;

      elsif ( not x66 and not x65 and not x67 and x21 and x9 and not x3 and x4 ) = '1' then
         current_group15m <= s40;

      elsif ( not x66 and not x65 and not x67 and x21 and x9 and not x3 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x65 and not x67 and x21 and not x9 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s150 =>
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

   when s151 =>
      if ( x66 and x62 and x61 and x13 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x66 and x62 and x61 and not x13 and x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x66 and x62 and x61 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x62 and not x61 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x62 and x63 and x17 and x13 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and not x62 and x63 and x17 and x13 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( x66 and not x62 and x63 and x17 and not x13 and x12 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x66 and not x62 and x63 and x17 and not x13 and x12 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( x66 and not x62 and x63 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x62 and x63 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x62 and not x63 and x19 and x13 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x66 and not x62 and not x63 and x19 and x13 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x66 and not x62 and not x63 and x19 and not x13 and x12 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x66 and not x62 and not x63 and x19 and not x13 and x12 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x66 and not x62 and not x63 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x62 and not x63 and not x19 ) = '1' then
         current_group15m <= s1;

      else
         y2 <= '1' ;
         y6 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      end if;

   when s152 =>
      if ( x64 and x63 ) = '1' then
         y3 <= '1' ;
         y22 <= '1' ;
         y37 <= '1' ;
         current_group15m <= s397;

      elsif ( x64 and not x63 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s20;

      elsif ( not x64 and x63 ) = '1' then
         current_group15m <= s1;

      else
         y15 <= '1' ;
         current_group15m <= s149;

      end if;

   when s153 =>
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

   when s154 =>
      if ( x67 and x22 and x17 and x18 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x67 and x22 and x17 and not x18 and x19 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x67 and x22 and x17 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and x22 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x22 and x18 and x13 and x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x67 and not x22 and x18 and x13 and not x23 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x67 and not x22 and x18 and not x13 and x12 and x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x67 and not x22 and x18 and not x13 and x12 and not x23 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x67 and not x22 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x22 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x61 and x60 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( not x67 and x61 and not x60 and x62 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x67 and x61 and not x60 and x62 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x67 and x61 and not x60 and x62 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x61 and not x60 and x62 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x61 and not x60 and not x62 and x15 ) = '1' then
         current_group15m <= s73;

      elsif ( not x67 and x61 and not x60 and not x62 and not x15 and x16 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s291;

      elsif ( not x67 and x61 and not x60 and not x62 and not x15 and not x16 ) = '1' then
         current_group15m <= s73;

      elsif ( not x67 and not x61 and x60 and x15 ) = '1' then
         current_group15m <= s73;

      elsif ( not x67 and not x61 and x60 and not x15 and x16 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s291;

      elsif ( not x67 and not x61 and x60 and not x15 and not x16 ) = '1' then
         current_group15m <= s73;

      elsif ( not x67 and not x61 and not x60 and x62 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x61 and not x60 and not x62 and x15 and x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( not x67 and not x61 and not x60 and not x62 and x15 and not x7 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x67 and not x61 and not x60 and not x62 and x15 and not x7 and not x11 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s254;

      elsif ( not x67 and not x61 and not x60 and not x62 and not x15 and x16 and x4 ) = '1' then
         current_group15m <= s40;

      elsif ( not x67 and not x61 and not x60 and not x62 and not x15 and x16 and not x4 and x11 and x9 ) = '1' then
         current_group15m <= s40;

      elsif ( not x67 and not x61 and not x60 and not x62 and not x15 and x16 and not x4 and x11 and not x9 and x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( not x67 and not x61 and not x60 and not x62 and not x15 and x16 and not x4 and x11 and not x9 and not x7 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s118;

      elsif ( not x67 and not x61 and not x60 and not x62 and not x15 and x16 and not x4 and not x11 and x9 and x7 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( not x67 and not x61 and not x60 and not x62 and not x15 and x16 and not x4 and not x11 and x9 and not x7 and x10 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( not x67 and not x61 and not x60 and not x62 and not x15 and x16 and not x4 and not x11 and x9 and not x7 and not x10 ) = '1' then
         current_group15m <= s40;

      elsif ( not x67 and not x61 and not x60 and not x62 and not x15 and x16 and not x4 and not x11 and not x9 and x7 and x8 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( not x67 and not x61 and not x60 and not x62 and not x15 and x16 and not x4 and not x11 and not x9 and x7 and not x8 ) = '1' then
         current_group15m <= s40;

      elsif ( not x67 and not x61 and not x60 and not x62 and not x15 and x16 and not x4 and not x11 and not x9 and not x7 and x12 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( not x67 and not x61 and not x60 and not x62 and not x15 and x16 and not x4 and not x11 and not x9 and not x7 and not x12 ) = '1' then
         current_group15m <= s40;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      end if;

   when s155 =>
      if ( x65 and x60 and x61 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s252;

      elsif ( x65 and x60 and not x61 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x60 and not x61 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x60 and not x61 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x60 and not x61 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and not x60 and x62 and x61 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x65 and not x60 and x62 and not x61 ) = '1' then
         current_group15m <= s316;

      elsif ( x65 and not x60 and not x62 and x61 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x60 and not x62 and x61 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x60 and not x62 and x61 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and not x60 and not x62 and x61 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and not x60 and not x62 and not x61 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and x21 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x65 and x21 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x65 and x21 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and x23 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and not x21 and x22 and x23 and x17 and not x14 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and not x21 and x22 and x23 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and x23 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and not x23 and x18 and x14 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x21 and x22 and not x23 and x18 and not x14 and x13 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x21 and x22 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      else
         y4 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s180;

      end if;

   when s156 =>
      if ( x63 and x64 and x18 and x15 and x8 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( x63 and x64 and x18 and x15 and not x8 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x63 and x64 and x18 and not x15 and x16 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( x63 and x64 and x18 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s135;

      elsif ( x63 and x64 and not x18 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s152;

      elsif ( x63 and not x64 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s213;

      else
         y15 <= '1' ;
         current_group15m <= s149;

      end if;

   when s157 =>
      if ( x65 and x21 and x67 and x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x65 and x21 and x67 and x8 and not x9 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x65 and x21 and x67 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x21 and x67 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x21 and not x67 and x18 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x65 and x21 and not x67 and not x18 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x21 and not x67 and not x18 and x19 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x21 and not x67 and not x18 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x21 and not x67 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x23 and x22 and x67 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and x23 and x22 and x67 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and x23 and x22 and x67 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x23 and x22 and x67 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x23 and x22 and not x67 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( x65 and not x21 and x23 and x22 and not x67 and not x19 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x21 and x23 and x22 and not x67 and not x19 and x17 and not x14 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x21 and x23 and x22 and not x67 and not x19 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x23 and x22 and not x67 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x23 and not x22 and x67 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and x23 and not x22 and x67 and x9 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and x23 and not x22 and x67 and x9 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x23 and not x22 and x67 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x23 and not x22 and not x67 and x20 and x14 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x21 and x23 and not x22 and not x67 and x20 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x21 and x23 and not x22 and not x67 and x20 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x23 and not x22 and not x67 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x23 and x67 and x8 and x22 and x9 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and not x23 and x67 and x8 and x22 and not x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and not x23 and x67 and x8 and x22 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x23 and x67 and x8 and not x22 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and not x23 and x67 and x8 and not x22 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and not x23 and x67 and x8 and not x22 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x23 and x67 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x23 and not x67 and x18 and x14 and x22 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x21 and not x23 and not x67 and x18 and x14 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x21 and not x23 and not x67 and x18 and not x14 and x13 and x22 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x21 and not x23 and not x67 and x18 and not x14 and x13 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x21 and not x23 and not x67 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x23 and not x67 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x62 and x61 and x13 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and x62 and x61 and not x13 and x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and x62 and x61 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x62 and not x61 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x62 and x63 and x17 and x13 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and not x62 and x63 and x17 and x13 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x62 and x63 and x17 and not x13 and x12 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and not x62 and x63 and x17 and not x13 and x12 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x62 and x63 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x62 and x63 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x62 and not x63 and x19 and x13 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x62 and not x63 and x19 and x13 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and not x62 and not x63 and x19 and not x13 and x12 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x62 and not x63 and x19 and not x13 and x12 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and not x62 and not x63 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s158 =>
      if ( x65 and x21 and x18 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x65 and x21 and not x18 and x19 and x14 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x21 and not x18 and x19 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x21 and not x18 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x21 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x23 and x22 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( x65 and not x21 and x23 and x22 and not x19 and x17 and x14 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x21 and x23 and x22 and not x19 and x17 and not x14 and x13 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( x65 and not x21 and x23 and x22 and not x19 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x23 and x22 and not x19 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x23 and not x22 and x20 and x14 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x21 and x23 and not x22 and x20 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( x65 and not x21 and x23 and not x22 and x20 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x23 and not x22 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x23 and x18 and x14 and x22 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x21 and not x23 and x18 and x14 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x21 and not x23 and x18 and not x14 and x13 and x22 ) = '1' then
         y37 <= '1' ;
         current_group15m <= s120;

      elsif ( x65 and not x21 and not x23 and x18 and not x14 and x13 and not x22 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x21 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x62 and x61 and x13 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and x62 and x61 and not x13 and x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and x62 and x61 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x62 and not x61 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x62 and x63 and x17 and x13 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and not x62 and x63 and x17 and x13 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x62 and x63 and x17 and not x13 and x12 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and not x62 and x63 and x17 and not x13 and x12 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x62 and x63 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x62 and x63 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x62 and not x63 and x19 and x13 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x62 and not x63 and x19 and x13 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and not x62 and not x63 and x19 and not x13 and x12 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and not x62 and not x63 and x19 and not x13 and x12 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and not x62 and not x63 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s159 =>
      if ( x62 and x61 and x13 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x62 and x61 and not x13 and x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x62 and x61 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x62 and not x61 ) = '1' then
         current_group15m <= s1;

      else
         y15 <= '1' ;
         current_group15m <= s149;

      end if;

   when s160 =>
      if ( x24 and x26 and x18 and x15 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( x24 and x26 and x18 and not x15 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( x24 and x26 and x18 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x24 and x26 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x24 and not x26 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( x24 and not x26 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( x24 and not x26 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x24 and not x26 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x25 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x25 and x19 and not x14 and not x13 and x26 ) = '1' then
         current_group15m <= s160;

      elsif ( not x24 and x25 and x19 and not x14 and not x13 and not x26 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and x26 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x24 and not x25 and x26 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x24 and not x25 and x26 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and x26 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and not x26 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x24 and not x25 and not x26 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x24 and not x25 and not x26 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s161 =>
      if ( x65 and x21 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x65 and not x21 and x22 and x8 and x9 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and x22 and x8 and not x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and x22 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x22 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x22 and x23 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and not x22 and x23 and x9 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and not x22 and x23 and x9 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x22 and x23 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x22 and not x23 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and not x22 and not x23 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and not x22 and not x23 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x22 and not x23 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x24 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s160;

      elsif ( not x65 and not x24 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x24 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x65 and not x24 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s161;

      else
         current_group15m <= s1;

      end if;

   when s162 =>
      if ( x24 and x26 ) = '1' then
         current_group15m <= s1;

      elsif ( x24 and not x26 ) = '1' then
         y11 <= '1' ;
         y16 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s281;

      elsif ( not x24 and x25 and x15 and x10 and x11 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s160;

      elsif ( not x24 and x25 and x15 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s398;

      elsif ( not x24 and x25 and x15 and x10 and not x11 and not x12 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s160;

      elsif ( not x24 and x25 and x15 and not x10 and x12 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s399;

      elsif ( not x24 and x25 and x15 and not x10 and not x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s48;

      elsif ( not x24 and x25 and not x15 and x16 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( not x24 and x25 and not x15 and not x16 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      elsif ( not x24 and not x25 and x26 ) = '1' then
         y11 <= '1' ;
         y16 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s281;

      elsif ( not x24 and not x25 and not x26 and x18 and x15 and x12 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and not x25 and not x26 and x18 and x15 and not x12 and x11 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and not x25 and not x26 and x18 and x15 and not x12 and not x11 and x10 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x24 and not x25 and not x26 and x18 and x15 and not x12 and not x11 and not x10 ) = '1' then
         y12 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s49;

      elsif ( not x24 and not x25 and not x26 and x18 and not x15 and x16 and x10 and x12 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s282;

      elsif ( not x24 and not x25 and not x26 and x18 and not x15 and x16 and x10 and not x12 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s392;

      elsif ( not x24 and not x25 and not x26 and x18 and not x15 and x16 and not x10 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s282;

      elsif ( not x24 and not x25 and not x26 and x18 and not x15 and not x16 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      else
         y11 <= '1' ;
         y16 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s281;

      end if;

   when s163 =>
      if ( x65 ) = '1' then
         y15 <= '1' ;
         y21 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s313;

      elsif ( not x65 and x66 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      end if;

   when s164 =>
      if ( x24 and x26 and x18 and x15 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( x24 and x26 and x18 and not x15 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( x24 and x26 and x18 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x24 and x26 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x24 and not x26 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and x26 and x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and x26 and not x18 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x24 and x25 and not x26 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x25 and not x26 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x25 and not x26 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and not x26 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and x26 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x24 and not x25 and x26 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x24 and not x25 and x26 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and x26 and not x18 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s165 =>
      if ( x24 and x26 and x18 and x15 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( x24 and x26 and x18 and not x15 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( x24 and x26 and x18 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x24 and x26 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x24 and not x26 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x24 and x25 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x25 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x25 and x19 and not x14 and not x13 and x26 ) = '1' then
         current_group15m <= s165;

      elsif ( not x24 and x25 and x19 and not x14 and not x13 and not x26 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and x26 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x24 and not x25 and x26 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x24 and not x25 and x26 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and x26 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and not x26 and x5 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x24 and not x25 and not x26 and not x5 and x18 and x15 and x12 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and not x25 and not x26 and not x5 and x18 and x15 and not x12 and x11 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and not x25 and not x26 and not x5 and x18 and x15 and not x12 and not x11 and x10 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x24 and not x25 and not x26 and not x5 and x18 and x15 and not x12 and not x11 and not x10 ) = '1' then
         y12 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s49;

      elsif ( not x24 and not x25 and not x26 and not x5 and x18 and not x15 and x16 and x10 and x12 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s282;

      elsif ( not x24 and not x25 and not x26 and not x5 and x18 and not x15 and x16 and x10 and not x12 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s392;

      elsif ( not x24 and not x25 and not x26 and not x5 and x18 and not x15 and x16 and not x10 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s282;

      elsif ( not x24 and not x25 and not x26 and not x5 and x18 and not x15 and not x16 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      else
         y11 <= '1' ;
         y16 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s281;

      end if;

   when s166 =>
      if ( x24 and x26 and x11 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s160;

      elsif ( x24 and x26 and not x11 and x18 and x15 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( x24 and x26 and not x11 and x18 and not x15 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( x24 and x26 and not x11 and x18 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x24 and x26 and not x11 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x24 and not x26 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( x24 and not x26 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( x24 and not x26 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x24 and not x26 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x26 and x25 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x26 and x25 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x26 and x25 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s166;

      elsif ( not x24 and x26 and x25 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x26 and not x25 and x10 and x12 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x24 and x26 and not x25 and x10 and x12 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x24 and x26 and not x25 and x10 and x12 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x26 and not x25 and x10 and x12 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x26 and not x25 and x10 and not x12 ) = '1' then
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s165;

      elsif ( not x24 and x26 and not x25 and not x10 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x24 and x26 and not x25 and not x10 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x24 and x26 and not x25 and not x10 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x26 and not x25 and not x10 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x26 and x10 and x12 and x25 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and not x26 and x10 and x12 and x25 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and not x26 and x10 and x12 and x25 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x26 and x10 and x12 and x25 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x26 and x10 and x12 and not x25 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x24 and not x26 and x10 and x12 and not x25 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x24 and not x26 and x10 and x12 and not x25 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x26 and x10 and x12 and not x25 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x26 and x10 and not x12 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x24 and not x26 and not x10 and x25 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and not x26 and not x10 and x25 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and not x26 and not x10 and x25 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x26 and not x10 and x25 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x26 and not x10 and not x25 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x24 and not x26 and not x10 and not x25 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x24 and not x26 and not x10 and not x25 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s167 =>
      if ( x24 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s282;

      else
         y8 <= '1' ;
         y17 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s164;

      end if;

   when s168 =>
      if ( x66 and x42 and x15 and x8 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( x66 and x42 and x15 and not x8 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x66 and x42 and not x15 and x16 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s151;

      elsif ( x66 and x42 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s135;

      elsif ( x66 and not x42 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s400;

      elsif ( not x66 and x24 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x24 and x25 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      else
         y15 <= '1' ;
         current_group15m <= s149;

      end if;

   when s169 =>
      if ( x65 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x4 ) = '1' then
         current_group15m <= s1;

      else
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      end if;

   when s170 =>
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

   when s171 =>
      if ( x24 and x26 and x4 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( x24 and x26 and not x4 and x20 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( x24 and x26 and not x4 and not x20 and x21 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( x24 and x26 and not x4 and not x20 and not x21 and x22 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( x24 and x26 and not x4 and not x20 and not x21 and not x22 and x23 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( x24 and x26 and not x4 and not x20 and not x21 and not x22 and not x23 and x16 and x11 ) = '1' then
         y12 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s49;

      elsif ( x24 and x26 and not x4 and not x20 and not x21 and not x22 and not x23 and x16 and not x11 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x24 and x26 and not x4 and not x20 and not x21 and not x22 and not x23 and not x16 and x17 and x13 and x11 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x24 and x26 and not x4 and not x20 and not x21 and not x22 and not x23 and not x16 and x17 and x13 and not x11 and x12 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( x24 and x26 and not x4 and not x20 and not x21 and not x22 and not x23 and not x16 and x17 and x13 and not x11 and not x12 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x24 and x26 and not x4 and not x20 and not x21 and not x22 and not x23 and not x16 and x17 and not x13 and x11 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( x24 and x26 and not x4 and not x20 and not x21 and not x22 and not x23 and not x16 and x17 and not x13 and not x11 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x24 and x26 and not x4 and not x20 and not x21 and not x22 and not x23 and not x16 and not x17 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s51;

      elsif ( x24 and not x26 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( x24 and not x26 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( x24 and not x26 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x24 and not x26 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x25 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x25 and x19 and not x14 and not x13 and x26 ) = '1' then
         current_group15m <= s171;

      elsif ( not x24 and x25 and x19 and not x14 and not x13 and not x26 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and x26 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x24 and not x25 and x26 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x24 and not x25 and x26 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and x26 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and not x26 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x24 and not x25 and not x26 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x24 and not x25 and not x26 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s172 =>
      if ( x67 and x24 and x26 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x67 and x24 and not x26 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( x67 and not x24 and x25 and x26 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x67 and not x24 and x25 and not x26 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( x67 and not x24 and not x25 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x67 and x3 and x4 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( not x67 and x3 and not x4 and x5 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( not x67 and x3 and not x4 and not x5 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s173 =>
      if ( x67 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s355;

      else
         y2 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s105;

      end if;

   when s174 =>
      if ( x65 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x24 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x65 and not x24 and x15 and x10 and x11 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s187;

      elsif ( not x65 and not x24 and x15 and x10 and not x11 and x12 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s185;

      elsif ( not x65 and not x24 and x15 and x10 and not x11 and not x12 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s160;

      elsif ( not x65 and not x24 and x15 and not x10 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s50;

      elsif ( not x65 and not x24 and not x15 and x16 and x10 and x12 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s282;

      elsif ( not x65 and not x24 and not x15 and x16 and x10 and not x12 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and not x24 and not x15 and x16 and not x10 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s282;

      else
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      end if;

   when s175 =>
      if ( x24 and x26 ) = '1' then
         y11 <= '1' ;
         y16 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s281;

      elsif ( x24 and not x26 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( x24 and not x26 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( x24 and not x26 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x24 and not x26 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and x26 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x24 and not x25 and x26 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x24 and not x25 and x26 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and x26 and not x18 ) = '1' then
         current_group15m <= s1;

      else
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      end if;

   when s176 =>
      if ( x21 and x9 and x3 ) = '1' then
         current_group15m <= s40;

      elsif ( x21 and x9 and not x3 and x4 ) = '1' then
         current_group15m <= s40;

      elsif ( x21 and x9 and not x3 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x10 and x19 and x15 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s177;

      elsif ( not x21 and x22 and x10 and x19 and not x15 ) = '1' then
         y2 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      elsif ( not x21 and x22 and x10 and not x19 and x20 and x15 and x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s178;

      elsif ( not x21 and x22 and x10 and not x19 and x20 and x15 and not x14 and x16 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s178;

      elsif ( not x21 and x22 and x10 and not x19 and x20 and x15 and not x14 and not x16 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and x10 and not x19 and x20 and x15 and not x14 and not x16 and x5 and not x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and x10 and not x19 and x20 and x15 and not x14 and not x16 and x5 and not x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x10 and not x19 and x20 and x15 and not x14 and not x16 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x10 and not x19 and x20 and not x15 and x14 and x18 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s178;

      elsif ( not x21 and x22 and x10 and not x19 and x20 and not x15 and x14 and not x18 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and x10 and not x19 and x20 and not x15 and x14 and not x18 and x5 and not x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and x10 and not x19 and x20 and not x15 and x14 and not x18 and x5 and not x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x10 and not x19 and x20 and not x15 and x14 and not x18 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x10 and not x19 and x20 and not x15 and not x14 and x17 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s178;

      elsif ( not x21 and x22 and x10 and not x19 and x20 and not x15 and not x14 and not x17 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and x10 and not x19 and x20 and not x15 and not x14 and not x17 and x5 and not x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and x10 and not x19 and x20 and not x15 and not x14 and not x17 and x5 and not x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x10 and not x19 and x20 and not x15 and not x14 and not x17 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x10 and not x19 and not x20 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s151;

      elsif ( not x21 and x22 and not x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and x19 and x15 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x21 and not x22 and x19 and not x15 ) = '1' then
         y2 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      elsif ( not x21 and not x22 and not x19 and x20 ) = '1' then
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s179;

      else
         y21 <= '1' ;
         current_group15m <= s151;

      end if;

   when s177 =>
      if ( x21 and x9 and x3 ) = '1' then
         current_group15m <= s40;

      elsif ( x21 and x9 and not x3 and x4 ) = '1' then
         current_group15m <= s40;

      elsif ( x21 and x9 and not x3 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and x5 and not x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and x5 and not x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x19 and x15 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x21 and not x22 and x19 and not x15 ) = '1' then
         y2 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      else
         y21 <= '1' ;
         current_group15m <= s151;

      end if;

   when s178 =>
      if ( x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( x5 and not x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( x5 and not x4 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s179 =>
      if ( x21 and x6 ) = '1' then
         y8 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s106;

      elsif ( x21 and not x6 and x8 and x19 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( x21 and not x6 and x8 and not x19 and x20 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s176;

      elsif ( x21 and not x6 and x8 and not x19 and not x20 ) = '1' then
         y17 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s377;

      elsif ( x21 and not x6 and not x8 ) = '1' then
         y8 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s378;

      elsif ( not x21 and x22 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x4 and x5 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and not x22 and x4 and not x5 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and not x22 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s180 =>
      if ( x21 and x16 and x15 and x10 and x12 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( x21 and x16 and x15 and x10 and not x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( x21 and x16 and x15 and not x10 and x11 and x12 ) = '1' then
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s339;

      elsif ( x21 and x16 and x15 and not x10 and x11 and not x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s331;

      elsif ( x21 and x16 and x15 and not x10 and not x11 and x12 and x13 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s335;

      elsif ( x21 and x16 and x15 and not x10 and not x11 and x12 and not x13 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x16 and x15 and not x10 and not x11 and x12 and not x13 and x18 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x16 and x15 and not x10 and not x11 and x12 and not x13 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x16 and x15 and not x10 and not x11 and not x12 and x14 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s335;

      elsif ( x21 and x16 and x15 and not x10 and not x11 and not x12 and not x14 and x18 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x16 and x15 and not x10 and not x11 and not x12 and not x14 and x18 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x16 and x15 and not x10 and not x11 and not x12 and not x14 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x16 and not x15 and x12 and x10 and x8 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x16 and not x15 and x12 and x10 and x8 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x16 and not x15 and x12 and x10 and x8 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x16 and not x15 and x12 and x10 and x8 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x16 and not x15 and x12 and x10 and not x8 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( x21 and x16 and not x15 and x12 and x10 and not x8 and not x3 and x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( x21 and x16 and not x15 and x12 and x10 and not x8 and not x3 and not x5 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( x21 and x16 and not x15 and x12 and not x10 and x7 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( x21 and x16 and not x15 and x12 and not x10 and x7 and not x3 and x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( x21 and x16 and not x15 and x12 and not x10 and x7 and not x3 and not x5 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( x21 and x16 and not x15 and x12 and not x10 and not x7 and x11 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( x21 and x16 and not x15 and x12 and not x10 and not x7 and x11 and not x3 and x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( x21 and x16 and not x15 and x12 and not x10 and not x7 and x11 and not x3 and not x5 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( x21 and x16 and not x15 and x12 and not x10 and not x7 and not x11 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x16 and not x15 and x12 and not x10 and not x7 and not x11 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x16 and not x15 and x12 and not x10 and not x7 and not x11 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x16 and not x15 and x12 and not x10 and not x7 and not x11 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x16 and not x15 and not x12 and x10 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( x21 and x16 and not x15 and not x12 and x10 and not x3 and x5 ) = '1' then
         y4 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s315;

      elsif ( x21 and x16 and not x15 and not x12 and x10 and not x3 and not x5 ) = '1' then
         y4 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s370;

      elsif ( x21 and x16 and not x15 and not x12 and not x10 and x11 and x9 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( x21 and x16 and not x15 and not x12 and not x10 and x11 and x9 and not x3 and x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( x21 and x16 and not x15 and not x12 and not x10 and x11 and x9 and not x3 and not x5 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( x21 and x16 and not x15 and not x12 and not x10 and x11 and not x9 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x16 and not x15 and not x12 and not x10 and x11 and not x9 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x16 and not x15 and not x12 and not x10 and x11 and not x9 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x16 and not x15 and not x12 and not x10 and x11 and not x9 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x16 and not x15 and not x12 and not x10 and not x11 and x8 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( x21 and x16 and not x15 and not x12 and not x10 and not x11 and x8 and not x3 and x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( x21 and x16 and not x15 and not x12 and not x10 and not x11 and x8 and not x3 and not x5 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( x21 and x16 and not x15 and not x12 and not x10 and not x11 and not x8 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x16 and not x15 and not x12 and not x10 and not x11 and not x8 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x16 and not x15 and not x12 and not x10 and not x11 and not x8 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x16 and not x15 and not x12 and not x10 and not x11 and not x8 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x16 and x15 and x10 and x11 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( x21 and not x16 and x15 and x10 and not x11 and x12 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s126;

      elsif ( x21 and not x16 and x15 and x10 and not x11 and not x12 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( x21 and not x16 and x15 and x10 and not x11 and not x12 and not x3 and x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( x21 and not x16 and x15 and x10 and not x11 and not x12 and not x3 and not x5 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( x21 and not x16 and x15 and not x10 and x11 and x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s285;

      elsif ( x21 and not x16 and x15 and not x10 and x11 and not x12 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x21 and not x16 and x15 and not x10 and not x11 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( x21 and not x16 and x15 and not x10 and not x11 and not x3 and x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( x21 and not x16 and x15 and not x10 and not x11 and not x3 and not x5 and x12 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s333;

      elsif ( x21 and not x16 and x15 and not x10 and not x11 and not x3 and not x5 and not x12 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s332;

      elsif ( x21 and not x16 and not x15 and x3 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s163;

      elsif ( x21 and not x16 and not x15 and not x3 and x5 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( x21 and not x16 and not x15 and not x3 and not x5 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s5;

      elsif ( not x21 and x22 and x23 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x21 and x22 and not x23 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x21 and not x22 and x23 and x19 and x14 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x21 and not x22 and x23 and x19 and not x14 and x13 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x21 and not x22 and x23 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x23 and x18 and x14 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x21 and not x22 and not x23 and x18 and not x14 and x13 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x21 and not x22 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s181 =>
         y8 <= '1' ;
         current_group15m <= s92;

   when s182 =>
      if ( x68 and x20 and x18 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x68 and x20 and x18 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x68 and x20 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x68 and x20 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x68 and not x20 and x21 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( x68 and not x20 and not x21 and x17 and x13 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( x68 and not x20 and not x21 and x17 and not x13 and x12 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( x68 and not x20 and not x21 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x68 and not x20 and not x21 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x68 and x24 and x26 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x68 and x24 and not x26 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x68 and x24 and not x26 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x68 and x24 and not x26 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x68 and x24 and not x26 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x68 and not x24 and x25 and x26 and x15 and x10 and x11 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s160;

      elsif ( not x68 and not x24 and x25 and x26 and x15 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s398;

      elsif ( not x68 and not x24 and x25 and x26 and x15 and x10 and not x11 and not x12 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s160;

      elsif ( not x68 and not x24 and x25 and x26 and x15 and not x10 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s399;

      elsif ( not x68 and not x24 and x25 and x26 and not x15 and x16 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s282;

      elsif ( not x68 and not x24 and x25 and x26 and not x15 and not x16 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      elsif ( not x68 and not x24 and x25 and not x26 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x68 and not x24 and not x25 and x26 and x19 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x68 and not x24 and not x25 and x26 and not x19 and x20 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x68 and not x24 and not x25 and x26 and not x19 and not x20 and x21 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x68 and not x24 and not x25 and x26 and not x19 and not x20 and not x21 and x22 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x68 and not x24 and not x25 and x26 and not x19 and not x20 and not x21 and not x22 and x16 and x11 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x68 and not x24 and not x25 and x26 and not x19 and not x20 and not x21 and not x22 and x16 and not x11 and x12 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x68 and not x24 and not x25 and x26 and not x19 and not x20 and not x21 and not x22 and x16 and not x11 and not x12 and x10 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x68 and not x24 and not x25 and x26 and not x19 and not x20 and not x21 and not x22 and x16 and not x11 and not x12 and not x10 ) = '1' then
         y12 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s49;

      elsif ( not x68 and not x24 and not x25 and x26 and not x19 and not x20 and not x21 and not x22 and not x16 and x17 and x10 and x12 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( not x68 and not x24 and not x25 and x26 and not x19 and not x20 and not x21 and not x22 and not x16 and x17 and x10 and not x12 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x68 and not x24 and not x25 and x26 and not x19 and not x20 and not x21 and not x22 and not x16 and x17 and not x10 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( not x68 and not x24 and not x25 and x26 and not x19 and not x20 and not x21 and not x22 and not x16 and not x17 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x68 and not x24 and not x25 and not x26 and x15 and x12 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x68 and not x24 and not x25 and not x26 and x15 and not x12 and x11 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x68 and not x24 and not x25 and not x26 and x15 and not x12 and not x11 and x10 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x68 and not x24 and not x25 and not x26 and x15 and not x12 and not x11 and not x10 ) = '1' then
         y12 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s49;

      elsif ( not x68 and not x24 and not x25 and not x26 and not x15 and x16 and x10 and x12 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s282;

      elsif ( not x68 and not x24 and not x25 and not x26 and not x15 and x16 and x10 and not x12 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s392;

      elsif ( not x68 and not x24 and not x25 and not x26 and not x15 and x16 and not x10 ) = '1' then
         y5 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s282;

      else
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      end if;

   when s183 =>
      if ( x24 and x4 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( x24 and not x4 and x20 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( x24 and not x4 and not x20 and x21 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( x24 and not x4 and not x20 and not x21 and x22 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( x24 and not x4 and not x20 and not x21 and not x22 and x23 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( x24 and not x4 and not x20 and not x21 and not x22 and not x23 and x16 and x11 ) = '1' then
         y12 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s49;

      elsif ( x24 and not x4 and not x20 and not x21 and not x22 and not x23 and x16 and not x11 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x24 and not x4 and not x20 and not x21 and not x22 and not x23 and not x16 and x17 and x13 and x11 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x24 and not x4 and not x20 and not x21 and not x22 and not x23 and not x16 and x17 and x13 and not x11 and x12 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( x24 and not x4 and not x20 and not x21 and not x22 and not x23 and not x16 and x17 and x13 and not x11 and not x12 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x24 and not x4 and not x20 and not x21 and not x22 and not x23 and not x16 and x17 and not x13 and x11 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( x24 and not x4 and not x20 and not x21 and not x22 and not x23 and not x16 and x17 and not x13 and not x11 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( x24 and not x4 and not x20 and not x21 and not x22 and not x23 and not x16 and not x17 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s51;

      elsif ( not x24 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s183;

      else
         current_group15m <= s1;

      end if;

   when s184 =>
         y11 <= '1' ;
         current_group15m <= s53;

   when s185 =>
      if ( x26 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s48;

      else
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      end if;

   when s186 =>
      if ( x68 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s401;

      elsif ( not x68 and x26 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      else
         y15 <= '1' ;
         y112 <= '1' ;
         current_group15m <= s46;

      end if;

   when s187 =>
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

   when s188 =>
      if ( x66 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x66 and x24 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x66 and not x24 and x26 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      else
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      end if;

   when s189 =>
      if ( x65 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      else
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s402;

      end if;

   when s190 =>
      if ( x66 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      else
         y5 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s167;

      end if;

   when s191 =>
      if ( x65 and x66 and x68 and x21 and x20 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s403;

      elsif ( x65 and x66 and x68 and x21 and not x20 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( x65 and x66 and x68 and not x21 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( x65 and x66 and not x68 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      elsif ( x65 and not x66 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( not x65 and x16 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      else
         y12 <= '1' ;
         current_group15m <= s100;

      end if;

   when s192 =>
      if ( x21 and x20 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x20 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x20 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x20 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x20 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x20 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x20 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x20 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x19 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x21 and x19 and not x14 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x21 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s193 =>
      if ( x21 and x20 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x20 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x20 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x20 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x20 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x20 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x20 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x20 and not x19 ) = '1' then
         current_group15m <= s1;

      else
         y10 <= '1' ;
         current_group15m <= s12;

      end if;

   when s194 =>
      if ( x21 and x20 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x20 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x20 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x20 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x20 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x21 and x19 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x21 and x19 and not x14 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x21 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s195 =>
      if ( x21 and x20 ) = '1' then
         y1 <= '1' ;
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s194;

      elsif ( x21 and not x20 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x20 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x20 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x20 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x19 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x21 and x19 and not x14 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x21 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s196 =>
      if ( x21 and x20 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x20 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x20 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x20 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x20 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      else
         y10 <= '1' ;
         current_group15m <= s12;

      end if;

   when s197 =>
      if ( x21 and x65 and x20 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x65 and x20 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x65 and x20 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x65 and x20 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x65 and not x20 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x21 and not x65 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and not x65 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and not x65 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x65 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x65 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x65 and x22 and x23 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x21 and not x65 and x22 and x23 and x17 and not x14 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x21 and not x65 and x22 and x23 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x65 and x22 and x23 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x65 and x22 and not x23 and x18 and x14 ) = '1' then
         current_group15m <= s40;

      elsif ( not x21 and not x65 and x22 and not x23 and x18 and not x14 and x13 ) = '1' then
         current_group15m <= s40;

      elsif ( not x21 and not x65 and x22 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x65 and x22 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x65 and not x22 and x23 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s180;

      else
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s404;

      end if;

   when s198 =>
      if ( x65 and x21 and x20 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x21 and x20 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x21 and x20 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x21 and x20 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x21 and not x20 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x21 and not x20 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x21 and not x20 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x21 and not x20 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x19 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x21 and x19 and not x14 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and not x21 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x20 and x18 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x20 and x18 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x20 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x20 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x20 and x21 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x20 and x21 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x20 and x21 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x20 and x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x20 and not x21 and x17 and x13 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x65 and not x20 and not x21 and x17 and not x13 and x12 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x65 and not x20 and not x21 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s199 =>
      if ( x21 and x20 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x20 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x20 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x20 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x20 and x10 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s302;

      elsif ( x21 and not x20 and not x10 and x11 and x12 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x20 and not x10 and x11 and x12 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x20 and not x10 and x11 and x12 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x20 and not x10 and x11 and x12 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x20 and not x10 and x11 and not x12 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s302;

      elsif ( x21 and not x20 and not x10 and not x11 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s302;

      elsif ( not x21 and x19 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x21 and x19 and not x14 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x21 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s200 =>
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s405;

   when s201 =>
      if ( x20 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x20 and x21 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      else
         y10 <= '1' ;
         current_group15m <= s12;

      end if;

   when s202 =>
      if ( x10 and x12 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s259;

      elsif ( x10 and not x12 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      else
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s259;

      end if;

   when s203 =>
      if ( x65 and x21 and x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x65 and x21 and x8 and not x9 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x65 and x21 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x21 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x23 and x22 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and x23 and x22 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and x23 and x22 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x23 and x22 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x23 and not x22 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and x23 and not x22 and x9 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and x23 and not x22 and x9 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and x23 and not x22 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x23 and x8 and x22 and x9 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and not x23 and x8 and x22 and not x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and not x23 and x8 and x22 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x23 and x8 and not x22 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and not x23 and x8 and not x22 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x21 and not x23 and x8 and not x22 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 and not x23 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x62 and x61 and x13 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and x66 and x62 and x61 and not x13 and x12 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and x66 and x62 and x61 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and x62 and not x61 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x62 and x63 and x17 and x13 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and x66 and not x62 and x63 and x17 and x13 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and x66 and not x62 and x63 and x17 and not x13 and x12 and x64 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x65 and x66 and not x62 and x63 and x17 and not x13 and x12 and not x64 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and x66 and not x62 and x63 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x62 and x63 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x62 and not x63 and x19 and x13 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x66 and not x62 and not x63 and x19 and x13 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x66 and not x62 and not x63 and x19 and not x13 and x12 and x64 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x65 and x66 and not x62 and not x63 and x19 and not x13 and x12 and not x64 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x66 and not x62 and not x63 and x19 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x62 and not x63 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x21 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      else
         y5 <= '1' ;
         current_group15m <= s101;

      end if;

   when s204 =>
         y15 <= '1' ;
         current_group15m <= s149;

   when s205 =>
      if ( x21 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x21 and x22 and x23 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x21 and x22 and not x23 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s147;

      else
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s147;

      end if;

   when s206 =>
      if ( x20 and x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x20 and not x15 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s59;

      elsif ( not x20 and x21 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x20 and x21 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x20 and x21 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x20 and x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x20 and not x21 and x17 and x13 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x20 and not x21 and x17 and not x13 and x12 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x20 and not x21 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s207 =>
      if ( x20 and x18 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x20 and x18 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x20 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x20 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x20 and x21 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x20 and x21 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x20 and x21 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x20 and x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x20 and not x21 and x17 and x13 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x20 and not x21 and x17 and not x13 and x12 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x20 and not x21 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s208 =>
      if ( x1 ) = '1' then
         y2 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s277;

      elsif ( not x1 and x17 and x15 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s198;

      elsif ( not x1 and x17 and not x15 and x16 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s59;

      elsif ( not x1 and x17 and not x15 and not x16 ) = '1' then
         y7 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s211;

      else
         y12 <= '1' ;
         y15 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s401;

      end if;

   when s209 =>
      if ( x20 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s393;

      else
         y2 <= '1' ;
         current_group15m <= s56;

      end if;

   when s210 =>
      if ( x65 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( not x65 and x66 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x66 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x66 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x66 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and x20 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s393;

      elsif ( not x65 and not x66 and not x20 and x21 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x66 and not x20 and x21 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x66 and not x20 and x21 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x20 and x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x66 and not x20 and not x21 and x17 and x13 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x65 and not x66 and not x20 and not x21 and x17 and not x13 and x12 ) = '1' then
         y1 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s148;

      elsif ( not x65 and not x66 and not x20 and not x21 and x17 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s211 =>
      if ( x66 and x21 and x19 and x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and x21 and x19 and not x15 and x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and x21 and x19 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x21 and x20 and x15 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x66 and not x21 and x20 and not x15 and x14 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x66 and not x21 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x21 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x20 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s393;

      elsif ( not x66 and not x20 and x21 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x66 and not x20 and x21 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x66 and not x20 and x21 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x20 and x21 and not x18 ) = '1' then
         current_group15m <= s1;

      else
         y2 <= '1' ;
         current_group15m <= s56;

      end if;

   when s212 =>
      if ( x21 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x21 and x22 and x23 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x21 and x22 and not x23 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s147;

      elsif ( not x21 and not x22 and x23 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s147;

      elsif ( not x21 and not x22 and not x23 and x18 and x14 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x21 and not x22 and not x23 and x18 and not x14 and x13 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( not x21 and not x22 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s213 =>
      if ( x64 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      else
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s152;

      end if;

   when s214 =>
      if ( x21 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      else
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s308;

      end if;

   when s215 =>
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

   when s216 =>
      if ( x21 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x21 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x21 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x21 and not x22 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x21 and not x22 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x21 and not x22 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s217 =>
      if ( x21 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x21 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x21 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x7 and x8 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x21 and x22 and x7 and not x8 and x9 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x21 and x22 and x7 and not x8 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x21 and not x22 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x21 and not x22 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s218 =>
      if ( x21 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x21 and x22 and x10 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s219;

      elsif ( not x21 and x22 and not x10 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s28;

      elsif ( not x21 and not x22 and x8 and x16 and x15 and x10 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s219;

      elsif ( not x21 and not x22 and x8 and x16 and x15 and not x10 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s309;

      elsif ( not x21 and not x22 and x8 and x16 and not x15 and x10 ) = '1' then
         y2 <= '1' ;
         y16 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s124;

      elsif ( not x21 and not x22 and x8 and x16 and not x15 and not x10 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s310;

      elsif ( not x21 and not x22 and x8 and not x16 and x17 and x10 and x15 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s219;

      elsif ( not x21 and not x22 and x8 and not x16 and x17 and x10 and not x15 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s308;

      elsif ( not x21 and not x22 and x8 and not x16 and x17 and not x10 ) = '1' then
         y2 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s79;

      elsif ( not x21 and not x22 and x8 and not x16 and not x17 and x10 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s219;

      elsif ( not x21 and not x22 and x8 and not x16 and not x17 and not x10 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s311;

      else
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      end if;

   when s219 =>
         y17 <= '1' ;
         current_group15m <= s77;

   when s220 =>
      if ( x21 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s311;

      elsif ( not x21 and x22 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x21 and not x22 and x3 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s218;

      elsif ( not x21 and not x22 and not x3 and x8 and x16 and x15 and x10 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s219;

      elsif ( not x21 and not x22 and not x3 and x8 and x16 and x15 and not x10 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s309;

      elsif ( not x21 and not x22 and not x3 and x8 and x16 and not x15 and x10 ) = '1' then
         y2 <= '1' ;
         y16 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s124;

      elsif ( not x21 and not x22 and not x3 and x8 and x16 and not x15 and not x10 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s310;

      elsif ( not x21 and not x22 and not x3 and x8 and not x16 and x17 and x10 and x15 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s219;

      elsif ( not x21 and not x22 and not x3 and x8 and not x16 and x17 and x10 and not x15 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s308;

      elsif ( not x21 and not x22 and not x3 and x8 and not x16 and x17 and not x10 ) = '1' then
         y2 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s79;

      elsif ( not x21 and not x22 and not x3 and x8 and not x16 and not x17 and x10 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s219;

      elsif ( not x21 and not x22 and not x3 and x8 and not x16 and not x17 and not x10 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s311;

      else
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      end if;

   when s221 =>
      if ( x21 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x21 and x22 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      else
         y2 <= '1' ;
         y16 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s124;

      end if;

   when s222 =>
         y17 <= '1' ;
         current_group15m <= s17;

   when s223 =>
      if ( x21 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s161;

      elsif ( not x21 and x22 and x8 and x9 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x8 and not x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x12 and x23 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s247;

      elsif ( not x21 and not x22 and x12 and not x23 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x21 and not x22 and not x12 and x23 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and not x12 and x23 and x9 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and not x12 and x23 and x9 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x12 and x23 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x12 and not x23 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and not x12 and not x23 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and not x12 and not x23 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s224 =>
      if ( x66 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      else
         y22 <= '1' ;
         current_group15m <= s4;

      end if;

   when s225 =>
         y2 <= '1' ;
         y6 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

   when s226 =>
      if ( x21 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x21 and x22 and x17 and x10 and x15 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s283;

      elsif ( not x21 and x22 and x17 and x10 and not x15 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( not x21 and x22 and x17 and not x10 ) = '1' then
         y13 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s284;

      elsif ( not x21 and x22 and not x17 and x10 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s219;

      elsif ( not x21 and x22 and not x17 and not x10 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s217;

      elsif ( not x21 and not x22 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x21 and not x22 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x21 and not x22 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s227 =>
      if ( x21 and x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and x8 and not x9 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x23 and x22 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x23 and x22 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x23 and x22 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x23 and x22 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x23 and not x22 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x23 and not x22 and x9 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x23 and not x22 and x9 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x23 and not x22 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x23 and x8 and x22 and x9 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x23 and x8 and x22 and not x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x23 and x8 and x22 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x23 and x8 and not x22 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x23 and x8 and not x22 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x23 and x8 and not x22 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s228 =>
      if ( x21 and x18 ) = '1' then
         y14 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s116;

      elsif ( x21 and not x18 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s117;

      elsif ( not x21 and x22 and x23 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x21 and x22 and x23 and not x12 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x23 and not x12 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x23 and not x12 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and not x12 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s243;

      else
         y14 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s116;

      end if;

   when s229 =>
      if ( x21 and x18 and x4 and x15 and x17 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x21 and x18 and x4 and x15 and not x17 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s231;

      elsif ( x21 and x18 and x4 and not x15 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s235;

      elsif ( x21 and x18 and not x4 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s231;

      elsif ( x21 and not x18 and x19 and x15 and x4 and x17 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x21 and not x18 and x19 and x15 and x4 and not x17 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s231;

      elsif ( x21 and not x18 and x19 and x15 and not x4 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s231;

      elsif ( x21 and not x18 and x19 and not x15 and x16 and x14 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s231;

      elsif ( x21 and not x18 and x19 and not x15 and x16 and not x14 and x17 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s231;

      elsif ( x21 and not x18 and x19 and not x15 and x16 and not x14 and not x17 and x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and not x18 and x19 and not x15 and x16 and not x14 and not x17 and x8 and not x9 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and not x18 and x19 and not x15 and x16 and not x14 and not x17 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 and x19 and not x15 and x16 and not x14 and not x17 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 and x19 and not x15 and not x16 and x17 and x12 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s231;

      elsif ( x21 and not x18 and x19 and not x15 and not x16 and x17 and not x12 and x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and not x18 and x19 and not x15 and not x16 and x17 and not x12 and x8 and not x9 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and not x18 and x19 and not x15 and not x16 and x17 and not x12 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 and x19 and not x15 and not x16 and x17 and not x12 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 and x19 and not x15 and not x16 and not x17 and x13 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s231;

      elsif ( x21 and not x18 and x19 and not x15 and not x16 and not x17 and not x13 and x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and not x18 and x19 and not x15 and not x16 and not x17 and not x13 and x8 and not x9 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and not x18 and x19 and not x15 and not x16 and not x17 and not x13 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 and x19 and not x15 and not x16 and not x17 and not x13 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 and not x19 and x4 ) = '1' then
         y15 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s36;

      elsif ( x21 and not x18 and not x19 and not x4 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s231;

      elsif ( not x21 and x23 and x22 and x6 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s231;

      elsif ( not x21 and x23 and x22 and not x6 and x7 and x18 and x15 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( not x21 and x23 and x22 and not x6 and x7 and x18 and not x15 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x21 and x23 and x22 and not x6 and x7 and not x18 and x19 and x15 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s247;

      elsif ( not x21 and x23 and x22 and not x6 and x7 and not x18 and x19 and not x15 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      elsif ( not x21 and x23 and x22 and not x6 and x7 and not x18 and not x19 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s33;

      elsif ( not x21 and x23 and x22 and not x6 and not x7 ) = '1' then
         y3 <= '1' ;
         y12 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s34;

      elsif ( not x21 and x23 and not x22 ) = '1' then
         y12 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s230;

      elsif ( not x21 and not x23 and x22 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s161;

      elsif ( not x21 and not x23 and not x22 and x6 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s231;

      elsif ( not x21 and not x23 and not x22 and not x6 and x7 and x18 and x15 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( not x21 and not x23 and not x22 and not x6 and x7 and x18 and not x15 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x21 and not x23 and not x22 and not x6 and x7 and not x18 and x19 and x15 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s247;

      elsif ( not x21 and not x23 and not x22 and not x6 and x7 and not x18 and x19 and not x15 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      elsif ( not x21 and not x23 and not x22 and not x6 and x7 and not x18 and not x19 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s33;

      else
         y3 <= '1' ;
         y12 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s34;

      end if;

   when s230 =>
      if ( x21 and x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and x8 and not x9 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x18 and x15 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( not x21 and x22 and x18 and not x15 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x21 and x22 and not x18 and x19 and x15 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x21 and x22 and not x18 and x19 and not x15 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x21 and x22 and not x18 and not x19 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( not x21 and not x22 and x23 and x19 and x16 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( not x21 and not x22 and x23 and x19 and not x16 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and x16 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s228;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x21 and not x22 and x23 and not x19 and not x20 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s231;

      elsif ( not x21 and not x22 and not x23 and x18 and x15 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( not x21 and not x22 and not x23 and x18 and not x15 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x21 and not x22 and not x23 and not x18 and x19 and x15 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s247;

      elsif ( not x21 and not x22 and not x23 and not x18 and x19 and not x15 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      else
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s33;

      end if;

   when s231 =>
      if ( x65 and x66 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and not x66 and x21 and x5 ) = '1' then
         y3 <= '1' ;
         y12 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s34;

      elsif ( x65 and not x66 and x21 and not x5 and x6 and x18 and x15 and x17 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and not x66 and x21 and not x5 and x6 and x18 and x15 and not x17 ) = '1' then
         y2 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s244;

      elsif ( x65 and not x66 and x21 and not x5 and x6 and x18 and not x15 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x65 and not x66 and x21 and not x5 and x6 and not x18 and x19 and x15 and x17 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and not x66 and x21 and not x5 and x6 and not x18 and x19 and x15 and not x17 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s246;

      elsif ( x65 and not x66 and x21 and not x5 and x6 and not x18 and x19 and not x15 ) = '1' then
         y8 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s227;

      elsif ( x65 and not x66 and x21 and not x5 and x6 and not x18 and not x19 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s31;

      elsif ( x65 and not x66 and x21 and not x5 and not x6 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s247;

      elsif ( x65 and not x66 and not x21 and x22 and x23 and x7 and x18 and x15 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( x65 and not x66 and not x21 and x22 and x23 and x7 and x18 and not x15 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x65 and not x66 and not x21 and x22 and x23 and x7 and not x18 and x19 and x15 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s247;

      elsif ( x65 and not x66 and not x21 and x22 and x23 and x7 and not x18 and x19 and not x15 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      elsif ( x65 and not x66 and not x21 and x22 and x23 and x7 and not x18 and not x19 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s33;

      elsif ( x65 and not x66 and not x21 and x22 and x23 and not x7 ) = '1' then
         y3 <= '1' ;
         y12 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s34;

      elsif ( x65 and not x66 and not x21 and x22 and not x23 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s161;

      elsif ( x65 and not x66 and not x21 and not x22 and x23 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s161;

      elsif ( x65 and not x66 and not x21 and not x22 and not x23 and x7 and x18 and x15 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( x65 and not x66 and not x21 and not x22 and not x23 and x7 and x18 and not x15 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( x65 and not x66 and not x21 and not x22 and not x23 and x7 and not x18 and x19 and x15 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s247;

      elsif ( x65 and not x66 and not x21 and not x22 and not x23 and x7 and not x18 and x19 and not x15 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      elsif ( x65 and not x66 and not x21 and not x22 and not x23 and x7 and not x18 and not x19 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s33;

      elsif ( x65 and not x66 and not x21 and not x22 and not x23 and not x7 ) = '1' then
         y3 <= '1' ;
         y12 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s34;

      else
         y17 <= '1' ;
         current_group15m <= s77;

      end if;

   when s232 =>
      if ( x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      else
         y2 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s322;

      end if;

   when s233 =>
      if ( x21 and x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and x8 and not x9 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x23 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x23 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s161;

      else
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s161;

      end if;

   when s234 =>
      if ( x21 and x65 and x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and x65 and x8 and not x9 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and x65 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x65 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x65 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( not x21 and x65 and x23 and x22 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x65 and x23 and x22 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x65 and x23 and x22 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x65 and x23 and x22 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x65 and x23 and not x22 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x65 and x23 and not x22 and x9 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x65 and x23 and not x22 and x9 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x65 and x23 and not x22 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x65 and not x23 and x8 and x22 and x9 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x65 and not x23 and x8 and x22 and not x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x65 and not x23 and x8 and x22 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x65 and not x23 and x8 and not x22 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x65 and not x23 and x8 and not x22 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x65 and not x23 and x8 and not x22 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x65 and not x23 and not x8 ) = '1' then
         current_group15m <= s1;

      else
         y5 <= '1' ;
         current_group15m <= s101;

      end if;

   when s235 =>
      if ( x21 and x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and x8 and not x9 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x23 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x23 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s161;

      elsif ( not x21 and not x22 and x23 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s161;

      elsif ( not x21 and not x22 and not x23 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and not x23 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and not x23 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s236 =>
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s28;

   when s237 =>
      if ( x21 and x18 and x15 and x17 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and x18 and x15 and not x17 ) = '1' then
         y2 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s244;

      elsif ( x21 and x18 and not x15 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x21 and not x18 and x19 and x15 and x17 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x18 and x19 and x15 and not x17 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s246;

      elsif ( x21 and not x18 and x19 and not x15 ) = '1' then
         y24 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s157;

      elsif ( x21 and not x18 and not x19 ) = '1' then
         y1 <= '1' ;
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s31;

      elsif ( not x21 and x22 and x23 and x18 and x15 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( not x21 and x22 and x23 and x18 and not x15 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x21 and x22 and x23 and not x18 and x19 and x15 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s247;

      elsif ( not x21 and x22 and x23 and not x18 and x19 and not x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x21 and x22 and x23 and not x18 and not x19 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s33;

      elsif ( not x21 and x22 and not x23 ) = '1' then
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s161;

      elsif ( not x21 and not x22 and x23 and x19 and x16 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( not x21 and not x22 and x23 and x19 and not x16 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and x16 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s228;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and x18 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and not x18 and x17 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and not x18 and not x17 and x5 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s283;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and not x18 and not x17 and not x5 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      elsif ( not x21 and not x22 and x23 and not x19 and not x20 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s231;

      elsif ( not x21 and not x22 and not x23 and x18 and x15 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( not x21 and not x22 and not x23 and x18 and not x15 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x21 and not x22 and not x23 and not x18 and x19 and x15 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s247;

      elsif ( not x21 and not x22 and not x23 and not x18 and x19 and not x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      else
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s33;

      end if;

   when s238 =>
      if ( x21 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s33;

      elsif ( not x21 and x22 and x23 and x15 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s240;

      elsif ( not x21 and x22 and x23 and not x15 and x19 and x18 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s240;

      elsif ( not x21 and x22 and x23 and not x15 and x19 and not x18 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x23 and not x15 and x19 and not x18 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x23 and not x15 and x19 and not x18 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and not x15 and x19 and not x18 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and not x15 and not x19 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s240;

      elsif ( not x21 and x22 and not x23 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x23 and x15 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s240;

      elsif ( not x21 and not x22 and not x23 and not x15 and x19 and x18 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s240;

      elsif ( not x21 and not x22 and not x23 and not x15 and x19 and not x18 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and not x23 and not x15 and x19 and not x18 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and not x23 and not x15 and x19 and not x18 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x23 and not x15 and x19 and not x18 and not x8 ) = '1' then
         current_group15m <= s1;

      else
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s240;

      end if;

   when s239 =>
      if ( x26 ) = '1' then
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s165;

      else
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s25;

      end if;

   when s240 =>
      if ( x21 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x21 and x22 and x23 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 and x6 and x18 and x15 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( not x21 and x22 and not x23 and x6 and x18 and not x15 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x21 and x22 and not x23 and x6 and not x18 and x19 and x15 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x21 and x22 and not x23 and x6 and not x18 and x19 and not x15 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x21 and x22 and not x23 and x6 and not x18 and not x19 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s229;

      elsif ( not x21 and x22 and not x23 and not x6 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s28;

      elsif ( not x21 and not x22 and x23 and x19 and x20 and x16 and x18 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( not x21 and not x22 and x23 and x19 and x20 and x16 and not x18 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x21 and not x22 and x23 and x19 and x20 and not x16 and x17 and x18 ) = '1' then
         y24 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s157;

      elsif ( not x21 and not x22 and x23 and x19 and x20 and not x16 and x17 and not x18 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         y20 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s227;

      elsif ( not x21 and not x22 and x23 and x19 and x20 and not x16 and not x17 and x18 and x11 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s247;

      elsif ( not x21 and not x22 and x23 and x19 and x20 and not x16 and not x17 and x18 and not x11 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and x23 and x19 and x20 and not x16 and not x17 and x18 and not x11 and x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and x19 and x20 and not x16 and not x17 and x18 and not x11 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and x19 and x20 and not x16 and not x17 and not x18 and x10 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s247;

      elsif ( not x21 and not x22 and x23 and x19 and x20 and not x16 and not x17 and not x18 and not x10 and x9 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and x23 and x19 and x20 and not x16 and not x17 and not x18 and not x10 and x9 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and x19 and x20 and not x16 and not x17 and not x18 and not x10 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and x19 and not x20 and x17 and x16 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s203;

      elsif ( not x21 and not x22 and x23 and x19 and not x20 and x17 and not x16 and x18 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x21 and not x22 and x23 and x19 and not x20 and x17 and not x16 and not x18 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s233;

      elsif ( not x21 and not x22 and x23 and x19 and not x20 and not x17 and x18 and x16 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s234;

      elsif ( not x21 and not x22 and x23 and x19 and not x20 and not x17 and x18 and not x16 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s235;

      elsif ( not x21 and not x22 and x23 and x19 and not x20 and not x17 and not x18 and x3 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x21 and not x22 and x23 and x19 and not x20 and not x17 and not x18 and not x3 and x5 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( not x21 and not x22 and x23 and x19 and not x20 and not x17 and not x18 and not x3 and not x5 and x16 ) = '1' then
         y5 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s227;

      elsif ( not x21 and not x22 and x23 and x19 and not x20 and not x17 and not x18 and not x3 and not x5 and not x16 ) = '1' then
         y16 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s227;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and x16 and x3 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and x16 and not x3 and x5 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and x16 and not x3 and not x5 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and x17 and x18 and x3 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and x17 and x18 and not x3 and x5 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and x17 and x18 and not x3 and not x5 ) = '1' then
         y8 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s227;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and x17 and not x18 and x15 and x3 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and x17 and not x18 and x15 and not x3 and x5 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and x17 and not x18 and x15 and not x3 and not x5 ) = '1' then
         y8 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s227;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and x17 and not x18 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and not x17 and x18 and x13 and x3 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and not x17 and x18 and x13 and not x3 and x5 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and not x17 and x18 and x13 and not x3 and not x5 ) = '1' then
         y8 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s227;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and not x17 and x18 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and not x17 and not x18 and x12 and x3 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and not x17 and not x18 and x12 and not x3 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and not x17 and not x18 and not x12 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and not x17 and not x18 and not x12 and x9 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and not x17 and not x18 and not x12 and x9 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and not x19 and x20 and not x16 and not x17 and not x18 and not x12 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and not x19 and not x20 and x3 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x21 and not x22 and x23 and not x19 and not x20 and not x3 and x5 ) = '1' then
         y12 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s237;

      elsif ( not x21 and not x22 and x23 and not x19 and not x20 and not x3 and not x5 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      else
         current_group15m <= s1;

      end if;

   when s241 =>
         y7 <= '1' ;
         current_group15m <= s338;

   when s242 =>
      if ( x65 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      else
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s51;

      end if;

   when s243 =>
      if ( x21 and x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and x8 and not x9 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x21 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s117;

      elsif ( not x21 and x22 and not x12 and x8 and x9 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and not x12 and x8 and not x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and not x12 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x12 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x12 and x23 ) = '1' then
         y6 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s247;

      elsif ( not x21 and not x22 and x12 and not x23 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x21 and not x22 and not x12 and x23 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and not x12 and x23 and x9 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and not x12 and x23 and x9 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x12 and x23 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x12 and not x23 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and not x12 and not x23 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and not x12 and not x23 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s244 =>
      if ( x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x8 and not x9 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s245 =>
         y3 <= '1' ;
         y12 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s406;

   when s246 =>
      if ( x65 and x67 ) = '1' then
         y8 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s407;

      elsif ( x65 and not x67 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x65 and x21 and x3 and x4 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( not x65 and x21 and x3 and not x4 and x5 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( not x65 and x21 and x3 and not x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and not x3 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and not x22 and x8 and x9 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x65 and not x21 and not x22 and x8 and not x9 and x10 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x65 and not x21 and not x22 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s247 =>
      if ( x21 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s238;

      elsif ( not x21 and x22 and x23 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x21 and x22 and x23 and not x12 and x8 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x23 and not x12 and x8 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and x22 and x23 and not x12 and x8 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and not x12 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 ) = '1' then
         y14 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s116;

      elsif ( not x21 and not x22 and x23 and x9 and x10 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and x23 and x9 and not x10 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x22 and x23 and x9 and not x10 and not x11 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and not x9 ) = '1' then
         current_group15m <= s1;

      else
         y6 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s223;

      end if;

   when s248 =>
      if ( x22 and x21 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( x22 and not x21 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s409;

      elsif ( not x22 and x19 and x21 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( not x22 and x19 and not x21 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s409;

      else
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      end if;

   when s249 =>
      if ( x21 and x18 and x16 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( x21 and x18 and not x16 and x13 and x15 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( x21 and x18 and not x16 and x13 and not x15 and x17 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s409;

      elsif ( x21 and x18 and not x16 and x13 and not x15 and not x17 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( x21 and x18 and not x16 and not x13 and x17 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s409;

      elsif ( x21 and x18 and not x16 and not x13 and not x17 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( x21 and not x18 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s409;

      elsif ( not x21 and x19 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( not x21 and not x19 and x22 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( not x21 and not x19 and not x22 and x20 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s409;

      elsif ( not x21 and not x19 and not x22 and not x20 and x16 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( not x21 and not x19 and not x22 and not x20 and not x16 and x15 and x13 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( not x21 and not x19 and not x22 and not x20 and not x16 and x15 and not x13 and x17 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s409;

      elsif ( not x21 and not x19 and not x22 and not x20 and not x16 and x15 and not x13 and not x17 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( not x21 and not x19 and not x22 and not x20 and not x16 and not x15 and x17 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s409;

      else
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      end if;

   when s250 =>
      if ( x65 and x60 and x61 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s68;

      elsif ( x65 and x60 and not x61 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      elsif ( x65 and not x60 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      elsif ( not x65 and x23 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s410;

      elsif ( not x65 and not x23 and x19 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s285;

      else
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s84;

      end if;

   when s251 =>
      if ( x60 and x61 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s256;

      elsif ( x60 and not x61 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      else
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      end if;

   when s252 =>
      if ( x60 and x7 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x60 and not x7 and x61 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x60 and not x7 and x61 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x60 and not x7 and x61 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x60 and not x7 and x61 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x60 and not x7 and not x61 ) = '1' then
         current_group15m <= s39;

      elsif ( not x60 and x61 and x62 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x60 and x61 and x62 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x60 and x61 and x62 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( not x60 and x61 and x62 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x60 and x61 and not x62 and x7 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( not x60 and x61 and not x62 and not x7 ) = '1' then
         current_group15m <= s39;

      elsif ( not x60 and not x61 and x62 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      else
         current_group15m <= s40;

      end if;

   when s253 =>
      if ( x60 and x61 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s257;

      elsif ( x60 and not x61 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      else
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      end if;

   when s254 =>
      if ( x65 and x60 and x61 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x60 and x61 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x60 and x61 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x60 and x61 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x60 and not x61 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x60 and not x61 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x60 and not x61 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x60 and not x61 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and not x60 and x61 and x62 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and not x60 and x61 and x62 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and not x60 and x61 and x62 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x60 and x61 and x62 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x60 and x61 and not x62 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x60 and x61 and not x62 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x60 and x61 and not x62 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and not x60 and x61 and not x62 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and not x60 and not x61 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and x20 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and not x20 and x18 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x20 and x18 and not x13 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x65 and not x20 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s255 =>
      if ( x67 and x22 and x4 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x67 and x22 and not x4 and x20 and x15 and x8 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x67 and x22 and not x4 and x20 and x15 and not x8 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x67 and x22 and not x4 and x20 and not x15 and x16 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s302;

      elsif ( x67 and x22 and not x4 and x20 and not x15 and not x16 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s122;

      elsif ( x67 and x22 and not x4 and not x20 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s368;

      elsif ( x67 and not x22 and x23 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x67 and not x22 and not x23 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x61 and x60 and x3 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s118;

      elsif ( not x67 and x61 and x60 and not x3 and x18 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s38;

      elsif ( not x67 and x61 and x60 and not x3 and not x18 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s319;

      elsif ( not x67 and x61 and not x60 and x62 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x67 and x61 and not x60 and x62 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x67 and x61 and not x60 and x62 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x61 and not x60 and x62 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x61 and not x60 and not x62 and x19 and x15 ) = '1' then
         current_group15m <= s73;

      elsif ( not x67 and x61 and not x60 and not x62 and x19 and not x15 and x16 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s291;

      elsif ( not x67 and x61 and not x60 and not x62 and x19 and not x15 and not x16 ) = '1' then
         current_group15m <= s73;

      elsif ( not x67 and x61 and not x60 and not x62 and not x19 ) = '1' then
         y4 <= '1' ;
         y13 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s64;

      elsif ( not x67 and not x61 and x60 and x19 and x15 ) = '1' then
         current_group15m <= s73;

      elsif ( not x67 and not x61 and x60 and x19 and not x15 and x16 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s291;

      elsif ( not x67 and not x61 and x60 and x19 and not x15 and not x16 ) = '1' then
         current_group15m <= s73;

      elsif ( not x67 and not x61 and x60 and not x19 ) = '1' then
         y4 <= '1' ;
         y13 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s64;

      elsif ( not x67 and not x61 and not x60 and x62 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and not x61 and not x60 and not x62 and x18 and x15 and x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( not x67 and not x61 and not x60 and not x62 and x18 and x15 and not x7 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x67 and not x61 and not x60 and not x62 and x18 and x15 and not x7 and not x11 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s254;

      elsif ( not x67 and not x61 and not x60 and not x62 and x18 and not x15 and x16 and x4 ) = '1' then
         current_group15m <= s40;

      elsif ( not x67 and not x61 and not x60 and not x62 and x18 and not x15 and x16 and not x4 and x11 and x9 ) = '1' then
         current_group15m <= s40;

      elsif ( not x67 and not x61 and not x60 and not x62 and x18 and not x15 and x16 and not x4 and x11 and not x9 and x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( not x67 and not x61 and not x60 and not x62 and x18 and not x15 and x16 and not x4 and x11 and not x9 and not x7 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s118;

      elsif ( not x67 and not x61 and not x60 and not x62 and x18 and not x15 and x16 and not x4 and not x11 and x9 and x7 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( not x67 and not x61 and not x60 and not x62 and x18 and not x15 and x16 and not x4 and not x11 and x9 and not x7 and x10 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( not x67 and not x61 and not x60 and not x62 and x18 and not x15 and x16 and not x4 and not x11 and x9 and not x7 and not x10 ) = '1' then
         current_group15m <= s40;

      elsif ( not x67 and not x61 and not x60 and not x62 and x18 and not x15 and x16 and not x4 and not x11 and not x9 and x7 and x8 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( not x67 and not x61 and not x60 and not x62 and x18 and not x15 and x16 and not x4 and not x11 and not x9 and x7 and not x8 ) = '1' then
         current_group15m <= s40;

      elsif ( not x67 and not x61 and not x60 and not x62 and x18 and not x15 and x16 and not x4 and not x11 and not x9 and not x7 and x12 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( not x67 and not x61 and not x60 and not x62 and x18 and not x15 and x16 and not x4 and not x11 and not x9 and not x7 and not x12 ) = '1' then
         current_group15m <= s40;

      elsif ( not x67 and not x61 and not x60 and not x62 and x18 and not x15 and not x16 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      else
         y4 <= '1' ;
         y13 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s64;

      end if;

   when s256 =>
      if ( x60 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s68;

      else
         y14 <= '1' ;
         current_group15m <= s155;

      end if;

   when s257 =>
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s68;

   when s258 =>
      if ( x60 and x61 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( x60 and not x61 and x2 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x60 and not x61 and not x2 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x60 and x61 and x62 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x60 and x61 and x62 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x60 and x61 and x62 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( not x60 and x61 and x62 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x60 and x61 and not x62 and x2 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x60 and x61 and not x62 and not x2 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x60 and not x61 and x62 and x7 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x60 and not x61 and x62 and not x7 ) = '1' then
         current_group15m <= s40;

      else
         y12 <= '1' ;
         current_group15m <= s100;

      end if;

   when s259 =>
      if ( x21 and x20 and x10 and x12 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x20 and x10 and x12 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x20 and x10 and x12 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x20 and x10 and x12 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x20 and x10 and not x12 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s302;

      elsif ( x21 and x20 and not x10 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x20 and not x10 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x20 and not x10 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x20 and not x10 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x20 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x20 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x21 and not x20 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x20 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x10 and x12 and x19 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x21 and x10 and x12 and x19 and not x14 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x21 and x10 and x12 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x10 and x12 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x10 and not x12 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( not x21 and not x10 and x19 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x21 and not x10 and x19 and not x14 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x21 and not x10 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s260 =>
      if ( x60 and x61 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x60 and x61 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x60 and x61 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x60 and x61 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x60 and not x61 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x60 and not x61 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x60 and not x61 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x60 and not x61 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( not x60 and x61 and x62 ) = '1' then
         current_group15m <= s1;

      elsif ( not x60 and x61 and not x62 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x60 and x61 and not x62 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x60 and x61 and not x62 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( not x60 and x61 and not x62 and not x18 ) = '1' then
         current_group15m <= s39;

      else
         current_group15m <= s40;

      end if;

   when s261 =>
      if ( x61 and x60 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x61 and x60 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x61 and x60 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x61 and x60 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x61 and not x60 and x62 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x61 and not x60 and x62 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x61 and not x60 and x62 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x61 and not x60 and x62 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x61 and not x60 and not x62 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x61 and not x60 and not x62 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x61 and not x60 and not x62 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x61 and not x60 and not x62 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( not x61 and x60 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x61 and x60 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x61 and x60 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( not x61 and x60 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( not x61 and not x60 and x62 and x19 and x15 and x12 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s292;

      elsif ( not x61 and not x60 and x62 and x19 and x15 and x12 and not x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s290;

      elsif ( not x61 and not x60 and x62 and x19 and x15 and not x12 and x7 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s63;

      elsif ( not x61 and not x60 and x62 and x19 and x15 and not x12 and not x7 ) = '1' then
         y2 <= '1' ;
         y10 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s263;

      elsif ( not x61 and not x60 and x62 and x19 and not x15 and x16 and x7 and x12 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s290;

      elsif ( not x61 and not x60 and x62 and x19 and not x15 and x16 and x7 and not x12 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s262;

      elsif ( not x61 and not x60 and x62 and x19 and not x15 and x16 and not x7 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s258;

      elsif ( not x61 and not x60 and x62 and x19 and not x15 and not x16 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x61 and not x60 and x62 and x19 and not x15 and not x16 and not x7 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x61 and not x60 and x62 and not x19 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s411;

      else
         current_group15m <= s40;

      end if;

   when s262 =>
      if ( x65 and x61 and x60 and x19 and x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x61 and x60 and x19 and not x13 and x14 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x65 and x61 and x60 and x19 and not x13 and not x14 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x61 and x60 and not x19 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and x61 and not x60 and x62 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x61 and not x60 and x62 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x65 and x61 and not x60 and x62 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x61 and not x60 and x62 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x61 and not x60 and not x62 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x61 and not x60 and not x62 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x61 and not x60 and not x62 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and x61 and not x60 and not x62 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and not x61 and x60 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x61 and x60 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x61 and x60 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and not x61 and x60 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( x65 and not x61 and not x60 and x62 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s258;

      elsif ( x65 and not x61 and not x60 and not x62 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and x21 and x10 and x5 and x16 and x15 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s399;

      elsif ( not x65 and x21 and x10 and x5 and x16 and not x15 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x21 and x10 and x5 and not x16 and x17 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s215;

      elsif ( not x65 and x21 and x10 and x5 and not x16 and not x17 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s215;

      elsif ( not x65 and x21 and x10 and not x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x21 and not x10 and x16 and x5 and x15 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s215;

      elsif ( not x65 and x21 and not x10 and x16 and x5 and not x15 ) = '1' then
         y13 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s284;

      elsif ( not x65 and x21 and not x10 and x16 and not x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x21 and not x10 and not x16 and x17 and x14 and x13 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x21 and not x10 and not x16 and x17 and x14 and not x13 and x15 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x21 and not x10 and not x16 and x17 and x14 and not x13 and not x15 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x21 and not x10 and not x16 and x17 and x14 and not x13 and not x15 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x21 and not x10 and not x16 and x17 and x14 and not x13 and not x15 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and not x10 and not x16 and x17 and x14 and not x13 and not x15 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and not x10 and not x16 and x17 and not x14 and x15 and x12 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x21 and not x10 and not x16 and x17 and not x14 and x15 and not x12 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x21 and not x10 and not x16 and x17 and not x14 and x15 and not x12 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x21 and not x10 and not x16 and x17 and not x14 and x15 and not x12 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and not x10 and not x16 and x17 and not x14 and x15 and not x12 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and not x10 and not x16 and x17 and not x14 and not x15 and x11 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x21 and not x10 and not x16 and x17 and not x14 and not x15 and not x11 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x21 and not x10 and not x16 and x17 and not x14 and not x15 and not x11 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x21 and not x10 and not x16 and x17 and not x14 and not x15 and not x11 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and not x10 and not x16 and x17 and not x14 and not x15 and not x11 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and not x10 and not x16 and not x17 and x5 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      elsif ( not x65 and x21 and not x10 and not x16 and not x17 and not x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and not x21 and x22 and x17 and x18 and x10 and x15 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s363;

      elsif ( not x65 and not x21 and x22 and x17 and x18 and x10 and not x15 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s13;

      elsif ( not x65 and not x21 and x22 and x17 and x18 and not x10 and x14 and x15 and x9 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s310;

      elsif ( not x65 and not x21 and x22 and x17 and x18 and not x10 and x14 and x15 and not x9 and x7 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and not x21 and x22 and x17 and x18 and not x10 and x14 and x15 and not x9 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and x17 and x18 and not x10 and x14 and not x15 and x8 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x65 and not x21 and x22 and x17 and x18 and not x10 and x14 and not x15 and not x8 and x7 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and not x21 and x22 and x17 and x18 and not x10 and x14 and not x15 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and x17 and x18 and not x10 and not x14 and x15 and x9 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s188;

      elsif ( not x65 and not x21 and x22 and x17 and x18 and not x10 and not x14 and x15 and not x9 and x8 and x7 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and not x21 and x22 and x17 and x18 and not x10 and not x14 and x15 and not x9 and x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and x17 and x18 and not x10 and not x14 and x15 and not x9 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and x17 and x18 and not x10 and not x14 and not x15 and x8 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s188;

      elsif ( not x65 and not x21 and x22 and x17 and x18 and not x10 and not x14 and not x15 and not x8 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and not x21 and x22 and x17 and not x18 and x14 and x10 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s335;

      elsif ( not x65 and not x21 and x22 and x17 and not x18 and x14 and not x10 and x15 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s410;

      elsif ( not x65 and not x21 and x22 and x17 and not x18 and x14 and not x10 and not x15 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and not x21 and x22 and x17 and not x18 and not x14 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( not x65 and not x21 and x22 and x17 and not x18 and not x14 and not x2 and x5 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s226;

      elsif ( not x65 and not x21 and x22 and x17 and not x18 and not x14 and not x2 and not x5 and x15 and x10 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s219;

      elsif ( not x65 and not x21 and x22 and x17 and not x18 and not x14 and not x2 and not x5 and x15 and not x10 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s309;

      elsif ( not x65 and not x21 and x22 and x17 and not x18 and not x14 and not x2 and not x5 and not x15 and x10 ) = '1' then
         y2 <= '1' ;
         y16 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s124;

      elsif ( not x65 and not x21 and x22 and x17 and not x18 and not x14 and not x2 and not x5 and not x15 and not x10 ) = '1' then
         y14 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s216;

      elsif ( not x65 and not x21 and x22 and not x17 and x2 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and x10 and x5 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s226;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and x10 and not x5 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s219;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and not x10 and x14 and x15 and x5 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s226;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and not x10 and x14 and x15 and not x5 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and not x10 and x14 and not x15 and x13 and x5 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s226;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and not x10 and x14 and not x15 and x13 and not x5 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and not x10 and x14 and not x15 and not x13 and x7 and x8 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and not x10 and x14 and not x15 and not x13 and x7 and not x8 and x9 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and not x10 and x14 and not x15 and not x13 and x7 and not x8 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and not x10 and x14 and not x15 and not x13 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and not x10 and not x14 and x15 and x12 and x5 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s226;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and not x10 and not x14 and x15 and x12 and not x5 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and not x10 and not x14 and x15 and not x12 and x7 and x8 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and not x10 and not x14 and x15 and not x12 and x7 and not x8 and x9 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and not x10 and not x14 and x15 and not x12 and x7 and not x8 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and not x10 and not x14 and x15 and not x12 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and not x10 and not x14 and not x15 and x11 and x5 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s226;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and not x10 and not x14 and not x15 and x11 and not x5 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and not x10 and not x14 and not x15 and not x11 and x7 and x8 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and not x10 and not x14 and not x15 and not x11 and x7 and not x8 and x9 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and not x10 and not x14 and not x15 and not x11 and x7 and not x8 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and x18 and not x10 and not x14 and not x15 and not x11 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and not x18 and x5 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and not x18 and not x5 and x10 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s219;

      elsif ( not x65 and not x21 and x22 and not x17 and not x2 and not x18 and not x5 and not x10 ) = '1' then
         y9 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s311;

      else
         current_group15m <= s1;

      end if;

   when s263 =>
      if ( x60 and x61 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x60 and not x61 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x60 and not x61 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x60 and not x61 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( x60 and not x61 and not x18 ) = '1' then
         current_group15m <= s39;

      elsif ( not x60 and x61 and x62 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x60 and x61 and x62 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x60 and x61 and x62 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( not x60 and x61 and x62 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x60 and x61 and not x62 and x18 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x60 and x61 and not x62 and x18 and not x13 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x60 and x61 and not x62 and x18 and not x13 and not x14 ) = '1' then
         current_group15m <= s39;

      elsif ( not x60 and x61 and not x62 and not x18 ) = '1' then
         current_group15m <= s39;

      else
         current_group15m <= s40;

      end if;

   when s264 =>
      if ( x65 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s68;

      else
         y4 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s370;

      end if;

   when s265 =>
      if ( x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x12 ) = '1' then
         y10 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s273;

      elsif ( not x21 and x22 and not x12 and x6 and x7 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x21 and x22 and not x12 and x6 and not x7 and x8 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x21 and x22 and not x12 and x6 and not x7 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x12 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x7 and x18 and x15 ) = '1' then
         y8 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s82;

      elsif ( not x21 and not x22 and x7 and x18 and not x15 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s374;

      elsif ( not x21 and not x22 and x7 and not x18 and x19 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s320;

      elsif ( not x21 and not x22 and x7 and not x18 and x19 and not x15 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x21 and not x22 and x7 and not x18 and not x19 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      else
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s385;

      end if;

   when s266 =>
      if ( x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x7 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x21 and x22 and not x7 and x8 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x21 and x22 and not x7 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x8 and x9 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x21 and not x22 and x8 and not x9 and x10 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x21 and not x22 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s267 =>
      if ( x65 and x2 and x18 and x19 and x14 and x17 and x20 and x16 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x65 and x2 and x18 and x19 and x14 and x17 and x20 and not x16 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s346;

      elsif ( x65 and x2 and x18 and x19 and x14 and x17 and not x20 and x16 ) = '1' then
         y13 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s347;

      elsif ( x65 and x2 and x18 and x19 and x14 and x17 and not x20 and not x16 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x65 and x2 and x18 and x19 and x14 and not x17 and x20 and x8 and x16 ) = '1' then
         y13 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s347;

      elsif ( x65 and x2 and x18 and x19 and x14 and not x17 and x20 and x8 and not x16 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and x18 and x19 and x14 and not x17 and x20 and not x8 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and x18 and x19 and x14 and not x17 and not x20 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and x18 and x19 and not x14 and x15 and x17 and x20 and x16 ) = '1' then
         y9 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and x18 and x19 and not x14 and x15 and x17 and x20 and not x16 ) = '1' then
         y4 <= '1' ;
         y12 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and x18 and x19 and not x14 and x15 and x17 and not x20 and x16 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s346;

      elsif ( x65 and x2 and x18 and x19 and not x14 and x15 and x17 and not x20 and not x16 ) = '1' then
         y9 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and x18 and x19 and not x14 and x15 and not x17 and x16 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and x18 and x19 and not x14 and x15 and not x17 and not x16 and x13 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and x18 and x19 and not x14 and x15 and not x17 and not x16 and not x13 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and x18 and x19 and not x14 and x15 and not x17 and not x16 and not x13 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and x18 and x19 and not x14 and x15 and not x17 and not x16 and not x13 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and x19 and not x14 and x15 and not x17 and not x16 and not x13 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and x19 and not x14 and not x15 and x17 and x16 and x7 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x65 and x2 and x18 and x19 and not x14 and not x15 and x17 and x16 and not x7 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and x18 and x19 and not x14 and not x15 and x17 and x16 and not x7 and x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and x19 and not x14 and not x15 and x17 and x16 and not x7 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and x19 and not x14 and not x15 and x17 and not x16 and x6 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x65 and x2 and x18 and x19 and not x14 and not x15 and x17 and not x16 and not x6 and x5 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and x18 and x19 and not x14 and not x15 and x17 and not x16 and not x6 and x5 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and x19 and not x14 and not x15 and x17 and not x16 and not x6 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and x19 and not x14 and not x15 and not x17 and x16 and x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and x18 and x19 and not x14 and not x15 and not x17 and x16 and not x12 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and x18 and x19 and not x14 and not x15 and not x17 and x16 and not x12 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and x18 and x19 and not x14 and not x15 and not x17 and x16 and not x12 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and x19 and not x14 and not x15 and not x17 and x16 and not x12 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and x19 and not x14 and not x15 and not x17 and not x16 and x11 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and x18 and x19 and not x14 and not x15 and not x17 and not x16 and not x11 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and x18 and x19 and not x14 and not x15 and not x17 and not x16 and not x11 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and x18 and x19 and not x14 and not x15 and not x17 and not x16 and not x11 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and x19 and not x14 and not x15 and not x17 and not x16 and not x11 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and not x19 and x17 and x20 and x14 and x13 ) = '1' then
         y10 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s349;

      elsif ( x65 and x2 and x18 and not x19 and x17 and x20 and x14 and not x13 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x65 and x2 and x18 and not x19 and x17 and x20 and not x14 and x13 ) = '1' then
         y2 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s349;

      elsif ( x65 and x2 and x18 and not x19 and x17 and x20 and not x14 and not x13 and x6 ) = '1' then
         y6 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s102;

      elsif ( x65 and x2 and x18 and not x19 and x17 and x20 and not x14 and not x13 and not x6 and x5 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and x18 and not x19 and x17 and x20 and not x14 and not x13 and not x6 and x5 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and not x19 and x17 and x20 and not x14 and not x13 and not x6 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and not x19 and x17 and not x20 and x15 and x14 ) = '1' then
         y10 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s349;

      elsif ( x65 and x2 and x18 and not x19 and x17 and not x20 and x15 and not x14 ) = '1' then
         y6 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s102;

      elsif ( x65 and x2 and x18 and not x19 and x17 and not x20 and not x15 and x14 ) = '1' then
         y15 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s350;

      elsif ( x65 and x2 and x18 and not x19 and x17 and not x20 and not x15 and not x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and x20 and x13 and x12 and x14 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and x20 and x13 and x12 and not x14 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and x20 and x13 and x12 and not x14 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and x20 and x13 and x12 and not x14 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and x20 and x13 and x12 and not x14 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and x20 and x13 and not x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and x20 and not x13 and x11 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and x20 and not x13 and x11 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and x20 and not x13 and x11 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and x20 and not x13 and x11 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and x20 and not x13 and not x11 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and not x20 and x15 and x12 and x8 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s241;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and not x20 and x15 and x12 and not x8 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and not x20 and x15 and not x12 and x14 and x8 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s241;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and not x20 and x15 and not x12 and x14 and not x8 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and not x20 and x15 and not x12 and not x14 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and not x20 and x15 and not x12 and not x14 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and not x20 and x15 and not x12 and not x14 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and not x20 and x15 and not x12 and not x14 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and not x20 and not x15 and x14 and x13 and x8 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s241;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and not x20 and not x15 and x14 and x13 and not x8 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and not x20 and not x15 and x14 and not x13 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and not x20 and not x15 and x14 and not x13 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and not x20 and not x15 and x14 and not x13 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and not x20 and not x15 and x14 and not x13 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and not x20 and not x15 and not x14 and x11 and x8 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s241;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and not x20 and not x15 and not x14 and x11 and not x8 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and not x20 and not x15 and not x14 and not x11 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and not x20 and not x15 and not x14 and not x11 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and not x20 and not x15 and not x14 and not x11 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and x18 and not x19 and not x17 and not x20 and not x15 and not x14 and not x11 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and not x18 and x17 and x19 and x15 and x14 and x20 ) = '1' then
         y29 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and x19 and x15 and x14 and not x20 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and x19 and x15 and not x14 and x16 and x20 and x13 ) = '1' then
         y29 <= '1' ;
         y31 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and x19 and x15 and not x14 and x16 and x20 and not x13 ) = '1' then
         y29 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and x19 and x15 and not x14 and x16 and not x20 and x13 ) = '1' then
         y29 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and x19 and x15 and not x14 and x16 and not x20 and not x13 ) = '1' then
         y4 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and x19 and x15 and not x14 and not x16 and x20 ) = '1' then
         y4 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and x19 and x15 and not x14 and not x16 and not x20 and x4 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s348;

      elsif ( x65 and x2 and not x18 and x17 and x19 and x15 and not x14 and not x16 and not x20 and not x4 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( x65 and x2 and not x18 and x17 and x19 and not x15 and x14 and x16 and x20 ) = '1' then
         y29 <= '1' ;
         y31 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and x19 and not x15 and x14 and x16 and not x20 ) = '1' then
         y29 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and x19 and not x15 and x14 and not x16 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and not x18 and x17 and x19 and not x15 and not x14 and x20 and x8 and x16 ) = '1' then
         y4 <= '1' ;
         y18 <= '1' ;
         y29 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and x19 and not x15 and not x14 and x20 and x8 and not x16 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and x19 and not x15 and not x14 and x20 and not x8 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and not x18 and x17 and x19 and not x15 and not x14 and not x20 and x8 and x16 ) = '1' then
         y4 <= '1' ;
         y17 <= '1' ;
         y29 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and x19 and not x15 and not x14 and not x20 and x8 and not x16 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and x19 and not x15 and not x14 and not x20 and not x8 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and x20 and x16 and x14 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and x20 and x16 and not x14 and x15 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and x20 and x16 and not x14 and x15 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and x20 and x16 and not x14 and x15 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and x20 and x16 and not x14 and x15 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and x20 and x16 and not x14 and not x15 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and x20 and not x16 and x13 and x14 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and x20 and not x16 and x13 and x14 and not x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and x20 and not x16 and x13 and not x14 and x4 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and x20 and not x16 and x13 and not x14 and not x4 ) = '1' then
         y4 <= '1' ;
         y12 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and x20 and not x16 and not x13 and x8 ) = '1' then
         y13 <= '1' ;
         y20 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s347;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and x20 and not x16 and not x13 and not x8 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and not x20 and x14 and x16 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s346;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and not x20 and x14 and not x16 and x15 and x13 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and not x20 and x14 and not x16 and x15 and not x13 ) = '1' then
         y4 <= '1' ;
         y12 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and not x20 and x14 and not x16 and not x15 ) = '1' then
         y9 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and not x20 and not x14 and x15 and x16 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and not x20 and not x14 and x15 and not x16 and x8 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         y19 <= '1' ;
         y21 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s351;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and not x20 and not x14 and x15 and not x16 and not x8 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and not x20 and not x14 and not x15 and x8 and x16 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and not x20 and not x14 and not x15 and x8 and x16 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and not x20 and not x14 and not x15 and x8 and x16 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and not x20 and not x14 and not x15 and x8 and x16 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and not x20 and not x14 and not x15 and x8 and not x16 ) = '1' then
         y2 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s349;

      elsif ( x65 and x2 and not x18 and x17 and not x19 and not x20 and not x14 and not x15 and not x8 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and x2 and not x18 and not x17 and x8 ) = '1' then
         y4 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s395;

      elsif ( x65 and x2 and not x18 and not x17 and not x8 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s412;

      elsif ( x65 and not x2 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x65 and x21 and x4 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( not x65 and x21 and not x4 and x5 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( not x65 and x21 and not x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and x6 and x7 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x65 and not x21 and x22 and x6 and not x7 and x8 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x65 and not x21 and x22 and x6 and not x7 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and not x22 and x8 and x9 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x65 and not x21 and not x22 and x8 and not x9 and x10 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x65 and not x21 and not x22 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s268 =>
         y10 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s273;

   when s269 =>
      if ( x21 and x66 and x19 and x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x21 and x66 and x19 and not x15 and x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x21 and x66 and x19 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x66 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x66 and x3 and x4 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( x21 and not x66 and x3 and not x4 and x5 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( x21 and not x66 and x3 and not x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x66 and not x3 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x66 and x20 and x15 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( not x21 and x66 and x20 and not x15 and x14 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( not x21 and x66 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x66 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x66 and x22 and x6 and x7 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x21 and not x66 and x22 and x6 and not x7 and x8 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x21 and not x66 and x22 and x6 and not x7 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x66 and x22 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x66 and not x22 and x8 and x9 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x21 and not x66 and not x22 and x8 and not x9 and x10 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x21 and not x66 and not x22 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s270 =>
      if ( x21 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s394;

      elsif ( not x21 and x6 and x7 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x21 and x6 and not x7 and x8 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x21 and x6 and not x7 and not x8 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s271 =>
         y5 <= '1' ;
         current_group15m <= s101;

   when s272 =>
      if ( x21 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      else
         y5 <= '1' ;
         current_group15m <= s101;

      end if;

   when s273 =>
      if ( x21 and x3 and x4 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( x21 and x3 and not x4 and x5 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( x21 and x3 and not x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x3 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x6 and x7 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x21 and x22 and x6 and not x7 and x8 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x21 and x22 and x6 and not x7 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x8 and x9 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x21 and not x22 and x8 and not x9 and x10 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x21 and not x22 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s274 =>
      if ( x21 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x21 and x22 and x5 and x18 and x17 and x12 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s271;

      elsif ( not x21 and x22 and x5 and x18 and x17 and not x12 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s271;

      elsif ( not x21 and x22 and x5 and x18 and not x17 and x12 ) = '1' then
         y6 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s386;

      elsif ( not x21 and x22 and x5 and x18 and not x17 and not x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s374;

      elsif ( not x21 and x22 and x5 and not x18 and x19 and x12 and x17 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s271;

      elsif ( not x21 and x22 and x5 and not x18 and x19 and x12 and not x17 ) = '1' then
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s388;

      elsif ( not x21 and x22 and x5 and not x18 and x19 and not x12 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( not x21 and x22 and x5 and not x18 and not x19 and x12 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s271;

      elsif ( not x21 and x22 and x5 and not x18 and not x19 and not x12 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x21 and x22 and not x5 ) = '1' then
         y14 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s376;

      elsif ( not x21 and not x22 and x18 and x8 and x9 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x21 and not x22 and x18 and x8 and not x9 and x10 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x21 and not x22 and x18 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x18 and not x8 ) = '1' then
         current_group15m <= s1;

      else
         y18 <= '1' ;
         current_group15m <= s114;

      end if;

   when s275 =>
      if ( x21 and x19 and x18 and x17 and x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s272;

      elsif ( x21 and x19 and x18 and x17 and not x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s272;

      elsif ( x21 and x19 and x18 and not x17 and x12 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x21 and x19 and x18 and not x17 and not x12 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s273;

      elsif ( x21 and x19 and not x18 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s274;

      elsif ( x21 and not x19 and x9 and x20 and x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s272;

      elsif ( x21 and not x19 and x9 and x20 and not x12 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s105;

      elsif ( x21 and not x19 and x9 and not x20 and x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s270;

      elsif ( x21 and not x19 and x9 and not x20 and not x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s109;

      elsif ( x21 and not x19 and not x9 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s274;

      elsif ( not x21 and x22 and x3 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s274;

      elsif ( not x21 and x22 and not x3 and x5 and x18 and x17 and x12 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s271;

      elsif ( not x21 and x22 and not x3 and x5 and x18 and x17 and not x12 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s271;

      elsif ( not x21 and x22 and not x3 and x5 and x18 and not x17 and x12 ) = '1' then
         y6 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s386;

      elsif ( not x21 and x22 and not x3 and x5 and x18 and not x17 and not x12 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s374;

      elsif ( not x21 and x22 and not x3 and x5 and not x18 and x19 and x12 and x17 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s271;

      elsif ( not x21 and x22 and not x3 and x5 and not x18 and x19 and x12 and not x17 ) = '1' then
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s388;

      elsif ( not x21 and x22 and not x3 and x5 and not x18 and x19 and not x12 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( not x21 and x22 and not x3 and x5 and not x18 and not x19 and x12 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s271;

      elsif ( not x21 and x22 and not x3 and x5 and not x18 and not x19 and not x12 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x21 and x22 and not x3 and not x5 ) = '1' then
         y14 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s376;

      elsif ( not x21 and not x22 and x18 and x15 ) = '1' then
         y8 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s82;

      elsif ( not x21 and not x22 and x18 and not x15 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s374;

      elsif ( not x21 and not x22 and not x18 and x19 and x15 and x5 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s413;

      elsif ( not x21 and not x22 and not x18 and x19 and x15 and not x5 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s320;

      elsif ( not x21 and not x22 and not x18 and x19 and not x15 ) = '1' then
         y4 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s273;

      else
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      end if;

   when s276 =>
      if ( x16 and x15 and x10 and x12 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x16 and x15 and x10 and not x12 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( x16 and x15 and not x10 and x11 and x12 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s126;

      elsif ( x16 and x15 and not x10 and x11 and not x12 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s192;

      elsif ( x16 and x15 and not x10 and not x11 and x12 and x13 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s125;

      elsif ( x16 and x15 and not x10 and not x11 and x12 and not x13 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x16 and x15 and not x10 and not x11 and x12 and not x13 and x17 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x16 and x15 and not x10 and not x11 and x12 and not x13 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x16 and x15 and not x10 and not x11 and not x12 and x14 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s125;

      elsif ( x16 and x15 and not x10 and not x11 and not x12 and not x14 and x17 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x16 and x15 and not x10 and not x11 and not x12 and not x14 and x17 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x16 and x15 and not x10 and not x11 and not x12 and not x14 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x16 and not x15 and x12 and x10 and x8 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x16 and not x15 and x12 and x10 and x8 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x16 and not x15 and x12 and x10 and x8 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x16 and not x15 and x12 and x10 and x8 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x16 and not x15 and x12 and x10 and not x8 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x16 and not x15 and x12 and x10 and not x8 and not x5 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s132;

      elsif ( x16 and not x15 and x12 and x10 and not x8 and not x5 and not x2 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s199;

      elsif ( x16 and not x15 and x12 and not x10 and x11 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x16 and not x15 and x12 and not x10 and x11 and not x5 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s132;

      elsif ( x16 and not x15 and x12 and not x10 and x11 and not x5 and not x2 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s199;

      elsif ( x16 and not x15 and x12 and not x10 and not x11 and x7 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x16 and not x15 and x12 and not x10 and not x11 and x7 and not x5 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s132;

      elsif ( x16 and not x15 and x12 and not x10 and not x11 and x7 and not x5 and not x2 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s199;

      elsif ( x16 and not x15 and x12 and not x10 and not x11 and not x7 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x16 and not x15 and x12 and not x10 and not x11 and not x7 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x16 and not x15 and x12 and not x10 and not x11 and not x7 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x16 and not x15 and x12 and not x10 and not x11 and not x7 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x16 and not x15 and not x12 and x10 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x16 and not x15 and not x12 and x10 and not x5 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s200;

      elsif ( x16 and not x15 and not x12 and x10 and not x5 and not x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s132;

      elsif ( x16 and not x15 and not x12 and not x10 and x11 and x9 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x16 and not x15 and not x12 and not x10 and x11 and x9 and not x5 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s132;

      elsif ( x16 and not x15 and not x12 and not x10 and x11 and x9 and not x5 and not x2 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s199;

      elsif ( x16 and not x15 and not x12 and not x10 and x11 and not x9 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x16 and not x15 and not x12 and not x10 and x11 and not x9 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x16 and not x15 and not x12 and not x10 and x11 and not x9 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x16 and not x15 and not x12 and not x10 and x11 and not x9 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x16 and not x15 and not x12 and not x10 and not x11 and x8 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( x16 and not x15 and not x12 and not x10 and not x11 and x8 and not x5 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s132;

      elsif ( x16 and not x15 and not x12 and not x10 and not x11 and x8 and not x5 and not x2 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s199;

      elsif ( x16 and not x15 and not x12 and not x10 and not x11 and not x8 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x16 and not x15 and not x12 and not x10 and not x11 and not x8 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x16 and not x15 and not x12 and not x10 and not x11 and not x8 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x16 and not x15 and not x12 and not x10 and not x11 and not x8 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x16 and x15 and x10 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( not x16 and x15 and x10 and not x5 and x11 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s132;

      elsif ( not x16 and x15 and x10 and not x5 and x11 and not x2 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x16 and x15 and x10 and not x5 and not x11 and x12 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s132;

      elsif ( not x16 and x15 and x10 and not x5 and not x11 and x12 and not x2 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s193;

      elsif ( not x16 and x15 and x10 and not x5 and not x11 and not x12 and x2 ) = '1' then
         y8 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s195;

      elsif ( not x16 and x15 and x10 and not x5 and not x11 and not x12 and not x2 ) = '1' then
         y1 <= '1' ;
         y8 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s192;

      elsif ( not x16 and x15 and not x10 and x11 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x16 and x15 and not x10 and not x11 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( not x16 and x15 and not x10 and not x11 and not x5 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s132;

      elsif ( not x16 and x15 and not x10 and not x11 and not x5 and not x2 and x12 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      elsif ( not x16 and x15 and not x10 and not x11 and not x5 and not x2 and not x12 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s198;

      elsif ( not x16 and not x15 and x5 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         current_group15m <= s10;

      elsif ( not x16 and not x15 and not x5 and x2 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s132;

      else
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s390;

      end if;

   when s277 =>
      if ( x20 and x17 and x15 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s198;

      elsif ( x20 and x17 and not x15 and x16 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s59;

      elsif ( x20 and x17 and not x15 and not x16 ) = '1' then
         y7 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s211;

      elsif ( x20 and not x17 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s401;

      elsif ( not x20 and x21 ) = '1' then
         y12 <= '1' ;
         y15 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s401;

      else
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s186;

      end if;

   when s278 =>
      if ( x65 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x24 and x26 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x67 and x24 and not x26 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and x67 and x24 and not x26 and not x4 and x19 and x16 and x11 and x12 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s188;

      elsif ( not x65 and x67 and x24 and not x26 and not x4 and x19 and x16 and x11 and not x12 and x13 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s172;

      elsif ( not x65 and x67 and x24 and not x26 and not x4 and x19 and x16 and x11 and not x12 and not x13 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x65 and x67 and x24 and not x26 and not x4 and x19 and x16 and not x11 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s160;

      elsif ( not x65 and x67 and x24 and not x26 and not x4 and x19 and not x16 and x17 and x11 and x13 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      elsif ( not x65 and x67 and x24 and not x26 and not x4 and x19 and not x16 and x17 and x11 and not x13 ) = '1' then
         y15 <= '1' ;
         y112 <= '1' ;
         current_group15m <= s46;

      elsif ( not x65 and x67 and x24 and not x26 and not x4 and x19 and not x16 and x17 and not x11 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      elsif ( not x65 and x67 and x24 and not x26 and not x4 and x19 and not x16 and not x17 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x65 and x67 and x24 and not x26 and not x4 and not x19 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and x67 and not x24 and x25 and x26 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( not x65 and x67 and not x24 and x25 and not x26 and x15 and x10 and x11 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s187;

      elsif ( not x65 and x67 and not x24 and x25 and not x26 and x15 and x10 and not x11 and x12 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s185;

      elsif ( not x65 and x67 and not x24 and x25 and not x26 and x15 and x10 and not x11 and not x12 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s160;

      elsif ( not x65 and x67 and not x24 and x25 and not x26 and x15 and not x10 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s50;

      elsif ( not x65 and x67 and not x24 and x25 and not x26 and not x15 and x16 and x10 and x12 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( not x65 and x67 and not x24 and x25 and not x26 and not x15 and x16 and x10 and not x12 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and x67 and not x24 and x25 and not x26 and not x15 and x16 and not x10 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( not x65 and x67 and not x24 and x25 and not x26 and not x15 and not x16 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      elsif ( not x65 and x67 and not x24 and not x25 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and x21 and x9 and x3 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x67 and x21 and x9 and not x3 and x4 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x67 and x21 and x9 and not x3 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and x21 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and x22 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x67 and not x21 and x22 and x5 and not x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x65 and not x67 and not x21 and x22 and x5 and not x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x67 and not x21 and x22 and not x5 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s279 =>
      if ( x66 and x21 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( x66 and not x21 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s344;

      elsif ( not x66 and x68 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      else
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s402;

      end if;

   when s280 =>
         y8 <= '1' ;
         y17 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s164;

   when s281 =>
      if ( x24 and x26 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s150;

      elsif ( x24 and not x26 and x16 and x11 and x12 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s188;

      elsif ( x24 and not x26 and x16 and x11 and not x12 and x13 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s172;

      elsif ( x24 and not x26 and x16 and x11 and not x12 and not x13 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x24 and not x26 and x16 and not x11 ) = '1' then
         y5 <= '1' ;
         y14 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s160;

      elsif ( x24 and not x26 and not x16 and x17 and x11 and x13 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      elsif ( x24 and not x26 and not x16 and x17 and x11 and not x13 ) = '1' then
         y15 <= '1' ;
         y112 <= '1' ;
         current_group15m <= s46;

      elsif ( x24 and not x26 and not x16 and x17 and not x11 ) = '1' then
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

      elsif ( x24 and not x26 and not x16 and not x17 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x24 and x25 ) = '1' then
         y36 <= '1' ;
         current_group15m <= s55;

      elsif ( not x24 and not x25 and x26 and x16 and x11 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x24 and not x25 and x26 and x16 and not x11 and x12 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x24 and not x25 and x26 and x16 and not x11 and not x12 and x10 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x24 and not x25 and x26 and x16 and not x11 and not x12 and not x10 ) = '1' then
         y12 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s49;

      elsif ( not x24 and not x25 and x26 and not x16 and x17 and x10 and x12 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( not x24 and not x25 and x26 and not x16 and x17 and x10 and not x12 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x24 and not x25 and x26 and not x16 and x17 and not x10 ) = '1' then
         y13 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s166;

      elsif ( not x24 and not x25 and x26 and not x16 and not x17 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      else
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      end if;

   when s282 =>
      if ( x24 and x26 and x18 and x15 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( x24 and x26 and x18 and not x15 and x14 ) = '1' then
         y6 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s162;

      elsif ( x24 and x26 and x18 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x24 and x26 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x24 and not x26 and x20 and x15 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( x24 and not x26 and x20 and not x15 and x14 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( x24 and not x26 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x24 and not x26 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x25 and x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( not x24 and x25 and x19 and not x14 and not x13 and x26 ) = '1' then
         current_group15m <= s282;

      elsif ( not x24 and x25 and x19 and not x14 and not x13 and not x26 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and x25 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and x26 and x18 and x14 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x24 and not x25 and x26 and x18 and not x14 and x13 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x24 and not x25 and x26 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and x26 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and not x26 and x10 and x12 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x24 and not x25 and not x26 and x10 and x12 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x24 and not x25 and not x26 and x10 and x12 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and not x26 and x10 and x12 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x24 and not x25 and not x26 and x10 and not x12 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x24 and not x25 and not x26 and not x10 and x17 and x14 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x24 and not x25 and not x26 and not x10 and x17 and not x14 and x13 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x24 and not x25 and not x26 and not x10 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s283 =>
      if ( x65 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s54;

      else
         y17 <= '1' ;
         current_group15m <= s77;

      end if;

   when s284 =>
      if ( x21 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x21 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x21 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      else
         y12 <= '1' ;
         current_group15m <= s100;

      end if;

   when s285 =>
      if ( x21 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x21 and x22 and x23 and x17 and not x14 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x21 and x22 and x23 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 and x18 and x14 ) = '1' then
         current_group15m <= s40;

      elsif ( not x21 and x22 and not x23 and x18 and not x14 and x13 ) = '1' then
         current_group15m <= s40;

      elsif ( not x21 and x22 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      else
         y4 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s180;

      end if;

   when s286 =>
      if ( x65 and x60 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s314;

      elsif ( x65 and not x60 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s356;

      elsif ( not x65 and x21 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x65 and x21 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x65 and x21 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and x23 and x10 and x12 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and not x21 and x22 and x23 and x10 and x12 and x17 and not x14 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and not x21 and x22 and x23 and x10 and x12 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and x23 and x10 and x12 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and x23 and x10 and not x12 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s341;

      elsif ( not x65 and not x21 and x22 and x23 and not x10 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and not x21 and x22 and x23 and not x10 and x17 and not x14 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x65 and not x21 and x22 and x23 and not x10 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and x23 and not x10 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and not x23 and x18 and x14 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x21 and x22 and not x23 and x18 and not x14 and x13 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and not x21 and x22 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      else
         y4 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s180;

      end if;

   when s287 =>
         y1 <= '1' ;
         y11 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s226;

   when s288 =>
      if ( x65 and x22 and x21 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x22 and x21 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x22 and x21 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x22 and x21 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x22 and not x21 and x18 and x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x22 and not x21 and x18 and not x19 and x10 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( x65 and x22 and not x21 and x18 and not x19 and not x10 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x22 and not x21 and x18 and not x19 and not x10 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x22 and not x21 and x18 and not x19 and not x10 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x22 and not x21 and x18 and not x19 and not x10 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x22 and not x21 and not x18 and x19 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x22 and not x21 and not x18 and x19 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x22 and not x21 and not x18 and x19 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x22 and not x21 and not x18 and not x19 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x22 and not x21 and not x18 and not x19 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x22 and not x21 and not x18 and not x19 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x22 and not x21 and not x18 and not x19 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x22 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x22 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and not x22 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x22 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x21 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x21 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x22 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and not x22 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and not x21 and not x22 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x65 and not x21 and not x22 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s289 =>
         y12 <= '1' ;
         current_group15m <= s210;

   when s290 =>
      if ( x65 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      else
         y17 <= '1' ;
         current_group15m <= s77;

      end if;

   when s291 =>
      if ( x65 and x60 ) = '1' then
         current_group15m <= s73;

      elsif ( x65 and not x60 and x61 ) = '1' then
         current_group15m <= s73;

      elsif ( x65 and not x60 and not x61 ) = '1' then
         current_group15m <= s40;

      else
         y17 <= '1' ;
         current_group15m <= s77;

      end if;

   when s292 =>
      if ( x65 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      else
         y17 <= '1' ;
         current_group15m <= s17;

      end if;

   when s293 =>
      if ( x66 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      else
         y12 <= '1' ;
         current_group15m <= s100;

      end if;

   when s294 =>
      if ( x21 ) = '1' then
         y35 <= '1' ;
         current_group15m <= s26;

      elsif ( not x21 and x23 and x22 ) = '1' then
         y20 <= '1' ;
         current_group15m <= s363;

      elsif ( not x21 and x23 and not x22 ) = '1' then
         y35 <= '1' ;
         current_group15m <= s26;

      elsif ( not x21 and not x23 and x22 and x17 and x15 and x9 ) = '1' then
         y4 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s119;

      elsif ( not x21 and not x23 and x22 and x17 and x15 and not x9 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( not x21 and not x23 and x22 and x17 and not x15 and x16 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( not x21 and not x23 and x22 and x17 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s205;

      elsif ( not x21 and not x23 and x22 and not x17 ) = '1' then
         y35 <= '1' ;
         current_group15m <= s26;

      elsif ( not x21 and not x23 and not x22 and x2 ) = '1' then
         y35 <= '1' ;
         current_group15m <= s26;

      elsif ( not x21 and not x23 and not x22 and not x2 and x17 and x15 and x9 ) = '1' then
         y6 <= '1' ;
         current_group15m <= s91;

      elsif ( not x21 and not x23 and not x22 and not x2 and x17 and x15 and not x9 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( not x21 and not x23 and not x22 and not x2 and x17 and not x15 and x16 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( not x21 and not x23 and not x22 and not x2 and x17 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s205;

      else
         y36 <= '1' ;
         current_group15m <= s55;

      end if;

   when s295 =>
         y9 <= '1' ;
         y10 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s240;

   when s296 =>
      if ( x66 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      else
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      end if;

   when s297 =>
      if ( x66 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x66 and x24 ) = '1' then
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s182;

      else
         y8 <= '1' ;
         current_group15m <= s92;

      end if;

   when s298 =>
      if ( x65 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s99;

      elsif ( not x65 and x63 and x1 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s156;

      elsif ( not x65 and x63 and not x1 and x18 and x15 and x8 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( not x65 and x63 and not x1 and x18 and x15 and not x8 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x65 and x63 and not x1 and x18 and not x15 and x16 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( not x65 and x63 and not x1 and x18 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s135;

      elsif ( not x65 and x63 and not x1 and not x18 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s152;

      else
         y3 <= '1' ;
         y22 <= '1' ;
         y37 <= '1' ;
         current_group15m <= s397;

      end if;

   when s299 =>
         y3 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s345;

   when s300 =>
      if ( x21 and x66 and x20 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x66 and x20 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x21 and x66 and x20 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x66 and x20 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x66 and not x20 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x21 and not x66 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x21 and not x66 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x21 and not x66 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x66 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x66 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x66 and x22 and x18 and x19 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x66 and x22 and x18 and x19 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x66 and x22 and x18 and x19 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x66 and x22 and x18 and not x19 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x66 and x22 and x18 and not x19 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x66 and x22 and x18 and not x19 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x66 and x22 and x18 and not x19 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x66 and x22 and not x18 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x66 and x22 and not x18 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x66 and x22 and not x18 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x66 and x22 and not x18 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x66 and not x22 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x66 and not x22 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x66 and not x22 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s301 =>
      if ( x65 and x21 and x20 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x21 and x20 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x21 and x20 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x21 and x20 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x21 and not x20 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x21 and not x20 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x21 and not x20 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x21 and not x20 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x21 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x65 and x19 ) = '1' then
         y4 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s304;

      elsif ( not x65 and not x19 and x20 and x15 and x10 and x11 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s334;

      elsif ( not x65 and not x19 and x20 and x15 and x10 and not x11 and x12 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s334;

      elsif ( not x65 and not x19 and x20 and x15 and x10 and not x11 and not x12 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x65 and not x19 and x20 and x15 and not x10 and x12 and x11 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      elsif ( not x65 and not x19 and x20 and x15 and not x10 and x12 and not x11 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x65 and not x19 and x20 and x15 and not x10 and not x12 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      elsif ( not x65 and not x19 and x20 and not x15 and x16 and x10 and x12 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and not x19 and x20 and not x15 and x16 and x10 and not x12 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s341;

      elsif ( not x65 and not x19 and x20 and not x15 and x16 and not x10 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and not x19 and x20 and not x15 and not x16 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s81;

      else
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      end if;

   when s302 =>
      if ( x65 and x67 and x22 and x17 and x18 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and x22 and x17 and not x18 and x19 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and x67 and x22 and x17 and not x18 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and x22 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x22 and x18 and x13 and x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and x67 and not x22 and x18 and x13 and not x23 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x67 and not x22 and x18 and not x13 and x12 and x23 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and x67 and not x22 and x18 and not x13 and x12 and not x23 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and x67 and not x22 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x22 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x21 and x20 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x67 and x21 and x20 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x67 and x21 and x20 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x21 and x20 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x21 and not x20 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and not x67 and x21 and not x20 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x65 and not x67 and x21 and not x20 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x21 and not x20 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and not x21 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s259;

      else
         y4 <= '1' ;
         y16 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s45;

      end if;

   when s303 =>
      if ( x20 and x21 and x17 and x14 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x20 and x21 and x17 and not x14 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x20 and x21 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x20 and x21 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( x20 and not x21 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      else
         y10 <= '1' ;
         current_group15m <= s12;

      end if;

   when s304 =>
      if ( x21 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x21 and x20 and x15 and x10 and x11 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s334;

      elsif ( not x21 and x20 and x15 and x10 and not x11 and x12 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s334;

      elsif ( not x21 and x20 and x15 and x10 and not x11 and not x12 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x21 and x20 and x15 and not x10 and x12 and x11 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      elsif ( not x21 and x20 and x15 and not x10 and x12 and not x11 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x21 and x20 and x15 and not x10 and not x12 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      elsif ( not x21 and x20 and not x15 and x16 and x10 and x12 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x21 and x20 and not x15 and x16 and x10 and not x12 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s341;

      elsif ( not x21 and x20 and not x15 and x16 and not x10 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x21 and x20 and not x15 and not x16 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s81;

      else
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      end if;

   when s305 =>
      if ( x68 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x68 and x21 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x68 and not x21 and x22 and x23 and x15 and x10 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( not x68 and not x21 and x22 and x23 and x15 and not x10 and x12 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x68 and not x21 and x22 and x23 and x15 and not x10 and not x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s285;

      elsif ( not x68 and not x21 and x22 and x23 and not x15 and x16 and x10 and x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( not x68 and not x21 and x22 and x23 and not x15 and x16 and x10 and not x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x68 and not x21 and x22 and x23 and not x15 and x16 and not x10 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( not x68 and not x21 and x22 and x23 and not x15 and not x16 ) = '1' then
         current_group15m <= s40;

      elsif ( not x68 and not x21 and x22 and not x23 and x6 and x15 and x11 and x10 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s334;

      elsif ( not x68 and not x21 and x22 and not x23 and x6 and x15 and x11 and not x10 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s285;

      elsif ( not x68 and not x21 and x22 and not x23 and x6 and x15 and not x11 and x12 and x10 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s334;

      elsif ( not x68 and not x21 and x22 and not x23 and x6 and x15 and not x11 and x12 and not x10 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x68 and not x21 and x22 and not x23 and x6 and x15 and not x11 and not x12 and x10 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( not x68 and not x21 and x22 and not x23 and x6 and x15 and not x11 and not x12 and not x10 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s285;

      elsif ( not x68 and not x21 and x22 and not x23 and x6 and not x15 and x16 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x68 and not x21 and x22 and not x23 and x6 and not x15 and not x16 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s180;

      elsif ( not x68 and not x21 and x22 and not x23 and not x6 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x68 and not x21 and not x22 and x23 and x15 and x7 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s81;

      elsif ( not x68 and not x21 and not x22 and x23 and x15 and not x7 and x9 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x68 and not x21 and not x22 and x23 and x15 and not x7 and not x9 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x68 and not x21 and not x22 and x23 and not x15 and x16 and x7 and x9 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x68 and not x21 and not x22 and x23 and not x15 and x16 and x7 and not x9 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( not x68 and not x21 and not x22 and x23 and not x15 and x16 and not x7 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x68 and not x21 and not x22 and x23 and not x15 and not x16 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      else
         y3 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s81;

      end if;

   when s306 =>
      if ( x21 and x20 and x18 and x15 and x10 and x11 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s192;

      elsif ( x21 and x20 and x18 and x15 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s193;

      elsif ( x21 and x20 and x18 and x15 and x10 and not x11 and not x12 ) = '1' then
         y1 <= '1' ;
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s194;

      elsif ( x21 and x20 and x18 and x15 and not x10 and x12 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s300;

      elsif ( x21 and x20 and x18 and x15 and not x10 and not x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s192;

      elsif ( x21 and x20 and x18 and not x15 and x16 and x10 and x12 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s259;

      elsif ( x21 and x20 and x18 and not x15 and x16 and x10 and not x12 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( x21 and x20 and x18 and not x15 and x16 and not x10 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s259;

      elsif ( x21 and x20 and x18 and not x15 and not x16 ) = '1' then
         y2 <= '1' ;
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s134;

      elsif ( x21 and x20 and not x18 ) = '1' then
         y4 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s307;

      elsif ( x21 and not x20 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s199;

      elsif ( not x21 and x18 and x15 and x10 and x11 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x21 and x18 and x15 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s301;

      elsif ( not x21 and x18 and x15 and x10 and not x11 and not x12 ) = '1' then
         y8 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s195;

      elsif ( not x21 and x18 and x15 and not x10 and x12 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s197;

      elsif ( not x21 and x18 and x15 and not x10 and not x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s192;

      elsif ( not x21 and x18 and not x15 and x16 and x10 and x12 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s259;

      elsif ( not x21 and x18 and not x15 and x16 and x10 and not x12 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s302;

      elsif ( not x21 and x18 and not x15 and x16 and not x10 ) = '1' then
         y1 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s259;

      elsif ( not x21 and x18 and not x15 and not x16 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s303;

      else
         y5 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s57;

      end if;

   when s307 =>
      if ( x21 ) = '1' then
         y2 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s121;

      else
         current_group15m <= s1;

      end if;

   when s308 =>
         y2 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s79;

   when s309 =>
      if ( x22 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      else
         y17 <= '1' ;
         current_group15m <= s17;

      end if;

   when s310 =>
      if ( x21 and x9 and x8 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x21 and x9 and not x8 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( x21 and x9 and not x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x8 and x7 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( not x21 and x22 and x8 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x4 and x5 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x21 and not x22 and x4 and not x5 and x6 ) = '1' then
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s29;

      elsif ( not x21 and not x22 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s311 =>
      if ( x21 and x16 and x15 and x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s214;

      elsif ( x21 and x16 and x15 and not x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s215;

      elsif ( x21 and x16 and not x15 and x10 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s114;

      elsif ( x21 and x16 and not x15 and not x10 ) = '1' then
         y14 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s216;

      elsif ( x21 and not x16 and x17 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s215;

      elsif ( x21 and not x16 and not x17 and x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s215;

      elsif ( x21 and not x16 and not x17 and not x10 ) = '1' then
         y11 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s218;

      else
         y17 <= '1' ;
         current_group15m <= s77;

      end if;

   when s312 =>
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s118;

   when s313 =>
         y8 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s267;

   when s314 =>
      if ( x67 and x22 and x15 and x8 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x67 and x22 and x15 and not x8 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x67 and x22 and not x15 and x16 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s302;

      elsif ( x67 and x22 and not x15 and not x16 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s122;

      elsif ( x67 and not x22 ) = '1' then
         y10 <= '1' ;
         y26 <= '1' ;
         y27 <= '1' ;
         current_group15m <= s2;

      elsif ( not x67 and x60 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s154;

      else
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      end if;

   when s315 =>
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

   when s316 =>
      if ( x60 ) = '1' then
         current_group15m <= s1;

      elsif ( not x60 and x61 ) = '1' then
         current_group15m <= s1;

      elsif ( not x60 and not x61 and x62 ) = '1' then
         y2 <= '1' ;
         y19 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s321;

      else
         current_group15m <= s40;

      end if;

   when s317 =>
      if ( x21 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s75;

      elsif ( not x21 and x16 and x10 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s67;

      elsif ( not x21 and x16 and not x10 ) = '1' then
         y5 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s113;

      elsif ( not x21 and not x16 and x17 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      else
         y5 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s115;

      end if;

   when s318 =>
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

   when s319 =>
      if ( x65 and x61 and x60 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s328;

      elsif ( x65 and x61 and not x60 and x62 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      elsif ( x65 and x61 and not x60 and not x62 and x2 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s255;

      elsif ( x65 and x61 and not x60 and not x62 and not x2 and x19 and x15 ) = '1' then
         current_group15m <= s73;

      elsif ( x65 and x61 and not x60 and not x62 and not x2 and x19 and not x15 and x16 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s291;

      elsif ( x65 and x61 and not x60 and not x62 and not x2 and x19 and not x15 and not x16 ) = '1' then
         current_group15m <= s73;

      elsif ( x65 and x61 and not x60 and not x62 and not x2 and not x19 ) = '1' then
         y4 <= '1' ;
         y13 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s64;

      elsif ( x65 and not x61 and x60 and x2 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s255;

      elsif ( x65 and not x61 and x60 and not x2 and x19 and x15 ) = '1' then
         current_group15m <= s73;

      elsif ( x65 and not x61 and x60 and not x2 and x19 and not x15 and x16 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s291;

      elsif ( x65 and not x61 and x60 and not x2 and x19 and not x15 and not x16 ) = '1' then
         current_group15m <= s73;

      elsif ( x65 and not x61 and x60 and not x2 and not x19 ) = '1' then
         y4 <= '1' ;
         y13 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s64;

      elsif ( x65 and not x61 and not x60 and x62 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and not x61 and not x60 and not x62 and x5 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s255;

      elsif ( x65 and not x61 and not x60 and not x62 and not x5 and x18 and x15 and x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x65 and not x61 and not x60 and not x62 and not x5 and x18 and x15 and not x7 and x11 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x65 and not x61 and not x60 and not x62 and not x5 and x18 and x15 and not x7 and not x11 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s254;

      elsif ( x65 and not x61 and not x60 and not x62 and not x5 and x18 and not x15 and x16 and x4 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and not x61 and not x60 and not x62 and not x5 and x18 and not x15 and x16 and not x4 and x11 and x9 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and not x61 and not x60 and not x62 and not x5 and x18 and not x15 and x16 and not x4 and x11 and not x9 and x7 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s128;

      elsif ( x65 and not x61 and not x60 and not x62 and not x5 and x18 and not x15 and x16 and not x4 and x11 and not x9 and not x7 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s118;

      elsif ( x65 and not x61 and not x60 and not x62 and not x5 and x18 and not x15 and x16 and not x4 and not x11 and x9 and x7 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x65 and not x61 and not x60 and not x62 and not x5 and x18 and not x15 and x16 and not x4 and not x11 and x9 and not x7 and x10 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x65 and not x61 and not x60 and not x62 and not x5 and x18 and not x15 and x16 and not x4 and not x11 and x9 and not x7 and not x10 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and not x61 and not x60 and not x62 and not x5 and x18 and not x15 and x16 and not x4 and not x11 and not x9 and x7 and x8 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x65 and not x61 and not x60 and not x62 and not x5 and x18 and not x15 and x16 and not x4 and not x11 and not x9 and x7 and not x8 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and not x61 and not x60 and not x62 and not x5 and x18 and not x15 and x16 and not x4 and not x11 and not x9 and not x7 and x12 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x65 and not x61 and not x60 and not x62 and not x5 and x18 and not x15 and x16 and not x4 and not x11 and not x9 and not x7 and not x12 ) = '1' then
         current_group15m <= s40;

      elsif ( x65 and not x61 and not x60 and not x62 and not x5 and x18 and not x15 and not x16 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( x65 and not x61 and not x60 and not x62 and not x5 and not x18 ) = '1' then
         y4 <= '1' ;
         y13 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s64;

      else
         y2 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s374;

      end if;

   when s320 =>
      if ( x65 ) = '1' then
         current_group15m <= s40;

      elsif ( not x65 and x66 and x23 and x18 and x15 and x7 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y9 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s81;

      elsif ( not x65 and x66 and x23 and x18 and x15 and not x7 and x9 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x65 and x66 and x23 and x18 and x15 and not x7 and not x9 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x65 and x66 and x23 and x18 and not x15 and x7 and x9 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s330;

      elsif ( not x65 and x66 and x23 and x18 and not x15 and x7 and not x9 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( not x65 and x66 and x23 and x18 and not x15 and not x7 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s330;

      elsif ( not x65 and x66 and x23 and not x18 ) = '1' then
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s84;

      elsif ( not x65 and x66 and not x23 and x9 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x65 and x66 and not x23 and not x9 and x7 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x65 and x66 and not x23 and not x9 and not x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      else
         y5 <= '1' ;
         current_group15m <= s343;

      end if;

   when s321 =>
      if ( x61 and x16 and x17 and x11 and x13 ) = '1' then
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s260;

      elsif ( x61 and x16 and x17 and x11 and not x13 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         y10 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s261;

      elsif ( x61 and x16 and x17 and not x11 and x12 and x13 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s262;

      elsif ( x61 and x16 and x17 and not x11 and x12 and not x13 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s254;

      elsif ( x61 and x16 and x17 and not x11 and not x12 and x13 and x15 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s355;

      elsif ( x61 and x16 and x17 and not x11 and not x12 and x13 and not x15 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x61 and x16 and x17 and not x11 and not x12 and x13 and not x15 and x18 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x61 and x16 and x17 and not x11 and not x12 and x13 and not x15 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x61 and x16 and x17 and not x11 and not x12 and not x13 and x14 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s355;

      elsif ( x61 and x16 and x17 and not x11 and not x12 and not x13 and not x14 and x18 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x61 and x16 and x17 and not x11 and not x12 and not x13 and not x14 and x18 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x61 and x16 and x17 and not x11 and not x12 and not x13 and not x14 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x61 and x16 and not x17 and x12 and x11 and x13 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( x61 and x16 and not x17 and x12 and x11 and x13 and not x3 and x2 ) = '1' then
         current_group15m <= s40;

      elsif ( x61 and x16 and not x17 and x12 and x11 and x13 and not x3 and not x2 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s224;

      elsif ( x61 and x16 and not x17 and x12 and x11 and not x13 ) = '1' then
         y3 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s255;

      elsif ( x61 and x16 and not x17 and x12 and not x11 and x13 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s7;

      elsif ( x61 and x16 and not x17 and x12 and not x11 and not x13 ) = '1' then
         y2 <= '1' ;
         y10 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s263;

      elsif ( x61 and x16 and not x17 and not x12 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( x61 and x16 and not x17 and not x12 and not x3 and x2 ) = '1' then
         current_group15m <= s40;

      elsif ( x61 and x16 and not x17 and not x12 and not x3 and not x2 and x13 and x11 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s58;

      elsif ( x61 and x16 and not x17 and not x12 and not x3 and not x2 and x13 and not x11 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x61 and x16 and not x17 and not x12 and not x3 and not x2 and not x13 and x11 ) = '1' then
         y4 <= '1' ;
         y13 <= '1' ;
         y24 <= '1' ;
         current_group15m <= s64;

      elsif ( x61 and x16 and not x17 and not x12 and not x3 and not x2 and not x13 and not x11 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x61 and not x16 and x3 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( x61 and not x16 and not x3 and x17 and x13 and x11 and x9 and x2 ) = '1' then
         current_group15m <= s40;

      elsif ( x61 and not x16 and not x3 and x17 and x13 and x11 and x9 and not x2 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s252;

      elsif ( x61 and not x16 and not x3 and x17 and x13 and x11 and not x9 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x61 and not x16 and not x3 and x17 and x13 and x11 and not x9 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x61 and not x16 and not x3 and x17 and x13 and x11 and not x9 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x61 and not x16 and not x3 and x17 and x13 and x11 and not x9 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x61 and not x16 and not x3 and x17 and x13 and not x11 and x12 and x2 ) = '1' then
         current_group15m <= s40;

      elsif ( x61 and not x16 and not x3 and x17 and x13 and not x11 and x12 and not x2 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s252;

      elsif ( x61 and not x16 and not x3 and x17 and x13 and not x11 and not x12 and x8 and x2 ) = '1' then
         current_group15m <= s40;

      elsif ( x61 and not x16 and not x3 and x17 and x13 and not x11 and not x12 and x8 and not x2 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s252;

      elsif ( x61 and not x16 and not x3 and x17 and x13 and not x11 and not x12 and not x8 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x61 and not x16 and not x3 and x17 and x13 and not x11 and not x12 and not x8 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x61 and not x16 and not x3 and x17 and x13 and not x11 and not x12 and not x8 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x61 and not x16 and not x3 and x17 and x13 and not x11 and not x12 and not x8 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x61 and not x16 and not x3 and x17 and not x13 and x11 ) = '1' then
         current_group15m <= s40;

      elsif ( x61 and not x16 and not x3 and x17 and not x13 and not x11 and x12 and x10 and x2 ) = '1' then
         current_group15m <= s40;

      elsif ( x61 and not x16 and not x3 and x17 and not x13 and not x11 and x12 and x10 and not x2 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s252;

      elsif ( x61 and not x16 and not x3 and x17 and not x13 and not x11 and x12 and not x10 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x61 and not x16 and not x3 and x17 and not x13 and not x11 and x12 and not x10 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x61 and not x16 and not x3 and x17 and not x13 and not x11 and x12 and not x10 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x61 and not x16 and not x3 and x17 and not x13 and not x11 and x12 and not x10 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x61 and not x16 and not x3 and x17 and not x13 and not x11 and not x12 and x7 and x2 ) = '1' then
         current_group15m <= s40;

      elsif ( x61 and not x16 and not x3 and x17 and not x13 and not x11 and not x12 and x7 and not x2 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s252;

      elsif ( x61 and not x16 and not x3 and x17 and not x13 and not x11 and not x12 and not x7 and x18 and x14 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x61 and not x16 and not x3 and x17 and not x13 and not x11 and not x12 and not x7 and x18 and not x14 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x61 and not x16 and not x3 and x17 and not x13 and not x11 and not x12 and not x7 and x18 and not x14 and not x15 ) = '1' then
         current_group15m <= s1;

      elsif ( x61 and not x16 and not x3 and x17 and not x13 and not x11 and not x12 and not x7 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( x61 and not x16 and not x3 and not x17 and x2 ) = '1' then
         current_group15m <= s40;

      elsif ( x61 and not x16 and not x3 and not x17 and not x2 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s74;

      elsif ( not x61 and x62 and x2 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         y10 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s261;

      elsif ( not x61 and x62 and not x2 and x19 and x15 and x12 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s292;

      elsif ( not x61 and x62 and not x2 and x19 and x15 and x12 and not x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s290;

      elsif ( not x61 and x62 and not x2 and x19 and x15 and not x12 and x7 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s63;

      elsif ( not x61 and x62 and not x2 and x19 and x15 and not x12 and not x7 ) = '1' then
         y2 <= '1' ;
         y10 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s263;

      elsif ( not x61 and x62 and not x2 and x19 and not x15 and x16 and x7 and x12 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s290;

      elsif ( not x61 and x62 and not x2 and x19 and not x15 and x16 and x7 and not x12 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s262;

      elsif ( not x61 and x62 and not x2 and x19 and not x15 and x16 and not x7 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s258;

      elsif ( not x61 and x62 and not x2 and x19 and not x15 and not x16 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x61 and x62 and not x2 and x19 and not x15 and not x16 and not x7 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x61 and x62 and not x2 and not x19 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s411;

      else
         current_group15m <= s1;

      end if;

   when s322 =>
         y5 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s262;

   when s323 =>
      if ( x3 and x4 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( x3 and not x4 and x5 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( x3 and not x4 and not x5 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s324 =>
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s414;

   when s325 =>
         current_group15m <= s40;

   when s326 =>
         y3 <= '1' ;
         current_group15m <= s89;

   when s327 =>
         y19 <= '1' ;
         current_group15m <= s11;

   when s328 =>
      if ( x65 and x60 and x61 ) = '1' then
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s38;

      elsif ( x65 and x60 and not x61 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s68;

      elsif ( x65 and not x60 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s68;

      elsif ( not x65 and x68 and x19 ) = '1' then
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s375;

      elsif ( not x65 and x68 and not x19 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x65 and not x68 and x21 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      else
         y8 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s378;

      end if;

   when s329 =>
      if ( x65 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s66;

      else
         y9 <= '1' ;
         current_group15m <= s27;

      end if;

   when s330 =>
      if ( x21 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x21 and x22 and x23 and x17 and not x14 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x21 and x22 and x23 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 and x18 and x14 ) = '1' then
         current_group15m <= s40;

      elsif ( not x21 and x22 and not x23 and x18 and not x14 and x13 ) = '1' then
         current_group15m <= s40;

      elsif ( not x21 and x22 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and x7 and x9 and x19 and x14 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x21 and not x22 and x23 and x7 and x9 and x19 and not x14 and x13 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x21 and not x22 and x23 and x7 and x9 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and x7 and x9 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and x7 and not x9 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s333;

      elsif ( not x21 and not x22 and x23 and not x7 and x19 and x14 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x21 and not x22 and x23 and not x7 and x19 and not x14 and x13 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x21 and not x22 and x23 and not x7 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and not x7 and not x19 ) = '1' then
         current_group15m <= s1;

      else
         y12 <= '1' ;
         current_group15m <= s100;

      end if;

   when s331 =>
      if ( x21 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 and x18 and x14 ) = '1' then
         current_group15m <= s40;

      elsif ( not x21 and x22 and not x23 and x18 and not x14 and x13 ) = '1' then
         current_group15m <= s40;

      elsif ( not x21 and x22 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and x19 and x14 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x21 and not x22 and x23 and x19 and not x14 and x13 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x21 and not x22 and x23 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and not x19 ) = '1' then
         current_group15m <= s1;

      else
         y12 <= '1' ;
         current_group15m <= s100;

      end if;

   when s332 =>
      if ( x21 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x23 and x22 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x21 and x23 and not x22 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s180;

      else
         y12 <= '1' ;
         current_group15m <= s100;

      end if;

   when s333 =>
      if ( x21 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s143;

      elsif ( not x21 and x22 and x23 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x21 and x22 and x23 and x17 and not x14 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x21 and x22 and x23 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x21 and not x22 and x23 and x19 and x14 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x21 and not x22 and x23 and x19 and not x14 and x13 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x21 and not x22 and x23 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and not x19 ) = '1' then
         current_group15m <= s1;

      else
         y3 <= '1' ;
         current_group15m <= s320;

      end if;

   when s334 =>
         y12 <= '1' ;
         current_group15m <= s100;

   when s335 =>
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s341;

   when s336 =>
      if ( x68 and x7 and x8 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( x68 and x7 and not x8 and x9 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( x68 and x7 and not x8 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x68 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x68 and x21 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s343;

      elsif ( not x68 and not x21 and x22 and x23 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x68 and not x21 and x22 and x23 and x17 and not x14 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x68 and not x21 and x22 and x23 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x68 and not x21 and x22 and x23 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x68 and not x21 and x22 and not x23 and x18 and x14 ) = '1' then
         current_group15m <= s40;

      elsif ( not x68 and not x21 and x22 and not x23 and x18 and not x14 and x13 ) = '1' then
         current_group15m <= s40;

      elsif ( not x68 and not x21 and x22 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x68 and not x21 and x22 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x68 and not x21 and not x22 and x23 ) = '1' then
         current_group15m <= s1;

      else
         y4 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s180;

      end if;

   when s337 =>
      if ( x23 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s333;

      else
         y3 <= '1' ;
         current_group15m <= s89;

      end if;

   when s338 =>
      if ( x65 and x66 ) = '1' then
         current_group15m <= s316;

      elsif ( x65 and not x66 and x67 and x8 and x9 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x65 and not x66 and x67 and x8 and not x9 and x10 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s136;

      elsif ( x65 and not x66 and x67 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and x67 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x19 and x18 and x14 ) = '1' then
         y6 <= '1' ;
         y8 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x19 and x18 and not x14 and x17 ) = '1' then
         y6 <= '1' ;
         y8 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x19 and x18 and not x14 and not x17 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x19 and x18 and not x14 and not x17 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and x19 and x18 and not x14 and not x17 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x19 and x18 and not x14 and not x17 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and x19 and not x18 ) = '1' then
         y6 <= '1' ;
         y8 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and not x19 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and not x19 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and not x66 and not x67 and not x19 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x66 and not x67 and not x19 and not x5 ) = '1' then
         current_group15m <= s1;

      else
         y7 <= '1' ;
         current_group15m <= s140;

      end if;

   when s339 =>
      if ( x21 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( x21 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and x4 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s53;

      elsif ( not x21 and x22 and x23 and not x4 and x18 and x15 and x10 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      elsif ( not x21 and x22 and x23 and not x4 and x18 and x15 and not x10 and x12 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x21 and x22 and x23 and not x4 and x18 and x15 and not x10 and not x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s285;

      elsif ( not x21 and x22 and x23 and not x4 and x18 and not x15 and x16 and x10 and x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s286;

      elsif ( not x21 and x22 and x23 and not x4 and x18 and not x15 and x16 and x10 and not x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x21 and x22 and x23 and not x4 and x18 and not x15 and x16 and not x10 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s286;

      elsif ( not x21 and x22 and x23 and not x4 and x18 and not x15 and not x16 ) = '1' then
         current_group15m <= s40;

      elsif ( not x21 and x22 and x23 and not x4 and not x18 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x21 and x22 and not x23 and x18 and x14 ) = '1' then
         current_group15m <= s40;

      elsif ( not x21 and x22 and not x23 and x18 and not x14 and x13 ) = '1' then
         current_group15m <= s40;

      elsif ( not x21 and x22 and not x23 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and x19 and x14 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x21 and not x22 and x23 and x19 and not x14 and x13 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x21 and not x22 and x23 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and not x19 ) = '1' then
         current_group15m <= s1;

      else
         y12 <= '1' ;
         current_group15m <= s100;

      end if;

   when s340 =>
      if ( x21 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      elsif ( not x21 and x22 and x15 and x10 and x16 and x12 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x21 and x22 and x15 and x10 and x16 and not x12 ) = '1' then
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s339;

      elsif ( not x21 and x22 and x15 and x10 and not x16 and x3 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x21 and x22 and x15 and x10 and not x16 and not x3 and x2 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( not x21 and x22 and x15 and x10 and not x16 and not x3 and not x2 and x11 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s126;

      elsif ( not x21 and x22 and x15 and x10 and not x16 and not x3 and not x2 and not x11 and x12 ) = '1' then
         y3 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s332;

      elsif ( not x21 and x22 and x15 and x10 and not x16 and not x3 and not x2 and not x11 and not x12 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s330;

      elsif ( not x21 and x22 and x15 and not x10 and x11 and x12 and x16 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s331;

      elsif ( not x21 and x22 and x15 and not x10 and x11 and x12 and not x16 and x3 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x21 and x22 and x15 and not x10 and x11 and x12 and not x16 and not x3 and x2 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( not x21 and x22 and x15 and not x10 and x11 and x12 and not x16 and not x3 and not x2 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s336;

      elsif ( not x21 and x22 and x15 and not x10 and x11 and not x12 and x16 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and x15 and not x10 and x11 and not x12 and not x16 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s333;

      elsif ( not x21 and x22 and x15 and not x10 and not x11 and x16 and x12 and x13 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s122;

      elsif ( not x21 and x22 and x15 and not x10 and not x11 and x16 and x12 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x15 and not x10 and not x11 and x16 and not x12 and x14 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s122;

      elsif ( not x21 and x22 and x15 and not x10 and not x11 and x16 and not x12 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x15 and not x10 and not x11 and not x16 and x3 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x21 and x22 and x15 and not x10 and not x11 and not x16 and not x3 and x2 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( not x21 and x22 and x15 and not x10 and not x11 and not x16 and not x3 and not x2 and x12 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x21 and x22 and x15 and not x10 and not x11 and not x16 and not x3 and not x2 and not x12 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s48;

      elsif ( not x21 and x22 and not x15 and x16 and x12 and x10 and x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x15 and x16 and x12 and x10 and not x8 and x3 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x21 and x22 and not x15 and x16 and x12 and x10 and not x8 and not x3 and x2 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( not x21 and x22 and not x15 and x16 and x12 and x10 and not x8 and not x3 and not x2 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( not x21 and x22 and not x15 and x16 and x12 and not x10 and x11 and x3 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x21 and x22 and not x15 and x16 and x12 and not x10 and x11 and not x3 and x2 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( not x21 and x22 and not x15 and x16 and x12 and not x10 and x11 and not x3 and not x2 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( not x21 and x22 and not x15 and x16 and x12 and not x10 and not x11 and x7 and x3 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x21 and x22 and not x15 and x16 and x12 and not x10 and not x11 and x7 and not x3 and x2 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s69;

      elsif ( not x21 and x22 and not x15 and x16 and x12 and not x10 and not x11 and x7 and not x3 and not x2 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( not x21 and x22 and not x15 and x16 and x12 and not x10 and not x11 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x15 and x16 and not x12 and x10 and x3 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x21 and x22 and not x15 and x16 and not x12 and x10 and not x3 and x2 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s264;

      elsif ( not x21 and x22 and not x15 and x16 and not x12 and x10 and not x3 and not x2 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( not x21 and x22 and not x15 and x16 and not x12 and not x10 and x11 and x9 and x3 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x21 and x22 and not x15 and x16 and not x12 and not x10 and x11 and x9 and not x3 and x2 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( not x21 and x22 and not x15 and x16 and not x12 and not x10 and x11 and x9 and not x3 and not x2 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( not x21 and x22 and not x15 and x16 and not x12 and not x10 and x11 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x15 and x16 and not x12 and not x10 and not x11 and x8 and x3 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x21 and x22 and not x15 and x16 and not x12 and not x10 and not x11 and x8 and not x3 and x2 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( not x21 and x22 and not x15 and x16 and not x12 and not x10 and not x11 and x8 and not x3 and not x2 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( not x21 and x22 and not x15 and x16 and not x12 and not x10 and not x11 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x15 and not x16 and x3 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x21 and x22 and not x15 and not x16 and not x3 and x2 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      elsif ( not x21 and x22 and not x15 and not x16 and not x3 and not x2 ) = '1' then
         y7 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s110;

      elsif ( not x21 and not x22 and x23 and x19 and x14 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x21 and not x22 and x23 and x19 and not x14 and x13 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x21 and not x22 and x23 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x23 and not x19 ) = '1' then
         current_group15m <= s1;

      else
         y12 <= '1' ;
         current_group15m <= s100;

      end if;

   when s341 =>
      if ( x68 and x7 and x8 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( x68 and x7 and not x8 and x9 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      elsif ( x68 and x7 and not x8 and not x9 ) = '1' then
         current_group15m <= s1;

      elsif ( x68 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( not x68 and x21 and x18 and x14 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x68 and x21 and x18 and not x14 and x13 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s144;

      elsif ( not x68 and x21 and x18 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x68 and x21 and not x18 ) = '1' then
         current_group15m <= s1;

      elsif ( not x68 and not x21 and x22 and x23 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x68 and not x21 and x22 and x23 and x17 and not x14 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x68 and not x21 and x22 and x23 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x68 and not x21 and x22 and x23 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x68 and not x21 and x22 and not x23 ) = '1' then
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s301;

      elsif ( not x68 and not x21 and not x22 and x23 and x19 and x14 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x68 and not x21 and not x22 and x23 and x19 and not x14 and x13 ) = '1' then
         y7 <= '1' ;
         y10 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s145;

      elsif ( not x68 and not x21 and not x22 and x23 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x68 and not x21 and not x22 and x23 and not x19 ) = '1' then
         current_group15m <= s1;

      else
         y4 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s180;

      end if;

   when s342 =>
      if ( x66 and x22 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s122;

      elsif ( x66 and not x22 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      else
         y1 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s142;

      end if;

   when s343 =>
      if ( x66 and x21 ) = '1' then
         y1 <= '1' ;
         current_group15m <= s22;

      elsif ( x66 and not x21 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s86;

      else
         y10 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s273;

      end if;

   when s344 =>
      if ( x21 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      elsif ( not x21 and x20 and x15 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( not x21 and x20 and not x15 and x14 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( not x21 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s345 =>
      if ( x68 and x15 and x10 and x11 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s192;

      elsif ( x68 and x15 and x10 and not x11 and x12 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s193;

      elsif ( x68 and x15 and x10 and not x11 and not x12 ) = '1' then
         y1 <= '1' ;
         y8 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s192;

      elsif ( x68 and x15 and not x10 and x12 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s300;

      elsif ( x68 and x15 and not x10 and not x12 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s192;

      elsif ( x68 and not x15 and x16 and x10 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x68 and not x15 and x16 and x10 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x68 and not x15 and x16 and x10 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x68 and not x15 and x16 and x10 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x68 and not x15 and x16 and not x10 and x12 and x11 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s199;

      elsif ( x68 and not x15 and x16 and not x10 and x12 and not x11 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x68 and not x15 and x16 and not x10 and x12 and not x11 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x68 and not x15 and x16 and not x10 and x12 and not x11 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x68 and not x15 and x16 and not x10 and x12 and not x11 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x68 and not x15 and x16 and not x10 and not x12 and x19 and x14 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x68 and not x15 and x16 and not x10 and not x12 and x19 and not x14 and x13 ) = '1' then
         y22 <= '1' ;
         current_group15m <= s4;

      elsif ( x68 and not x15 and x16 and not x10 and not x12 and x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( x68 and not x15 and x16 and not x10 and not x12 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x68 and not x15 and not x16 ) = '1' then
         y5 <= '1' ;
         y7 <= '1' ;
         y8 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s201;

      else
         y1 <= '1' ;
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s72;

      end if;

   when s346 =>
      if ( x67 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x67 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x67 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x67 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x67 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x67 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x67 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s347 =>
      if ( x19 and x20 and x11 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x19 and x20 and not x11 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x19 and x20 and not x11 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x19 and x20 and not x11 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x19 and x20 and not x11 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( x19 and not x20 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x19 and not x20 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x19 and not x20 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x19 and not x20 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x19 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x19 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x19 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s348 =>
      if ( x19 and x17 and x20 and x14 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( x19 and x17 and x20 and not x14 ) = '1' then
         y4 <= '1' ;
         y29 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s351;

      elsif ( x19 and x17 and not x20 and x14 ) = '1' then
         y4 <= '1' ;
         y18 <= '1' ;
         y29 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s351;

      elsif ( x19 and x17 and not x20 and not x14 and x15 ) = '1' then
         y16 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s352;

      elsif ( x19 and x17 and not x20 and not x14 and not x15 and x16 ) = '1' then
         y29 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s351;

      elsif ( x19 and x17 and not x20 and not x14 and not x15 and not x16 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s351;

      elsif ( x19 and not x17 and x18 ) = '1' then
         y2 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s349;

      elsif ( x19 and not x17 and not x18 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( not x19 and x20 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( not x19 and not x20 and x17 and x16 ) = '1' then
         y29 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s351;

      elsif ( not x19 and not x20 and x17 and not x16 and x15 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x19 and not x20 and x17 and not x16 and not x15 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( not x19 and not x20 and not x17 and x18 and x4 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s415;

      elsif ( not x19 and not x20 and not x17 and x18 and not x4 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s338;

      else
         y4 <= '1' ;
         current_group15m <= s43;

      end if;

   when s349 =>
      if ( x19 and x11 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x19 and not x11 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x19 and not x11 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x19 and not x11 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x19 and not x11 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x19 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x19 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x19 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s350 =>
      if ( x19 and x14 and x20 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s338;

      elsif ( x19 and x14 and not x20 ) = '1' then
         y2 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s416;

      elsif ( x19 and not x14 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s338;

      elsif ( not x19 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x19 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x19 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s351 =>
      if ( x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s352 =>
      if ( x19 and x20 and x9 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s415;

      elsif ( x19 and x20 and not x9 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( x19 and not x20 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x19 and not x20 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x19 and not x20 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x19 and not x20 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x19 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x19 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x19 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s353 =>
      if ( x65 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 ) = '1' then
         y17 <= '1' ;
         current_group15m <= s77;

      else
         y4 <= '1' ;
         y5 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s344;

      end if;

   when s354 =>
         y14 <= '1' ;
         current_group15m <= s417;

   when s355 =>
      if ( x65 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      else
         y15 <= '1' ;
         y112 <= '1' ;
         current_group15m <= s46;

      end if;

   when s356 =>
      if ( x65 and x60 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s63;

      elsif ( x65 and not x60 and x61 and x62 ) = '1' then
         y1 <= '1' ;
         y4 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s411;

      elsif ( x65 and not x60 and x61 and not x62 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s63;

      elsif ( x65 and not x60 and not x61 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      else
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      end if;

   when s357 =>
      if ( x65 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      else
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      end if;

   when s358 =>
      if ( x21 and x18 and x10 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x21 and x18 and not x10 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x21 and x18 and not x10 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x21 and x18 and not x10 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x18 and not x10 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x21 and not x18 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x21 and not x18 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and x22 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and x22 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x20 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x22 and x20 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x22 and x20 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x20 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x20 and x19 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x22 and not x20 and x19 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x22 and not x20 and x19 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x20 and x19 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x20 and not x19 and x10 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( not x21 and not x22 and not x20 and not x19 and not x10 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x22 and not x20 and not x19 and not x10 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x22 and not x20 and not x19 and not x10 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s359 =>
      if ( x21 and x16 and x13 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x21 and x16 and not x13 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s360;

      elsif ( x21 and not x16 and x17 and x18 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s418;

      elsif ( x21 and not x16 and x17 and x18 and not x3 and x13 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s249;

      elsif ( x21 and not x16 and x17 and x18 and not x3 and not x13 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( x21 and not x16 and x17 and not x18 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( x21 and not x16 and not x17 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s146;

      elsif ( not x21 and x22 and x16 and x19 and x18 and x10 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x21 and x22 and x16 and x19 and x18 and not x10 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s362;

      elsif ( not x21 and x22 and x16 and x19 and not x18 and x13 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and x16 and x19 and not x18 and not x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x21 and x22 and x16 and not x19 and x13 ) = '1' then
         y3 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s146;

      elsif ( not x21 and x22 and x16 and not x19 and not x13 and x18 and x15 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and x16 and not x19 and not x13 and x18 and not x15 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( not x21 and x22 and x16 and not x19 and not x13 and not x18 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x21 and x22 and not x16 and x17 and x18 and x19 and x10 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s418;

      elsif ( not x21 and x22 and not x16 and x17 and x18 and x19 and x10 and not x3 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

      elsif ( not x21 and x22 and not x16 and x17 and x18 and x19 and not x10 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s146;

      elsif ( not x21 and x22 and not x16 and x17 and x18 and not x19 and x13 and x3 ) = '1' then
         y3 <= '1' ;
         y8 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s419;

      elsif ( not x21 and x22 and not x16 and x17 and x18 and not x19 and x13 and not x3 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

      elsif ( not x21 and x22 and not x16 and x17 and x18 and not x19 and not x13 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x21 and x22 and not x16 and x17 and not x18 and x13 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s418;

      elsif ( not x21 and x22 and not x16 and x17 and not x18 and x13 and not x3 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

      elsif ( not x21 and x22 and not x16 and x17 and not x18 and not x13 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( not x21 and x22 and not x16 and x17 and not x18 and not x13 and not x19 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( not x21 and x22 and not x16 and not x17 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s146;

      elsif ( not x21 and not x22 and x19 and x17 and x13 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and not x22 and x19 and x17 and not x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x21 and not x22 and x19 and not x17 and x18 and x13 and x3 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

      elsif ( not x21 and not x22 and x19 and not x17 and x18 and x13 and not x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s418;

      elsif ( not x21 and not x22 and x19 and not x17 and x18 and not x13 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( not x21 and not x22 and x19 and not x17 and not x18 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s146;

      elsif ( not x21 and not x22 and not x19 and x16 and x13 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( not x21 and not x22 and not x19 and x16 and not x13 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s360;

      elsif ( not x21 and not x22 and not x19 and not x16 and x17 and x20 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( not x21 and not x22 and not x19 and not x16 and x17 and not x20 and x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s418;

      elsif ( not x21 and not x22 and not x19 and not x16 and x17 and not x20 and not x3 and x13 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s249;

      elsif ( not x21 and not x22 and not x19 and not x16 and x17 and not x20 and not x3 and not x13 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      else
         y8 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s146;

      end if;

   when s360 =>
      if ( x21 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x21 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x21 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x19 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and x22 and x19 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and x22 and x19 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x19 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x19 and x18 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and x22 and not x19 and x18 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and x22 and not x19 and x18 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x19 and x18 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x19 and not x18 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s300;

      elsif ( not x21 and not x22 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x22 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x22 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s361 =>
      if ( x22 and x19 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x22 and x19 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x22 and x19 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x22 and x19 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x22 and not x19 and x18 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x22 and not x19 and x18 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x22 and not x19 and x18 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x22 and not x19 and x18 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x22 and not x19 and not x18 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x22 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x22 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x22 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s362 =>
      if ( x22 and x19 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x22 and x19 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x22 and x19 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x22 and x19 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x22 and not x19 and x18 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( x22 and not x19 and not x18 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x22 and not x19 and not x18 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x22 and not x19 and not x18 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x22 and not x19 and not x18 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x22 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x22 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x22 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s363 =>
      if ( x65 and x67 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x67 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x65 and x67 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and x67 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x67 and x21 ) = '1' then
         y4 <= '1' ;
         y22 <= '1' ;
         y38 <= '1' ;
         current_group15m <= s95;

      elsif ( x65 and not x67 and not x21 ) = '1' then
         y35 <= '1' ;
         current_group15m <= s26;

      else
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s288;

      end if;

   when s364 =>
      if ( x19 and x18 and x14 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s338;

      elsif ( x19 and x18 and not x14 and x17 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s338;

      elsif ( x19 and x18 and not x14 and not x17 and x20 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s30;

      elsif ( x19 and x18 and not x14 and not x17 and not x20 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( x19 and not x18 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s338;

      else
         y7 <= '1' ;
         current_group15m <= s140;

      end if;

   when s365 =>
         y9 <= '1' ;
         current_group15m <= s27;

   when s366 =>
      if ( x20 and x15 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s198;

      elsif ( x20 and not x15 and x16 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s59;

      elsif ( x20 and not x15 and not x16 ) = '1' then
         y7 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s211;

      elsif ( not x20 and x21 and x17 and x15 and x8 ) = '1' then
         y8 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s254;

      elsif ( not x20 and x21 and x17 and x15 and not x8 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s198;

      elsif ( not x20 and x21 and x17 and not x15 and x16 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x20 and x21 and x17 and not x15 and not x16 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s209;

      elsif ( not x20 and x21 and not x17 ) = '1' then
         current_group15m <= s40;

      elsif ( not x20 and not x21 and x3 ) = '1' then
         current_group15m <= s40;

      elsif ( not x20 and not x21 and not x3 and x18 and x15 and x8 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( not x20 and not x21 and not x3 and x18 and x15 and not x8 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s198;

      elsif ( not x20 and not x21 and not x3 and x18 and not x15 and x16 ) = '1' then
         y10 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s47;

      elsif ( not x20 and not x21 and not x3 and x18 and not x15 and not x16 ) = '1' then
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s209;

      else
         current_group15m <= s39;

      end if;

   when s367 =>
      if ( x61 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( not x61 and x15 and x12 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s292;

      elsif ( not x61 and x15 and x12 and not x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s290;

      elsif ( not x61 and x15 and not x12 and x7 ) = '1' then
         y7 <= '1' ;
         y14 <= '1' ;
         y23 <= '1' ;
         current_group15m <= s63;

      elsif ( not x61 and x15 and not x12 and not x7 ) = '1' then
         y2 <= '1' ;
         y10 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s263;

      elsif ( not x61 and not x15 and x16 and x7 and x12 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s290;

      elsif ( not x61 and not x15 and x16 and x7 and not x12 ) = '1' then
         y5 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s262;

      elsif ( not x61 and not x15 and x16 and not x7 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s258;

      elsif ( not x61 and not x15 and not x16 and x7 ) = '1' then
         y12 <= '1' ;
         current_group15m <= s100;

      else
         y3 <= '1' ;
         current_group15m <= s89;

      end if;

   when s368 =>
      if ( x22 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s314;

      elsif ( not x22 and x19 and x15 and x8 ) = '1' then
         y11 <= '1' ;
         current_group15m <= s8;

      elsif ( not x22 and x19 and x15 and not x8 ) = '1' then
         y4 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s111;

      elsif ( not x22 and x19 and not x15 and x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s50;

      elsif ( not x22 and x19 and not x15 and not x16 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      else
         y5 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s314;

      end if;

   when s369 =>
      if ( x4 ) = '1' then
         y3 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s168;

      elsif ( not x4 and x42 and x15 and x8 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s140;

      elsif ( not x4 and x42 and x15 and not x8 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x4 and x42 and not x15 and x16 ) = '1' then
         y21 <= '1' ;
         current_group15m <= s151;

      elsif ( not x4 and x42 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s135;

      else
         y2 <= '1' ;
         y12 <= '1' ;
         y14 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s400;

      end if;

   when s370 =>
      if ( x21 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s155;

      elsif ( not x21 and x22 and x23 and x17 and x14 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x21 and x22 and x23 and x17 and not x14 and x13 ) = '1' then
         y1 <= '1' ;
         y7 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s87;

      elsif ( not x21 and x22 and x23 and x17 and not x14 and not x13 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and x23 and not x17 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x23 ) = '1' then
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s341;

      else
         y4 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s180;

      end if;

   when s371 =>
      if ( x22 ) = '1' then
         y2 <= '1' ;
         y6 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      elsif ( not x22 and x21 ) = '1' then
         y2 <= '1' ;
         y6 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      elsif ( not x22 and not x21 and x4 and x5 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x22 and not x21 and x4 and not x5 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x22 and not x21 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s372 =>
         y2 <= '1' ;
         y11 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s123;

   when s373 =>
      if ( x21 ) = '1' then
         y2 <= '1' ;
         y6 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      elsif ( not x21 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x5 and not x4 and x22 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x5 and not x4 and x22 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x5 and not x4 and not x22 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x5 and x22 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x5 and not x22 and x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and not x5 and not x22 and x4 and not x6 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s374 =>
      if ( x66 and x16 and x21 and x7 and x10 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s67;

      elsif ( x66 and x16 and x21 and x7 and not x10 ) = '1' then
         y5 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s113;

      elsif ( x66 and x16 and x21 and not x7 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s67;

      elsif ( x66 and x16 and not x21 and x7 and x10 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s75;

      elsif ( x66 and x16 and not x21 and x7 and not x10 ) = '1' then
         y4 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s395;

      elsif ( x66 and x16 and not x21 and not x7 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s75;

      elsif ( x66 and not x16 and x17 and x9 and x21 and x10 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s67;

      elsif ( x66 and not x16 and x17 and x9 and x21 and not x10 and x13 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s67;

      elsif ( x66 and not x16 and x17 and x9 and x21 and not x10 and not x13 and x19 and x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and not x16 and x17 and x9 and x21 and not x10 and not x13 and x19 and not x15 and x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and not x16 and x17 and x9 and x21 and not x10 and not x13 and x19 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and x17 and x9 and x21 and not x10 and not x13 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and x17 and x9 and not x21 and x10 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s75;

      elsif ( x66 and not x16 and x17 and x9 and not x21 and not x10 and x13 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s75;

      elsif ( x66 and not x16 and x17 and x9 and not x21 and not x10 and not x13 and x20 and x15 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x66 and not x16 and x17 and x9 and not x21 and not x10 and not x13 and x20 and not x15 and x14 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x66 and not x16 and x17 and x9 and not x21 and not x10 and not x13 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and x17 and x9 and not x21 and not x10 and not x13 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and x17 and not x9 and x21 and x10 and x11 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s67;

      elsif ( x66 and not x16 and x17 and not x9 and x21 and x10 and not x11 and x19 and x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and not x16 and x17 and not x9 and x21 and x10 and not x11 and x19 and not x15 and x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and not x16 and x17 and not x9 and x21 and x10 and not x11 and x19 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and x17 and not x9 and x21 and x10 and not x11 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and x17 and not x9 and x21 and not x10 and x12 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s67;

      elsif ( x66 and not x16 and x17 and not x9 and x21 and not x10 and not x12 and x19 and x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and not x16 and x17 and not x9 and x21 and not x10 and not x12 and x19 and not x15 and x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( x66 and not x16 and x17 and not x9 and x21 and not x10 and not x12 and x19 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and x17 and not x9 and x21 and not x10 and not x12 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and x17 and not x9 and not x21 and x10 and x11 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s75;

      elsif ( x66 and not x16 and x17 and not x9 and not x21 and x10 and not x11 and x20 and x15 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x66 and not x16 and x17 and not x9 and not x21 and x10 and not x11 and x20 and not x15 and x14 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x66 and not x16 and x17 and not x9 and not x21 and x10 and not x11 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and x17 and not x9 and not x21 and x10 and not x11 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and x17 and not x9 and not x21 and not x10 and x12 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s75;

      elsif ( x66 and not x16 and x17 and not x9 and not x21 and not x10 and not x12 and x20 and x15 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x66 and not x16 and x17 and not x9 and not x21 and not x10 and not x12 and x20 and not x15 and x14 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( x66 and not x16 and x17 and not x9 and not x21 and not x10 and not x12 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and x17 and not x9 and not x21 and not x10 and not x12 and not x20 ) = '1' then
         current_group15m <= s1;

      elsif ( x66 and not x16 and not x17 and x7 ) = '1' then
         y4 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s353;

      elsif ( x66 and not x16 and not x17 and not x7 and x21 ) = '1' then
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s67;

      elsif ( x66 and not x16 and not x17 and not x7 and not x21 ) = '1' then
         y4 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s75;

      elsif ( not x66 and x21 and x3 and x4 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( not x66 and x21 and x3 and not x4 and x5 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( not x66 and x21 and x3 and not x4 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and x21 and not x3 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x21 and x22 and x6 and x7 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x66 and not x21 and x22 and x6 and not x7 and x8 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( not x66 and not x21 and x22 and x6 and not x7 and not x8 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x21 and x22 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x66 and not x21 and not x22 and x8 and x9 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x66 and not x21 and not x22 and x8 and not x9 and x10 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s88;

      elsif ( not x66 and not x21 and not x22 and x8 and not x9 and not x10 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s375 =>
      if ( x21 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s413;

      elsif ( not x21 and not x22 and x5 ) = '1' then
         y13 <= '1' ;
         current_group15m <= s265;

      elsif ( not x21 and not x22 and not x5 and x7 and x18 and x15 ) = '1' then
         y8 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s82;

      elsif ( not x21 and not x22 and not x5 and x7 and x18 and not x15 ) = '1' then
         y2 <= '1' ;
         y4 <= '1' ;
         current_group15m <= s374;

      elsif ( not x21 and not x22 and not x5 and x7 and not x18 and x19 and x15 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s320;

      elsif ( not x21 and not x22 and not x5 and x7 and not x18 and x19 and not x15 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( not x21 and not x22 and not x5 and x7 and not x18 and not x19 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      else
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s385;

      end if;

   when s376 =>
      if ( x21 ) = '1' then
         y18 <= '1' ;
         current_group15m <= s203;

      elsif ( not x21 and x22 ) = '1' then
         y1 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s142;

      else
         y18 <= '1' ;
         current_group15m <= s114;

      end if;

   when s377 =>
      if ( x22 and x21 ) = '1' then
         y2 <= '1' ;
         y6 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      elsif ( x22 and not x21 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( x22 and not x21 and x5 and not x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( x22 and not x21 and x5 and not x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x22 and not x21 and not x5 ) = '1' then
         current_group15m <= s1;

      else
         y2 <= '1' ;
         y6 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      end if;

   when s378 =>
      if ( x21 ) = '1' then
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s126;

      elsif ( not x21 and x22 and x5 and x4 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and x5 and not x4 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and x5 and not x4 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x22 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and x19 and x15 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s103;

      elsif ( not x21 and not x22 and x19 and not x15 and x12 ) = '1' then
         y2 <= '1' ;
         y6 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s123;

      elsif ( not x21 and not x22 and x19 and not x15 and not x12 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s103;

      elsif ( not x21 and not x22 and not x19 and x20 and x14 and x15 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s103;

      elsif ( not x21 and not x22 and not x19 and x20 and x14 and not x15 and x18 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s103;

      elsif ( not x21 and not x22 and not x19 and x20 and x14 and not x15 and not x18 and x4 and x5 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and not x22 and not x19 and x20 and x14 and not x15 and not x18 and x4 and not x5 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and not x22 and not x19 and x20 and x14 and not x15 and not x18 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x19 and x20 and x14 and not x15 and not x18 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x19 and x20 and not x14 and x15 and x16 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s103;

      elsif ( not x21 and not x22 and not x19 and x20 and not x14 and x15 and not x16 and x4 and x5 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and not x22 and not x19 and x20 and not x14 and x15 and not x16 and x4 and not x5 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and not x22 and not x19 and x20 and not x14 and x15 and not x16 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x19 and x20 and not x14 and x15 and not x16 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x19 and x20 and not x14 and not x15 and x17 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s103;

      elsif ( not x21 and not x22 and not x19 and x20 and not x14 and not x15 and not x17 and x4 and x5 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and not x22 and not x19 and x20 and not x14 and not x15 and not x17 and x4 and not x5 and x6 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and not x22 and not x19 and x20 and not x14 and not x15 and not x17 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x19 and x20 and not x14 and not x15 and not x17 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x19 and not x20 and x12 ) = '1' then
         y6 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s225;

      else
         y2 <= '1' ;
         y3 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s103;

      end if;

   when s379 =>
         y8 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s106;

   when s380 =>
         y21 <= '1' ;
         current_group15m <= s7;

   when s381 =>
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

   when s382 =>
         y11 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s52;

   when s383 =>
         y4 <= '1' ;
         current_group15m <= s43;

   when s384 =>
         y18 <= '1' ;
         current_group15m <= s394;

   when s385 =>
      if ( x21 and x8 ) = '1' then
         y3 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s275;

      elsif ( x21 and not x8 and x19 and x18 and x17 and x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s272;

      elsif ( x21 and not x8 and x19 and x18 and x17 and not x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s272;

      elsif ( x21 and not x8 and x19 and x18 and not x17 and x12 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x21 and not x8 and x19 and x18 and not x17 and not x12 ) = '1' then
         y4 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s273;

      elsif ( x21 and not x8 and x19 and not x18 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s274;

      elsif ( x21 and not x8 and not x19 and x9 and x20 and x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s272;

      elsif ( x21 and not x8 and not x19 and x9 and x20 and not x12 ) = '1' then
         y2 <= '1' ;
         y9 <= '1' ;
         y10 <= '1' ;
         current_group15m <= s105;

      elsif ( x21 and not x8 and not x19 and x9 and not x20 and x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s270;

      elsif ( x21 and not x8 and not x19 and x9 and not x20 and not x12 ) = '1' then
         y16 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s109;

      elsif ( x21 and not x8 and not x19 and not x9 ) = '1' then
         y9 <= '1' ;
         y17 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s274;

      elsif ( not x21 and x22 ) = '1' then
         current_group15m <= s1;

      else
         y6 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s102;

      end if;

   when s386 =>
      if ( x6 and x7 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( x6 and not x7 and x8 ) = '1' then
         y8 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s138;

      elsif ( x6 and not x7 and not x8 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s387 =>
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s388;

   when s388 =>
         y13 <= '1' ;
         current_group15m <= s265;

   when s389 =>
         y3 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s255;

   when s390 =>
      if ( x21 and x20 ) = '1' then
         y5 <= '1' ;
         y6 <= '1' ;
         current_group15m <= s133;

      elsif ( x21 and not x20 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      else
         y10 <= '1' ;
         current_group15m <= s12;

      end if;

   when s391 =>
      if ( x3 ) = '1' then
         y3 <= '1' ;
         y7 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s420;

      elsif ( not x3 and x8 and x21 and x16 and x13 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( not x3 and x8 and x21 and x16 and not x13 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s360;

      elsif ( not x3 and x8 and x21 and not x16 and x17 and x18 and x13 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s249;

      elsif ( not x3 and x8 and x21 and not x16 and x17 and x18 and not x13 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( not x3 and x8 and x21 and not x16 and x17 and not x18 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( not x3 and x8 and x21 and not x16 and not x17 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s146;

      elsif ( not x3 and x8 and not x21 and x22 and x16 and x19 and x18 and x10 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x3 and x8 and not x21 and x22 and x16 and x19 and x18 and not x10 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s362;

      elsif ( not x3 and x8 and not x21 and x22 and x16 and x19 and not x18 and x13 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x3 and x8 and not x21 and x22 and x16 and x19 and not x18 and not x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x3 and x8 and not x21 and x22 and x16 and not x19 and x13 ) = '1' then
         y3 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s146;

      elsif ( not x3 and x8 and not x21 and x22 and x16 and not x19 and not x13 and x18 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( not x3 and x8 and not x21 and x22 and x16 and not x19 and not x13 and not x18 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x3 and x8 and not x21 and x22 and not x16 and x17 and x19 and x18 and x10 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

      elsif ( not x3 and x8 and not x21 and x22 and not x16 and x17 and x19 and x18 and not x10 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s146;

      elsif ( not x3 and x8 and not x21 and x22 and not x16 and x17 and x19 and not x18 and x13 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

      elsif ( not x3 and x8 and not x21 and x22 and not x16 and x17 and x19 and not x18 and not x13 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( not x3 and x8 and not x21 and x22 and not x16 and x17 and not x19 and x13 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

      elsif ( not x3 and x8 and not x21 and x22 and not x16 and x17 and not x19 and not x13 and x18 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x3 and x8 and not x21 and x22 and not x16 and x17 and not x19 and not x13 and not x18 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( not x3 and x8 and not x21 and x22 and not x16 and not x17 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s146;

      elsif ( not x3 and x8 and not x21 and not x22 and x19 and x17 and x13 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x3 and x8 and not x21 and not x22 and x19 and x17 and not x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x3 and x8 and not x21 and not x22 and x19 and not x17 and x18 and x13 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

      elsif ( not x3 and x8 and not x21 and not x22 and x19 and not x17 and x18 and not x13 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( not x3 and x8 and not x21 and not x22 and x19 and not x17 and not x18 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s146;

      elsif ( not x3 and x8 and not x21 and not x22 and not x19 and x16 and x13 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( not x3 and x8 and not x21 and not x22 and not x19 and x16 and not x13 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s360;

      elsif ( not x3 and x8 and not x21 and not x22 and not x19 and not x16 and x17 and x20 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( not x3 and x8 and not x21 and not x22 and not x19 and not x16 and x17 and not x20 and x13 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s249;

      elsif ( not x3 and x8 and not x21 and not x22 and not x19 and not x16 and x17 and not x20 and not x13 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( not x3 and x8 and not x21 and not x22 and not x19 and not x16 and not x17 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s146;

      else
         y3 <= '1' ;
         y8 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s421;

      end if;

   when s392 =>
      if ( x68 ) = '1' then
         y6 <= '1' ;
         y7 <= '1' ;
         current_group15m <= s76;

      else
         y5 <= '1' ;
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s282;

      end if;

   when s393 =>
      if ( x20 and x18 and x13 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x20 and x18 and not x13 and x12 ) = '1' then
         y9 <= '1' ;
         current_group15m <= s27;

      elsif ( x20 and x18 and not x13 and not x12 ) = '1' then
         current_group15m <= s1;

      elsif ( x20 and not x18 ) = '1' then
         current_group15m <= s1;

      else
         y2 <= '1' ;
         current_group15m <= s56;

      end if;

   when s394 =>
         y4 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s273;

   when s395 =>
      if ( x65 and x5 and x6 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x5 and not x6 and x7 ) = '1' then
         y5 <= '1' ;
         current_group15m <= s101;

      elsif ( x65 and x5 and not x6 and not x7 ) = '1' then
         current_group15m <= s1;

      elsif ( x65 and not x5 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and x19 and x15 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and x21 and x19 and not x15 and x14 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s92;

      elsif ( not x65 and x21 and x19 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and x21 and not x19 ) = '1' then
         current_group15m <= s1;

      elsif ( not x65 and not x21 and x20 and x15 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( not x65 and not x21 and x20 and not x15 and x14 ) = '1' then
         y27 <= '1' ;
         current_group15m <= s3;

      elsif ( not x65 and not x21 and x20 and not x15 and not x14 ) = '1' then
         current_group15m <= s1;

      else
         current_group15m <= s1;

      end if;

   when s396 =>
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s375;

   when s397 =>
      if ( x63 and x15 and x8 ) = '1' then
         y2 <= '1' ;
         y3 <= '1' ;
         current_group15m <= s23;

      elsif ( x63 and x15 and not x8 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x63 and not x15 and x16 ) = '1' then
         y19 <= '1' ;
         current_group15m <= s11;

      elsif ( x63 and not x15 and not x16 ) = '1' then
         y13 <= '1' ;
         y14 <= '1' ;
         y29 <= '1' ;
         current_group15m <= s135;

      else
         current_group15m <= s1;

      end if;

   when s398 =>
      if ( x19 and x14 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( x19 and not x14 and x13 ) = '1' then
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s175;

      elsif ( x19 and not x14 and not x13 ) = '1' then
         current_group15m <= s398;

      else
         current_group15m <= s1;

      end if;

   when s399 =>
      if ( x66 ) = '1' then
         y15 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s137;

      else
         y11 <= '1' ;
         current_group15m <= s53;

      end if;

   when s400 =>
         y3 <= '1' ;
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s130;

   when s401 =>
      if ( x20 ) = '1' then
         y2 <= '1' ;
         y7 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s366;

      else
         current_group15m <= s1;

      end if;

   when s402 =>
      if ( x25 and x24 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( x25 and not x24 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      else
         y24 <= '1' ;
         current_group15m <= s278;

      end if;

   when s403 =>
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s59;

   when s404 =>
      if ( x3 ) = '1' then
         y4 <= '1' ;
         y5 <= '1' ;
         current_group15m <= s250;

      elsif ( not x3 and x19 ) = '1' then
         y14 <= '1' ;
         current_group15m <= s285;

      else
         y14 <= '1' ;
         y21 <= '1' ;
         y22 <= '1' ;
         current_group15m <= s84;

      end if;

   when s405 =>
      if ( x21 and x20 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( x21 and not x20 ) = '1' then
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s302;

      else
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s302;

      end if;

   when s406 =>
         y8 <= '1' ;
         current_group15m <= s246;

   when s407 =>
         y20 <= '1' ;
         current_group15m <= s13;

   when s408 =>
      if ( x21 and x18 and x16 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s1;

      elsif ( x21 and x18 and not x16 and x17 and x13 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s1;

      elsif ( x21 and x18 and not x16 and x17 and not x13 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x21 and x18 and not x16 and x17 and not x13 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x21 and x18 and not x16 and x17 and not x13 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x18 and not x16 and x17 and not x13 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and x18 and not x16 and not x17 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s1;

      elsif ( x21 and not x18 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x21 and not x18 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( x21 and not x18 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( x21 and not x18 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and x19 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s1;

      elsif ( not x21 and not x19 and x22 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s1;

      elsif ( not x21 and not x19 and not x22 and x20 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x19 and not x22 and x20 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x19 and not x22 and x20 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x19 and not x22 and x20 and not x4 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x19 and not x22 and not x20 and x16 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s1;

      elsif ( not x21 and not x19 and not x22 and not x20 and not x16 and x13 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s1;

      elsif ( not x21 and not x19 and not x22 and not x20 and not x16 and not x13 and x17 and x4 and x5 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x19 and not x22 and not x20 and not x16 and not x13 and x17 and x4 and not x5 and x6 ) = '1' then
         y10 <= '1' ;
         current_group15m <= s12;

      elsif ( not x21 and not x19 and not x22 and not x20 and not x16 and not x13 and x17 and x4 and not x5 and not x6 ) = '1' then
         current_group15m <= s1;

      elsif ( not x21 and not x19 and not x22 and not x20 and not x16 and not x13 and x17 and not x4 ) = '1' then
         current_group15m <= s1;

      else
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s1;

      end if;

   when s409 =>
      if ( x21 and x18 and x13 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x21 and x18 and not x13 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s1;

      elsif ( x21 and not x18 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s1;

      elsif ( not x21 and x22 and x18 and x19 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x21 and x22 and x18 and not x19 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( not x21 and x22 and not x18 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s146;

      elsif ( not x21 and not x22 and x19 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s146;

      elsif ( not x21 and not x22 and not x19 and x13 and x20 ) = '1' then
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s1;

      elsif ( not x21 and not x22 and not x19 and x13 and not x20 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      else
         y5 <= '1' ;
         y16 <= '1' ;
         y17 <= '1' ;
         current_group15m <= s1;

      end if;

   when s410 =>
         y9 <= '1' ;
         y14 <= '1' ;
         current_group15m <= s336;

   when s411 =>
      if ( x61 ) = '1' then
         current_group15m <= s1;

      else
         y2 <= '1' ;
         y8 <= '1' ;
         current_group15m <= s367;

      end if;

   when s412 =>
      if ( x4 and x19 and x20 and x14 ) = '1' then
         y16 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s422;

      elsif ( x4 and x19 and x20 and not x14 and x16 ) = '1' then
         y16 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s422;

      elsif ( x4 and x19 and x20 and not x14 and not x16 and x17 ) = '1' then
         y16 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s352;

      elsif ( x4 and x19 and x20 and not x14 and not x16 and not x17 ) = '1' then
         y16 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s422;

      elsif ( x4 and x19 and not x20 ) = '1' then
         y16 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s422;

      elsif ( x4 and not x19 ) = '1' then
         y16 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s422;

      elsif ( not x4 and x9 and x17 and x19 and x20 and x14 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( not x4 and x9 and x17 and x19 and x20 and not x14 and x16 ) = '1' then
         y4 <= '1' ;
         y29 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s351;

      elsif ( not x4 and x9 and x17 and x19 and x20 and not x14 and not x16 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s415;

      elsif ( not x4 and x9 and x17 and x19 and not x20 and x14 ) = '1' then
         y4 <= '1' ;
         y18 <= '1' ;
         y29 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s351;

      elsif ( not x4 and x9 and x17 and x19 and not x20 and not x14 and x16 ) = '1' then
         y29 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s351;

      elsif ( not x4 and x9 and x17 and x19 and not x20 and not x14 and not x16 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s351;

      elsif ( not x4 and x9 and x17 and not x19 and x16 ) = '1' then
         y29 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s351;

      elsif ( not x4 and x9 and x17 and not x19 and not x16 and x20 ) = '1' then
         y9 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s351;

      elsif ( not x4 and x9 and x17 and not x19 and not x16 and not x20 and x15 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x4 and x9 and x17 and not x19 and not x16 and not x20 and not x15 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( not x4 and x9 and not x17 and x18 and x19 and x14 and x16 ) = '1' then
         y2 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s349;

      elsif ( not x4 and x9 and not x17 and x18 and x19 and x14 and not x16 ) = '1' then
         y2 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s416;

      elsif ( not x4 and x9 and not x17 and x18 and x19 and not x14 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s338;

      elsif ( not x4 and x9 and not x17 and x18 and not x19 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s338;

      elsif ( not x4 and x9 and not x17 and not x18 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( not x4 and not x9 and x19 and x20 and x17 and x16 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s415;

      elsif ( not x4 and not x9 and x19 and x20 and x17 and not x16 and x14 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s415;

      elsif ( not x4 and not x9 and x19 and x20 and x17 and not x16 and not x14 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( not x4 and not x9 and x19 and x20 and not x17 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s415;

      elsif ( not x4 and not x9 and x19 and not x20 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s415;

      elsif ( not x4 and not x9 and not x19 and x20 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s415;

      elsif ( not x4 and not x9 and not x19 and not x20 and x17 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s415;

      elsif ( not x4 and not x9 and not x19 and not x20 and not x17 and x18 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s241;

      else
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s415;

      end if;

   when s413 =>
      if ( x22 ) = '1' then
         y3 <= '1' ;
         y14 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s385;

      else
         y3 <= '1' ;
         current_group15m <= s320;

      end if;

   when s414 =>
         y7 <= '1' ;
         current_group15m <= s140;

   when s415 =>
      if ( x17 and x19 and x20 and x14 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( x17 and x19 and x20 and not x14 and x16 ) = '1' then
         y4 <= '1' ;
         y29 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s351;

      elsif ( x17 and x19 and x20 and not x14 and not x16 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( x17 and x19 and not x20 and x14 ) = '1' then
         y4 <= '1' ;
         y18 <= '1' ;
         y29 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s351;

      elsif ( x17 and x19 and not x20 and not x14 and x16 ) = '1' then
         y29 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s351;

      elsif ( x17 and x19 and not x20 and not x14 and not x16 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s351;

      elsif ( x17 and not x19 and x16 ) = '1' then
         y29 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s351;

      elsif ( x17 and not x19 and not x16 and x20 ) = '1' then
         y9 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s351;

      elsif ( x17 and not x19 and not x16 and not x20 and x15 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( x17 and not x19 and not x16 and not x20 and not x15 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( not x17 and x18 and x19 and x14 and x16 ) = '1' then
         y2 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s349;

      elsif ( not x17 and x18 and x19 and x14 and not x16 ) = '1' then
         y2 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s416;

      elsif ( not x17 and x18 and x19 and not x14 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s338;

      elsif ( not x17 and x18 and not x19 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s338;

      else
         y4 <= '1' ;
         current_group15m <= s43;

      end if;

   when s416 =>
      if ( x20 ) = '1' then
         y8 <= '1' ;
         current_group15m <= s246;

      else
         y6 <= '1' ;
         y20 <= '1' ;
         current_group15m <= s102;

      end if;

   when s417 =>
         y4 <= '1' ;
         y5 <= '1' ;
         y9 <= '1' ;
         current_group15m <= s80;

   when s418 =>
      if ( x21 and x13 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s249;

      elsif ( x21 and not x13 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( not x21 and x19 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

      elsif ( not x21 and not x19 and x22 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

      elsif ( not x21 and not x19 and not x22 and x13 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s249;

      else
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      end if;

   when s419 =>
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

   when s420 =>
      if ( x8 and x21 and x16 and x13 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x8 and x21 and x16 and not x13 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s360;

      elsif ( x8 and x21 and not x16 and x17 and x18 and x13 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s249;

      elsif ( x8 and x21 and not x16 and x17 and x18 and not x13 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( x8 and x21 and not x16 and x17 and not x18 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( x8 and x21 and not x16 and not x17 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s146;

      elsif ( x8 and not x21 and x22 and x16 and x19 and x18 and x10 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( x8 and not x21 and x22 and x16 and x19 and x18 and not x10 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s362;

      elsif ( x8 and not x21 and x22 and x16 and x19 and not x18 and x13 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( x8 and not x21 and x22 and x16 and x19 and not x18 and not x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x8 and not x21 and x22 and x16 and not x19 and x13 ) = '1' then
         y3 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s146;

      elsif ( x8 and not x21 and x22 and x16 and not x19 and not x13 and x18 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( x8 and not x21 and x22 and x16 and not x19 and not x13 and not x18 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( x8 and not x21 and x22 and not x16 and x17 and x19 and x18 and x10 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

      elsif ( x8 and not x21 and x22 and not x16 and x17 and x19 and x18 and not x10 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s146;

      elsif ( x8 and not x21 and x22 and not x16 and x17 and x19 and not x18 and x13 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

      elsif ( x8 and not x21 and x22 and not x16 and x17 and x19 and not x18 and not x13 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( x8 and not x21 and x22 and not x16 and x17 and not x19 and x13 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

      elsif ( x8 and not x21 and x22 and not x16 and x17 and not x19 and not x13 and x18 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( x8 and not x21 and x22 and not x16 and x17 and not x19 and not x13 and not x18 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( x8 and not x21 and x22 and not x16 and not x17 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s146;

      elsif ( x8 and not x21 and not x22 and x19 and x17 and x13 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( x8 and not x21 and not x22 and x19 and x17 and not x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( x8 and not x21 and not x22 and x19 and not x17 and x18 and x13 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

      elsif ( x8 and not x21 and not x22 and x19 and not x17 and x18 and not x13 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( x8 and not x21 and not x22 and x19 and not x17 and not x18 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s146;

      elsif ( x8 and not x21 and not x22 and not x19 and x16 and x13 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x8 and not x21 and not x22 and not x19 and x16 and not x13 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s360;

      elsif ( x8 and not x21 and not x22 and not x19 and not x16 and x17 and x20 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( x8 and not x21 and not x22 and not x19 and not x16 and x17 and not x20 and x13 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s249;

      elsif ( x8 and not x21 and not x22 and not x19 and not x16 and x17 and not x20 and not x13 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( x8 and not x21 and not x22 and not x19 and not x16 and not x17 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s146;

      else
         y3 <= '1' ;
         y8 <= '1' ;
         y12 <= '1' ;
         y13 <= '1' ;
         current_group15m <= s421;

      end if;

   when s421 =>
      if ( x21 and x16 and x13 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x21 and x16 and not x13 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s360;

      elsif ( x21 and not x16 and x17 and x18 and x13 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s249;

      elsif ( x21 and not x16 and x17 and x18 and not x13 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( x21 and not x16 and x17 and not x18 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( x21 and not x16 and not x17 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s146;

      elsif ( not x21 and x22 and x16 and x19 and x18 and x10 ) = '1' then
         y3 <= '1' ;
         current_group15m <= s89;

      elsif ( not x21 and x22 and x16 and x19 and x18 and not x10 ) = '1' then
         y5 <= '1' ;
         y8 <= '1' ;
         y11 <= '1' ;
         y12 <= '1' ;
         current_group15m <= s362;

      elsif ( not x21 and x22 and x16 and x19 and not x18 and x13 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and x22 and x16 and x19 and not x18 and not x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x21 and x22 and x16 and not x19 and x13 ) = '1' then
         y3 <= '1' ;
         y16 <= '1' ;
         current_group15m <= s146;

      elsif ( not x21 and x22 and x16 and not x19 and not x13 and x18 ) = '1' then
         y5 <= '1' ;
         y12 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s146;

      elsif ( not x21 and x22 and x16 and not x19 and not x13 and not x18 ) = '1' then
         y24 <= '1' ;
         current_group15m <= s278;

      elsif ( not x21 and x22 and not x16 and x17 and x18 and x19 and x10 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

      elsif ( not x21 and x22 and not x16 and x17 and x18 and x19 and not x10 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y18 <= '1' ;
         y19 <= '1' ;
         current_group15m <= s146;

      elsif ( not x21 and x22 and not x16 and x17 and x18 and not x19 and x13 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

      elsif ( not x21 and x22 and not x16 and x17 and x18 and not x19 and not x13 ) = '1' then
         y16 <= '1' ;
         current_group15m <= s16;

      elsif ( not x21 and x22 and not x16 and x17 and not x18 and x13 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

      elsif ( not x21 and x22 and not x16 and x17 and not x18 and not x13 and x19 ) = '1' then
         y7 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s146;

      elsif ( not x21 and x22 and not x16 and x17 and not x18 and not x13 and not x19 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( not x21 and x22 and not x16 and not x17 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s146;

      elsif ( not x21 and not x22 and x19 and x17 and x13 ) = '1' then
         y15 <= '1' ;
         current_group15m <= s149;

      elsif ( not x21 and not x22 and x19 and x17 and not x13 ) = '1' then
         y23 <= '1' ;
         current_group15m <= s83;

      elsif ( not x21 and not x22 and x19 and not x17 and x18 and x13 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s248;

      elsif ( not x21 and not x22 and x19 and not x17 and x18 and not x13 ) = '1' then
         y7 <= '1' ;
         y11 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s358;

      elsif ( not x21 and not x22 and x19 and not x17 and not x18 ) = '1' then
         y8 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s146;

      elsif ( not x21 and not x22 and not x19 and x16 and x13 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( not x21 and not x22 and not x19 and x16 and not x13 ) = '1' then
         y7 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s360;

      elsif ( not x21 and not x22 and not x19 and not x16 and x17 and x20 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      elsif ( not x21 and not x22 and not x19 and not x16 and x17 and not x20 and x13 ) = '1' then
         y1 <= '1' ;
         y25 <= '1' ;
         current_group15m <= s249;

      elsif ( not x21 and not x22 and not x19 and not x16 and x17 and not x20 and not x13 ) = '1' then
         y2 <= '1' ;
         y12 <= '1' ;
         y15 <= '1' ;
         current_group15m <= s408;

      else
         y8 <= '1' ;
         y9 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s146;

      end if;

   when s422 =>
      if ( x9 and x17 and x19 and x20 and x14 ) = '1' then
         y2 <= '1' ;
         current_group15m <= s56;

      elsif ( x9 and x17 and x19 and x20 and not x14 ) = '1' then
         y4 <= '1' ;
         y29 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s351;

      elsif ( x9 and x17 and x19 and not x20 and x14 ) = '1' then
         y4 <= '1' ;
         y18 <= '1' ;
         y29 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s351;

      elsif ( x9 and x17 and x19 and not x20 and not x14 and x16 ) = '1' then
         y29 <= '1' ;
         y31 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s351;

      elsif ( x9 and x17 and x19 and not x20 and not x14 and not x16 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         y18 <= '1' ;
         current_group15m <= s351;

      elsif ( x9 and x17 and not x19 and x16 ) = '1' then
         y29 <= '1' ;
         y30 <= '1' ;
         current_group15m <= s351;

      elsif ( x9 and x17 and not x19 and not x16 and x20 ) = '1' then
         y9 <= '1' ;
         y26 <= '1' ;
         current_group15m <= s351;

      elsif ( x9 and x17 and not x19 and not x16 and not x20 and x15 ) = '1' then
         y4 <= '1' ;
         y11 <= '1' ;
         current_group15m <= s112;

      elsif ( x9 and x17 and not x19 and not x16 and not x20 and not x15 ) = '1' then
         y25 <= '1' ;
         current_group15m <= s78;

      elsif ( x9 and not x17 and x18 and x19 and x14 and x16 ) = '1' then
         y2 <= '1' ;
         y14 <= '1' ;
         y19 <= '1' ;
         y29 <= '1' ;
         y30 <= '1' ;
         y32 <= '1' ;
         current_group15m <= s349;

      elsif ( x9 and not x17 and x18 and x19 and x14 and not x16 ) = '1' then
         y2 <= '1' ;
         y21 <= '1' ;
         current_group15m <= s416;

      elsif ( x9 and not x17 and x18 and x19 and not x14 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s338;

      elsif ( x9 and not x17 and x18 and not x19 ) = '1' then
         y7 <= '1' ;
         current_group15m <= s338;

      elsif ( x9 and not x17 and not x18 ) = '1' then
         y4 <= '1' ;
         current_group15m <= s43;

      elsif ( not x9 and x19 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s415;

      elsif ( not x9 and not x19 and x20 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s415;

      elsif ( not x9 and not x19 and not x20 and x17 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s415;

      elsif ( not x9 and not x19 and not x20 and not x17 and x18 ) = '1' then
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s241;

      else
         y17 <= '1' ;
         y20 <= '1' ;
         y28 <= '1' ;
         current_group15m <= s415;

      end if;

   end case;
   end proc_group15m;

   begin
      if ( rst = '1' ) then
	y1   <= '0' ;	y2   <= '0' ;	y3   <= '0' ;	y4   <= '0' ;
	y5   <= '0' ;	y6   <= '0' ;	y7   <= '0' ;	y8   <= '0' ;
	y9   <= '0' ;	y10  <= '0' ;	y11  <= '0' ;	y12  <= '0' ;
	y13  <= '0' ;	y14  <= '0' ;	y15  <= '0' ;	y16  <= '0' ;
	y17  <= '0' ;	y18  <= '0' ;	y19  <= '0' ;	y20  <= '0' ;
	y21  <= '0' ;	y22  <= '0' ;	y23  <= '0' ;	y24  <= '0' ;
	y25  <= '0' ;	y26  <= '0' ;	y27  <= '0' ;	y28  <= '0' ;
	y29  <= '0' ;	y30  <= '0' ;	y31  <= '0' ;	y32  <= '0' ;
	y33  <= '0' ;	y34  <= '0' ;	y35  <= '0' ;	y36  <= '0' ;
	y37  <= '0' ;	y38  <= '0' ;	y112 <= '0' ;
	current_group15m <= s1;
      elsif (clk'event and clk ='1') then
        proc_group15m;
      end if;
   end process;
end ARC;
