module group15m ( clk,rst,
	x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15,
	x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x42, x45, x51, x59, x60,
	x61, x62, x63, x64, x65, x66, x67, x68, 
	y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15,
	y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30,
	y31, y32, y33, y34, y35, y36, y37, y38, y112);

input clk, rst, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15,
	x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x42, x45, x51, x59, x60,
	x61, x62, x63, x64, x65, x66, x67, x68;
output y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15,
	y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30,
	y31, y32, y33, y34, y35, y36, y37, y38, y112;
reg y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15,
	y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30,
	y31, y32, y33, y34, y35, y36, y37, y38, y112;

parameter s1=1, s2=2, s3=3, s4=4, s5=5, s6=6, s7=7, s8=8, s9=9, s10=10,
	s11=11, s12=12, s13=13, s14=14, s15=15, s16=16, s17=17, s18=18, s19=19, s20=20,
	s21=21, s22=22, s23=23, s24=24, s25=25, s26=26, s27=27, s28=28, s29=29, s30=30,
	s31=31, s32=32, s33=33, s34=34, s35=35, s36=36, s37=37, s38=38, s39=39, s40=40,
	s41=41, s42=42, s43=43, s44=44, s45=45, s46=46, s47=47, s48=48, s49=49, s50=50,
	s51=51, s52=52, s53=53, s54=54, s55=55, s56=56, s57=57, s58=58, s59=59, s60=60,
	s61=61, s62=62, s63=63, s64=64, s65=65, s66=66, s67=67, s68=68, s69=69, s70=70,
	s71=71, s72=72, s73=73, s74=74, s75=75, s76=76, s77=77, s78=78, s79=79, s80=80,
	s81=81, s82=82, s83=83, s84=84, s85=85, s86=86, s87=87, s88=88, s89=89, s90=90,
	s91=91, s92=92, s93=93, s94=94, s95=95, s96=96, s97=97, s98=98, s99=99, s100=100,
	s101=101, s102=102, s103=103, s104=104, s105=105, s106=106, s107=107, s108=108, s109=109, s110=110,
	s111=111, s112=112, s113=113, s114=114, s115=115, s116=116, s117=117, s118=118, s119=119, s120=120,
	s121=121, s122=122, s123=123, s124=124, s125=125, s126=126, s127=127, s128=128, s129=129, s130=130,
	s131=131, s132=132, s133=133, s134=134, s135=135, s136=136, s137=137, s138=138, s139=139, s140=140,
	s141=141, s142=142, s143=143, s144=144, s145=145, s146=146, s147=147, s148=148, s149=149, s150=150,
	s151=151, s152=152, s153=153, s154=154, s155=155, s156=156, s157=157, s158=158, s159=159, s160=160,
	s161=161, s162=162, s163=163, s164=164, s165=165, s166=166, s167=167, s168=168, s169=169, s170=170,
	s171=171, s172=172, s173=173, s174=174, s175=175, s176=176, s177=177, s178=178, s179=179, s180=180,
	s181=181, s182=182, s183=183, s184=184, s185=185, s186=186, s187=187, s188=188, s189=189, s190=190,
	s191=191, s192=192, s193=193, s194=194, s195=195, s196=196, s197=197, s198=198, s199=199, s200=200,
	s201=201, s202=202, s203=203, s204=204, s205=205, s206=206, s207=207, s208=208, s209=209, s210=210,
	s211=211, s212=212, s213=213, s214=214, s215=215, s216=216, s217=217, s218=218, s219=219, s220=220,
	s221=221, s222=222, s223=223, s224=224, s225=225, s226=226, s227=227, s228=228, s229=229, s230=230,
	s231=231, s232=232, s233=233, s234=234, s235=235, s236=236, s237=237, s238=238, s239=239, s240=240,
	s241=241, s242=242, s243=243, s244=244, s245=245, s246=246, s247=247, s248=248, s249=249, s250=250,
	s251=251, s252=252, s253=253, s254=254, s255=255, s256=256, s257=257, s258=258, s259=259, s260=260,
	s261=261, s262=262, s263=263, s264=264, s265=265, s266=266, s267=267, s268=268, s269=269, s270=270,
	s271=271, s272=272, s273=273, s274=274, s275=275, s276=276, s277=277, s278=278, s279=279, s280=280,
	s281=281, s282=282, s283=283, s284=284, s285=285, s286=286, s287=287, s288=288, s289=289, s290=290,
	s291=291, s292=292, s293=293, s294=294, s295=295, s296=296, s297=297, s298=298, s299=299, s300=300,
	s301=301, s302=302, s303=303, s304=304, s305=305, s306=306, s307=307, s308=308, s309=309, s310=310,
	s311=311, s312=312, s313=313, s314=314, s315=315, s316=316, s317=317, s318=318, s319=319, s320=320,
	s321=321, s322=322, s323=323, s324=324, s325=325, s326=326, s327=327, s328=328, s329=329, s330=330,
	s331=331, s332=332, s333=333, s334=334, s335=335, s336=336, s337=337, s338=338, s339=339, s340=340,
	s341=341, s342=342, s343=343, s344=344, s345=345, s346=346, s347=347, s348=348, s349=349, s350=350,
	s351=351, s352=352, s353=353, s354=354, s355=355, s356=356, s357=357, s358=358, s359=359, s360=360,
	s361=361, s362=362, s363=363, s364=364, s365=365, s366=366, s367=367, s368=368, s369=369, s370=370,
	s371=371, s372=372, s373=373, s374=374, s375=375, s376=376, s377=377, s378=378, s379=379, s380=380,
	s381=381, s382=382, s383=383, s384=384, s385=385, s386=386, s387=387, s388=388, s389=389, s390=390,
	s391=391, s392=392, s393=393, s394=394, s395=395, s396=396, s397=397, s398=398, s399=399, s400=400,
	s401=401, s402=402, s403=403, s404=404, s405=405, s406=406, s407=407, s408=408, s409=409, s410=410,
	s411=411, s412=412, s413=413, s414=414, s415=415, s416=416, s417=417, s418=418, s419=419, s420=420,
	s421=421, s422=422;
integer pr_state;
integer nx_state;

always@ ( posedge rst or negedge clk )
begin
	if ( rst == 1'b1 )
		pr_state = s1;
	else
		pr_state = nx_state;
end

always@ ( pr_state or x1 or x2 or x3 or x4 or x5 or x6 or x7 or x8 or x9 or x10 or x11 or x12 or x13 or x14 or x15 or 
	x16 or x17 or x18 or x19 or x20 or x21 or x22 or x23 or x24 or x25 or x26 or x42 or x45 or x51 or x59 or x60 or 
	x61 or x62 or x63 or x64 or x65 or x66 or x67 or x68)
	begin
			y1 = 1'b0;	y2 = 1'b0;	y3 = 1'b0;	y4 = 1'b0;	
			y5 = 1'b0;	y6 = 1'b0;	y7 = 1'b0;	y8 = 1'b0;	
			y9 = 1'b0;	y10 = 1'b0;	y11 = 1'b0;	y12 = 1'b0;	
			y13 = 1'b0;	y14 = 1'b0;	y15 = 1'b0;	y16 = 1'b0;	
			y17 = 1'b0;	y18 = 1'b0;	y19 = 1'b0;	y20 = 1'b0;	
			y21 = 1'b0;	y22 = 1'b0;	y23 = 1'b0;	y24 = 1'b0;	
			y25 = 1'b0;	y26 = 1'b0;	y27 = 1'b0;	y28 = 1'b0;	
			y29 = 1'b0;	y30 = 1'b0;	y31 = 1'b0;	y32 = 1'b0;	
			y33 = 1'b0;	y34 = 1'b0;	y35 = 1'b0;	y36 = 1'b0;	
			y37 = 1'b0;	y38 = 1'b0;	y112 = 1'b0;	
		case ( pr_state )
				s1 : if( x67 && x66 && x65 && x22 && x5 && x21 && x1 )
						begin
							y10 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s2;
						end
					else if( x67 && x66 && x65 && x22 && x5 && x21 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && x65 && x22 && x5 && ~x21 && x1 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x67 && x66 && x65 && x22 && x5 && ~x21 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && x65 && x22 && ~x5 && x6 && x1 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x67 && x66 && x65 && x22 && ~x5 && x6 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && x65 && x22 && ~x5 && ~x6 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s5;
						end
					else if( x67 && x66 && x65 && x22 && ~x5 && ~x6 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && x65 && ~x22 && x4 && x17 && x23 && x1 )
						begin
							y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s1;
						end
					else if( x67 && x66 && x65 && ~x22 && x4 && x17 && x23 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && x65 && ~x22 && x4 && x17 && ~x23 && x1 )
						begin
							y3 = 1'b1;	y11 = 1'b1;	
							nx_state = s6;
						end
					else if( x67 && x66 && x65 && ~x22 && x4 && x17 && ~x23 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && x65 && ~x22 && x4 && ~x17 && x23 && x1 )
						begin
							y3 = 1'b1;	y11 = 1'b1;	
							nx_state = s6;
						end
					else if( x67 && x66 && x65 && ~x22 && x4 && ~x17 && x23 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && x65 && ~x22 && x4 && ~x17 && ~x23 && x1 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x67 && x66 && x65 && ~x22 && x4 && ~x17 && ~x23 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && x65 && ~x22 && ~x4 && x5 && x23 && x1 )
						begin
							y11 = 1'b1;	
							nx_state = s8;
						end
					else if( x67 && x66 && x65 && ~x22 && ~x4 && x5 && x23 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && x65 && ~x22 && ~x4 && x5 && ~x23 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y10 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s9;
						end
					else if( x67 && x66 && x65 && ~x22 && ~x4 && x5 && ~x23 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && x65 && ~x22 && ~x4 && ~x5 && x23 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x67 && x66 && x65 && ~x22 && ~x4 && ~x5 && x23 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && x65 && ~x22 && ~x4 && ~x5 && ~x23 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s5;
						end
					else if( x67 && x66 && x65 && ~x22 && ~x4 && ~x5 && ~x23 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && ~x65 && x68 && x1 && x21 && x6 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( x67 && x66 && ~x65 && x68 && x1 && x21 && ~x6 && x5 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x67 && x66 && ~x65 && x68 && x1 && x21 && ~x6 && x5 && ~x18 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x67 && x66 && ~x65 && x68 && x1 && x21 && ~x6 && ~x5 && x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s14;
						end
					else if( x67 && x66 && ~x65 && x68 && x1 && x21 && ~x6 && ~x5 && ~x4 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s15;
						end
					else if( x67 && x66 && ~x65 && x68 && x1 && ~x21 && x4 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( x67 && x66 && ~x65 && x68 && x1 && ~x21 && ~x4 && x5 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x67 && x66 && ~x65 && x68 && x1 && ~x21 && ~x4 && x5 && ~x18 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x67 && x66 && ~x65 && x68 && x1 && ~x21 && ~x4 && ~x5 && x6 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x67 && x66 && ~x65 && x68 && x1 && ~x21 && ~x4 && ~x5 && ~x6 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s15;
						end
					else if( x67 && x66 && ~x65 && x68 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && ~x65 && ~x68 && x62 && x5 && x51 && x1 )
						begin
							y17 = 1'b1;	
							nx_state = s17;
						end
					else if( x67 && x66 && ~x65 && ~x68 && x62 && x5 && x51 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && ~x65 && ~x68 && x62 && x5 && ~x51 && x1 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	
							nx_state = s1;
						end
					else if( x67 && x66 && ~x65 && ~x68 && x62 && x5 && ~x51 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && ~x65 && ~x68 && x62 && ~x5 && x2 && x1 )
						begin
							y14 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s18;
						end
					else if( x67 && x66 && ~x65 && ~x68 && x62 && ~x5 && x2 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && ~x65 && ~x68 && x62 && ~x5 && ~x2 && x1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s19;
						end
					else if( x67 && x66 && ~x65 && ~x68 && x62 && ~x5 && ~x2 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && x64 && x4 && x5 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s20;
						end
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && x64 && x4 && ~x5 )
						nx_state = s1;
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && x64 && ~x4 && x5 && x3 )
						begin
							y34 = 1'b1;	
							nx_state = s21;
						end
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && x64 && ~x4 && x5 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s22;
						end
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && x64 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && ~x64 && x2 && x1 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && ~x64 && x2 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && ~x64 && ~x2 && x4 && x1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && ~x64 && ~x2 && x4 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && ~x64 && ~x2 && ~x4 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s22;
						end
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && x63 && ~x64 && ~x2 && ~x4 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && x64 && x5 && x17 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s22;
						end
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && x64 && x5 && x17 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && x64 && x5 && ~x17 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && x64 && x5 && ~x17 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && x64 && ~x5 && x2 && x1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && x64 && ~x5 && x2 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && x64 && ~x5 && ~x2 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && x64 && ~x5 && ~x2 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && ~x64 && x5 && x18 && x1 )
						begin
							y35 = 1'b1;	
							nx_state = s26;
						end
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && ~x64 && x5 && x18 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && ~x64 && x5 && ~x18 && x1 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && ~x64 && x5 && ~x18 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && ~x64 && ~x5 && x2 && x1 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && ~x64 && ~x5 && x2 && ~x1 )
						nx_state = s1;
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && ~x64 && ~x5 && ~x2 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s22;
						end
					else if( x67 && x66 && ~x65 && ~x68 && ~x62 && ~x63 && ~x64 && ~x5 && ~x2 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && x65 && x68 && x21 && x7 && x1 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x67 && ~x66 && x65 && x68 && x21 && x7 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && x65 && x68 && x21 && ~x7 && x11 && x2 && x1 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s28;
						end
					else if( x67 && ~x66 && x65 && x68 && x21 && ~x7 && x11 && x2 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && x65 && x68 && x21 && ~x7 && x11 && ~x2 && x1 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x67 && ~x66 && x65 && x68 && x21 && ~x7 && x11 && ~x2 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && x65 && x68 && x21 && ~x7 && ~x11 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x67 && ~x66 && x65 && x68 && x21 && ~x7 && ~x11 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && x65 && x68 && ~x21 && x22 && x23 && x9 && x1 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x67 && ~x66 && x65 && x68 && ~x21 && x22 && x23 && x9 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && x65 && x68 && ~x21 && x22 && x23 && ~x9 && x2 && x3 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s31;
						end
					else if( x67 && ~x66 && x65 && x68 && ~x21 && x22 && x23 && ~x9 && x2 && x3 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && x65 && x68 && ~x21 && x22 && x23 && ~x9 && x2 && ~x3 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x67 && ~x66 && x65 && x68 && ~x21 && x22 && x23 && ~x9 && x2 && ~x3 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && x65 && x68 && ~x21 && x22 && x23 && ~x9 && ~x2 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s32;
						end
					else if( x67 && ~x66 && x65 && x68 && ~x21 && x22 && x23 && ~x9 && ~x2 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && x65 && x68 && ~x21 && x22 && ~x23 && x4 && x7 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x67 && ~x66 && x65 && x68 && ~x21 && x22 && ~x23 && x4 && ~x7 && x2 && x1 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s33;
						end
					else if( x67 && ~x66 && x65 && x68 && ~x21 && x22 && ~x23 && x4 && ~x7 && x2 && ~x1 )
						begin
							y3 = 1'b1;	y12 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s34;
						end
					else if( x67 && ~x66 && x65 && x68 && ~x21 && x22 && ~x23 && x4 && ~x7 && ~x2 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s35;
						end
					else if( x67 && ~x66 && x65 && x68 && ~x21 && x22 && ~x23 && ~x4 )
						nx_state = s1;
					else if( x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && x23 && x7 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && x23 && x7 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && x23 && ~x7 && x2 && x8 && x1 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s36;
						end
					else if( x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && x23 && ~x7 && x2 && x8 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && x23 && ~x7 && x2 && ~x8 && x1 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s33;
						end
					else if( x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && x23 && ~x7 && x2 && ~x8 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && x23 && ~x7 && ~x2 && x1 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && x23 && ~x7 && ~x2 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && ~x23 && x9 && x1 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && ~x23 && x9 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && ~x23 && ~x9 && x2 && x3 && x1 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s31;
						end
					else if( x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && ~x23 && ~x9 && x2 && x3 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && ~x23 && ~x9 && x2 && ~x3 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && ~x23 && ~x9 && x2 && ~x3 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && ~x23 && ~x9 && ~x2 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s32;
						end
					else if( x67 && ~x66 && x65 && x68 && ~x21 && ~x22 && ~x23 && ~x9 && ~x2 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && x65 && ~x68 && x9 && x1 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	y12 = 1'b1;	
							nx_state = s37;
						end
					else if( x67 && ~x66 && x65 && ~x68 && x9 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && x65 && ~x68 && ~x9 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s38;
						end
					else if( x67 && ~x66 && x65 && ~x68 && ~x9 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && x68 && x20 && x4 && x19 && x2 )
						nx_state = s39;
					else if( x67 && ~x66 && ~x65 && x68 && x20 && x4 && x19 && ~x2 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && x68 && x20 && x4 && ~x19 && x2 )
						nx_state = s40;
					else if( x67 && ~x66 && ~x65 && x68 && x20 && x4 && ~x19 && ~x2 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && x68 && x20 && ~x4 && x3 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							nx_state = s41;
						end
					else if( x67 && ~x66 && ~x65 && x68 && x20 && ~x4 && x3 && ~x2 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && x68 && x20 && ~x4 && ~x3 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x67 && ~x66 && ~x65 && x68 && x20 && ~x4 && ~x3 && ~x2 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && x68 && ~x20 && x21 && x4 && x19 && x1 )
						begin
							y3 = 1'b1;	y20 = 1'b1;	
							nx_state = s42;
						end
					else if( x67 && ~x66 && ~x65 && x68 && ~x20 && x21 && x4 && x19 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && x68 && ~x20 && x21 && x4 && ~x19 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( x67 && ~x66 && ~x65 && x68 && ~x20 && x21 && x4 && ~x19 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && x68 && ~x20 && x21 && ~x4 && x5 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s44;
						end
					else if( x67 && ~x66 && ~x65 && x68 && ~x20 && x21 && ~x4 && x5 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && x68 && ~x20 && x21 && ~x4 && ~x5 && x1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( x67 && ~x66 && ~x65 && x68 && ~x20 && x21 && ~x4 && ~x5 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x5 && x1 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( x67 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && x5 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x5 && x4 && x1 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y21 = 1'b1;	
							nx_state = s45;
						end
					else if( x67 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x5 && x4 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x5 && ~x4 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s44;
						end
					else if( x67 && ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x5 && ~x4 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && ~x68 && x24 && x26 && x6 && x1 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s46;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && x24 && x26 && x6 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && ~x68 && x24 && x26 && ~x6 && x5 && x1 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && x24 && x26 && ~x6 && x5 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && ~x68 && x24 && x26 && ~x6 && ~x5 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && x24 && x26 && ~x6 && ~x5 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && ~x68 && x24 && ~x26 && x5 && x18 && x1 )
						begin
							y14 = 1'b1;	
							nx_state = s48;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && x24 && ~x26 && x5 && x18 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && ~x68 && x24 && ~x26 && x5 && ~x18 && x1 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s49;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && x24 && ~x26 && x5 && ~x18 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && ~x68 && x24 && ~x26 && ~x5 && x2 && x1 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s50;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && x24 && ~x26 && ~x5 && x2 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && ~x68 && x24 && ~x26 && ~x5 && ~x2 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && x24 && ~x26 && ~x5 && ~x2 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && x26 && x6 && x2 && x17 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s50;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && x26 && x6 && x2 && ~x17 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s46;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && x26 && x6 && ~x2 && x5 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s51;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && x26 && x6 && ~x2 && ~x5 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s19;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && x26 && ~x6 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x3 && x17 && x1 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x3 && x17 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x3 && ~x17 && x1 )
						begin
							y14 = 1'b1;	
							nx_state = s48;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x3 && ~x17 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && ~x3 && x4 && x1 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && ~x3 && x4 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && ~x3 && ~x4 && x1 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && ~x3 && ~x4 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && x6 && x1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && x6 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && ~x6 && x5 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && ~x6 && x5 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && ~x6 && ~x5 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && ~x6 && ~x5 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && ~x26 && x6 && x19 && x1 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && ~x26 && x6 && x19 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && ~x26 && x6 && ~x19 && x1 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && ~x26 && x6 && ~x19 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && ~x26 && ~x6 && x2 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && ~x26 && ~x6 && x2 && ~x1 )
						nx_state = s1;
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && ~x26 && ~x6 && ~x2 && x1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( x67 && ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && ~x26 && ~x6 && ~x2 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && x68 && x1 && x21 && x20 && x3 && x19 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x67 && x66 && x65 && x68 && x1 && x21 && x20 && x3 && ~x19 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s57;
						end
					else if( ~x67 && x66 && x65 && x68 && x1 && x21 && x20 && ~x3 && x4 )
						begin
							y22 = 1'b1;	
							nx_state = s58;
						end
					else if( ~x67 && x66 && x65 && x68 && x1 && x21 && x20 && ~x3 && ~x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x67 && x66 && x65 && x68 && x1 && x21 && ~x20 && x6 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s58;
						end
					else if( ~x67 && x66 && x65 && x68 && x1 && x21 && ~x20 && x6 && ~x17 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x67 && x66 && x65 && x68 && x1 && x21 && ~x20 && ~x6 && x4 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s60;
						end
					else if( ~x67 && x66 && x65 && x68 && x1 && x21 && ~x20 && ~x6 && ~x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x67 && x66 && x65 && x68 && x1 && ~x21 && x6 && x20 && x17 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x67 && x66 && x65 && x68 && x1 && ~x21 && x6 && x20 && ~x17 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	
							nx_state = s61;
						end
					else if( ~x67 && x66 && x65 && x68 && x1 && ~x21 && x6 && ~x20 && x17 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	
							nx_state = s61;
						end
					else if( ~x67 && x66 && x65 && x68 && x1 && ~x21 && x6 && ~x20 && ~x17 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x67 && x66 && x65 && x68 && x1 && ~x21 && ~x6 && x5 )
						begin
							y22 = 1'b1;	
							nx_state = s58;
						end
					else if( ~x67 && x66 && x65 && x68 && x1 && ~x21 && ~x6 && ~x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x67 && x66 && x65 && x68 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && x61 && x60 && x5 && x4 && x17 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x67 && x66 && x65 && ~x68 && x61 && x60 && x5 && x4 && ~x17 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x67 && x66 && x65 && ~x68 && x61 && x60 && x5 && ~x4 && x6 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y24 = 1'b1;	
							nx_state = s64;
						end
					else if( ~x67 && x66 && x65 && ~x68 && x61 && x60 && x5 && ~x4 && ~x6 )
						begin
							y3 = 1'b1;	
							nx_state = s65;
						end
					else if( ~x67 && x66 && x65 && ~x68 && x61 && x60 && ~x5 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && x62 && x59 && x19 && x1 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && x62 && x59 && x19 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && x62 && x59 && ~x19 && x1 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s67;
						end
					else if( ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && x62 && x59 && ~x19 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && x62 && ~x59 && x6 && x1 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s68;
						end
					else if( ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && x62 && ~x59 && x6 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && x62 && ~x59 && ~x6 && x1 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s69;
						end
					else if( ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && x62 && ~x59 && ~x6 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && ~x62 && x3 && x17 && x1 )
						nx_state = s70;
					else if( ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && ~x62 && x3 && x17 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && ~x62 && x3 && ~x17 && x1 )
						nx_state = s71;
					else if( ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && ~x62 && x3 && ~x17 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && ~x62 && ~x3 && x6 && x1 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && ~x62 && ~x3 && x6 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && ~x62 && ~x3 && ~x6 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( ~x67 && x66 && x65 && ~x68 && x61 && ~x60 && ~x62 && ~x3 && ~x6 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && x60 && x3 && x17 && x1 )
						nx_state = s70;
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && x60 && x3 && x17 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && x60 && x3 && ~x17 && x1 )
						nx_state = s71;
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && x60 && x3 && ~x17 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && x60 && ~x3 && x6 && x1 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && x60 && ~x3 && x6 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && x60 && ~x3 && ~x6 && x1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && x60 && ~x3 && ~x6 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && x62 && x3 && x1 )
						nx_state = s71;
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && x62 && x3 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && x62 && ~x3 && x5 && x1 )
						nx_state = s73;
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && x62 && ~x3 && x5 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && x62 && ~x3 && ~x5 && x15 && x16 && x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s74;
						end
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && x62 && ~x3 && ~x5 && x15 && x16 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && x62 && ~x3 && ~x5 && x15 && ~x16 && x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && x62 && ~x3 && ~x5 && x15 && ~x16 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && x62 && ~x3 && ~x5 && ~x15 && x1 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && x62 && ~x3 && ~x5 && ~x15 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && ~x62 && x6 && x1 )
						nx_state = s71;
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && ~x62 && x6 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && ~x62 && ~x6 && x2 && x1 )
						nx_state = s73;
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && ~x62 && ~x6 && x2 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && ~x62 && ~x6 && ~x2 && x1 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x67 && x66 && x65 && ~x68 && ~x61 && ~x60 && ~x62 && ~x6 && ~x2 && ~x1 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && x1 && x21 && x68 && x3 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x67 && x66 && ~x65 && x1 && x21 && x68 && ~x3 && x18 && x19 )
						begin
							y25 = 1'b1;	y26 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x67 && x66 && ~x65 && x1 && x21 && x68 && ~x3 && x18 && ~x19 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x67 && x66 && ~x65 && x1 && x21 && x68 && ~x3 && ~x18 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s79;
						end
					else if( ~x67 && x66 && ~x65 && x1 && x21 && ~x68 && x6 && x17 )
						nx_state = s40;
					else if( ~x67 && x66 && ~x65 && x1 && x21 && ~x68 && x6 && ~x17 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s80;
						end
					else if( ~x67 && x66 && ~x65 && x1 && x21 && ~x68 && ~x6 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s81;
						end
					else if( ~x67 && x66 && ~x65 && x1 && x21 && ~x68 && ~x6 && ~x2 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x67 && x66 && ~x65 && x1 && ~x21 && x22 && x68 && x3 )
						begin
							y8 = 1'b1;	y18 = 1'b1;	
							nx_state = s82;
						end
					else if( ~x67 && x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x3 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && x23 && x5 && x19 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x67 && x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && x23 && x5 && ~x19 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y13 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x67 && x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && x23 && ~x5 && x6 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s84;
						end
					else if( ~x67 && x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && x23 && ~x5 && ~x6 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x67 && x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && ~x23 && x4 && x17 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x67 && x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && ~x23 && x4 && ~x17 )
						begin
							y1 = 1'b1;	
							nx_state = s22;
						end
					else if( ~x67 && x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && ~x23 && ~x4 && x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x67 && x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && ~x23 && ~x4 && ~x5 )
						begin
							y2 = 1'b1;	
							nx_state = s85;
						end
					else if( ~x67 && x66 && ~x65 && x1 && ~x21 && ~x22 && x68 && x9 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s28;
						end
					else if( ~x67 && x66 && ~x65 && x1 && ~x21 && ~x22 && x68 && ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x67 && x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x5 && x17 )
						begin
							y1 = 1'b1;	
							nx_state = s22;
						end
					else if( ~x67 && x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x5 && ~x17 && x23 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x67 && x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x5 && ~x17 && ~x23 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x67 && x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && ~x5 && x6 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x67 && x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && ~x5 && ~x6 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x67 && x66 && ~x65 && ~x1 && x22 && x19 && x20 && x21 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && x22 && x19 && x20 && ~x21 && x68 && x3 )
						begin
							y25 = 1'b1;	y26 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x67 && x66 && ~x65 && ~x1 && x22 && x19 && x20 && ~x21 && x68 && ~x3 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && x22 && x19 && x20 && ~x21 && ~x68 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && x22 && x19 && ~x20 && x21 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && x22 && x19 && ~x20 && ~x21 && x68 && x3 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x67 && x66 && ~x65 && ~x1 && x22 && x19 && ~x20 && ~x21 && x68 && ~x3 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && x22 && x19 && ~x20 && ~x21 && ~x68 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && x22 && ~x19 && x21 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && x22 && ~x19 && ~x21 && x68 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x67 && x66 && ~x65 && ~x1 && x22 && ~x19 && ~x21 && x68 && ~x3 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && x22 && ~x19 && ~x21 && ~x68 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && x21 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && x17 && x10 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && x17 && ~x10 && x68 && x16 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && x17 && ~x10 && x68 && ~x16 && x15 && x14 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && x17 && ~x10 && x68 && ~x16 && x15 && ~x14 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && x17 && ~x10 && x68 && ~x16 && x15 && ~x14 && ~x3 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && x17 && ~x10 && x68 && ~x16 && ~x15 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && x17 && ~x10 && x68 && ~x16 && ~x15 && ~x3 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && x17 && ~x10 && ~x68 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && x14 && x68 && x16 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && x14 && x68 && x16 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && x14 && x68 && x16 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && x14 && x68 && ~x16 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && x14 && ~x68 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && x15 && x16 && x10 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && x15 && x16 && ~x10 && x68 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && x15 && x16 && ~x10 && x68 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && x15 && x16 && ~x10 && x68 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && x15 && x16 && ~x10 && x68 && ~x4 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && x15 && x16 && ~x10 && ~x68 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && x15 && ~x16 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && ~x15 && x68 && x16 && x10 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && ~x15 && x68 && x16 && ~x10 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && ~x15 && x68 && x16 && ~x10 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && ~x15 && x68 && x16 && ~x10 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && ~x15 && x68 && ~x16 )
						nx_state = s1;
					else if( ~x67 && x66 && ~x65 && ~x1 && ~x22 && ~x21 && ~x17 && ~x14 && ~x15 && ~x68 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && x68 && x10 && x1 )
						begin
							y28 = 1'b1;	y29 = 1'b1;	
							nx_state = s90;
						end
					else if( ~x67 && ~x66 && x65 && x68 && x10 && ~x1 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && x68 && ~x10 && x1 )
						begin
							y3 = 1'b1;	
							nx_state = s65;
						end
					else if( ~x67 && ~x66 && x65 && x68 && ~x10 && ~x1 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && x21 && x4 && x20 && x1 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && x21 && x4 && x20 && ~x1 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && x21 && x4 && ~x20 && x18 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && x21 && x4 && ~x20 && ~x18 && x1 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && x21 && x4 && ~x20 && ~x18 && ~x1 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && x21 && ~x4 && x3 && x1 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && x21 && ~x4 && x3 && ~x1 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && x21 && ~x4 && ~x3 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && x21 && ~x4 && ~x3 && ~x1 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && x2 && x20 && x23 && x1 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && x2 && x20 && x23 && ~x1 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && x2 && x20 && ~x23 )
						begin
							y28 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && x2 && ~x20 && x23 && x19 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && x2 && ~x20 && x23 && ~x19 && x1 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && x2 && ~x20 && x23 && ~x19 && ~x1 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && x2 && ~x20 && ~x23 && x4 && x19 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && x2 && ~x20 && ~x23 && x4 && ~x19 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && x2 && ~x20 && ~x23 && ~x4 && x3 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && x2 && ~x20 && ~x23 && ~x4 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x2 && x3 && x23 && x1 )
						begin
							y31 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x2 && x3 && x23 && ~x1 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x2 && x3 && ~x23 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x2 && ~x3 && x23 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x2 && ~x3 && x23 && ~x1 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && x22 && ~x2 && ~x3 && ~x23 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && x19 && x23 && x1 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && x19 && x23 && ~x1 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && x19 && ~x23 && x1 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							nx_state = s97;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && x19 && ~x23 && ~x1 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && x4 && x23 && x18 && x1 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && x4 && x23 && x18 && ~x1 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && x4 && x23 && ~x18 && x1 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							nx_state = s97;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && x4 && x23 && ~x18 && ~x1 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && x4 && ~x23 && x20 && x1 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s98;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && x4 && ~x23 && x20 && ~x1 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && x4 && ~x23 && ~x20 && x1 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && x4 && ~x23 && ~x20 && ~x1 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && ~x4 && x3 && x23 && x1 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && ~x4 && x3 && x23 && ~x1 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && ~x4 && x3 && ~x23 && x1 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && ~x4 && x3 && ~x23 && ~x1 )
						nx_state = s1;
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && ~x4 && ~x3 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x67 && ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x19 && ~x4 && ~x3 && ~x1 )
						nx_state = s1;
					else if( ~x67 && ~x66 && ~x65 && x1 && x21 && x68 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && x21 && x68 && ~x6 && x10 && x11 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s102;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && x21 && x68 && ~x6 && x10 && ~x11 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && x21 && x68 && ~x6 && ~x10 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && x21 && ~x68 && x10 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && x21 && ~x68 && ~x10 && x12 && x11 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && x21 && ~x68 && ~x10 && x12 && ~x11 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && x21 && ~x68 && ~x10 && ~x12 && x2 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && x21 && ~x68 && ~x10 && ~x12 && ~x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && x9 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s105;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && x10 && x18 && x19 && x11 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && x10 && x18 && x19 && ~x11 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s102;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && x10 && x18 && ~x19 && x12 && x16 && x11 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && x10 && x18 && ~x19 && x12 && x16 && ~x11 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s102;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && x10 && x18 && ~x19 && x12 && ~x16 && x11 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s102;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && x10 && x18 && ~x19 && x12 && ~x16 && ~x11 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && x10 && x18 && ~x19 && ~x12 && x11 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && x10 && x18 && ~x19 && ~x12 && ~x11 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s102;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && x10 && ~x18 && x11 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s102;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && x10 && ~x18 && ~x11 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && x68 && ~x9 && ~x10 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && x3 )
						begin
							y8 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s106;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && ~x3 && x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y9 = 1'b1;	
							nx_state = s107;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && ~x3 && x11 && ~x2 )
						nx_state = s40;
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && ~x3 && ~x11 && x9 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && x22 && ~x68 && ~x3 && ~x11 && ~x9 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && x68 && x11 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && x68 && ~x11 )
						nx_state = s1;
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && x20 && x13 && x9 && x11 )
						nx_state = s40;
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && x20 && x13 && x9 && ~x11 && x2 )
						nx_state = s1;
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && x20 && x13 && x9 && ~x11 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && x20 && x13 && ~x9 && x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && x20 && x13 && ~x9 && ~x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && x20 && ~x13 && x2 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && x20 && ~x13 && ~x2 && x9 && x11 )
						nx_state = s40;
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && x20 && ~x13 && ~x2 && x9 && ~x11 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && x20 && ~x13 && ~x2 && ~x9 && x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && x20 && ~x13 && ~x2 && ~x9 && ~x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && ~x20 && x2 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && ~x20 && ~x2 && x9 && x11 )
						nx_state = s40;
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && ~x20 && ~x2 && x9 && ~x11 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && ~x20 && ~x2 && ~x9 && x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && x19 && ~x20 && ~x2 && ~x9 && ~x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && ~x19 && x2 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && ~x19 && ~x2 && x9 && x11 )
						nx_state = s40;
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && ~x19 && ~x2 && x9 && ~x11 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && ~x19 && ~x2 && ~x9 && x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x67 && ~x66 && ~x65 && x1 && ~x21 && ~x22 && ~x68 && ~x19 && ~x2 && ~x9 && ~x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x67 && ~x66 && ~x65 && ~x1 && x68 && x22 )
						nx_state = s1;
					else if( ~x67 && ~x66 && ~x65 && ~x1 && x68 && ~x22 && x21 )
						nx_state = s1;
					else if( ~x67 && ~x66 && ~x65 && ~x1 && x68 && ~x22 && ~x21 && x11 && x3 && x6 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x67 && ~x66 && ~x65 && ~x1 && x68 && ~x22 && ~x21 && x11 && x3 && ~x6 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x67 && ~x66 && ~x65 && ~x1 && x68 && ~x22 && ~x21 && x11 && ~x3 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x67 && ~x66 && ~x65 && ~x1 && x68 && ~x22 && ~x21 && ~x11 )
						nx_state = s1;
					else if( ~x67 && ~x66 && ~x65 && ~x1 && ~x68 )
						nx_state = s1;
					else nx_state = s1;
				s2 : if( x22 )
						nx_state = s1;
					else if( ~x22 && x15 && x8 )
						begin
							y11 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x22 && x15 && ~x8 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s111;
						end
					else if( ~x22 && ~x15 && x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x22 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else nx_state = s2;
				s3 : if( x65 )
						nx_state = s1;
					else if( ~x65 && x21 && x16 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s113;
						end
					else if( ~x65 && x21 && x16 && ~x10 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && x21 && ~x16 )
						begin
							y5 = 1'b1;	y17 = 1'b1;	
							nx_state = s115;
						end
					else if( ~x65 && ~x21 )
						nx_state = s1;
					else nx_state = s3;
				s4 : if( x65 && x67 && x66 && x22 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y10 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s9;
						end
					else if( x65 && x67 && x66 && ~x22 && x23 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y10 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s9;
						end
					else if( x65 && x67 && x66 && ~x22 && ~x23 )
						nx_state = s1;
					else if( x65 && x67 && ~x66 && x21 && x18 )
						begin
							y14 = 1'b1;	y19 = 1'b1;	
							nx_state = s116;
						end
					else if( x65 && x67 && ~x66 && x21 && ~x18 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s117;
						end
					else if( x65 && x67 && ~x66 && ~x21 && x22 && x8 && x23 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x66 && ~x21 && x22 && x8 && x23 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x66 && ~x21 && x22 && x8 && x23 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && x67 && ~x66 && ~x21 && x22 && x8 && ~x23 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x66 && ~x21 && x22 && x8 && ~x23 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x66 && ~x21 && x22 && x8 && ~x23 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x65 && x67 && ~x66 && ~x21 && x22 && ~x8 )
						nx_state = s1;
					else if( x65 && x67 && ~x66 && ~x21 && ~x22 && x23 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x66 && ~x21 && ~x22 && x23 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x66 && ~x21 && ~x22 && x23 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && x67 && ~x66 && ~x21 && ~x22 && x23 && ~x9 )
						nx_state = s1;
					else if( x65 && x67 && ~x66 && ~x21 && ~x22 && ~x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x66 && ~x21 && ~x22 && ~x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x66 && ~x21 && ~x22 && ~x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && x67 && ~x66 && ~x21 && ~x22 && ~x23 && ~x8 )
						nx_state = s1;
					else if( x65 && ~x67 && x66 && x68 )
						nx_state = s1;
					else if( x65 && ~x67 && x66 && ~x68 && x61 && x60 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x67 && x66 && ~x68 && x61 && x60 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x67 && x66 && ~x68 && x61 && x60 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && ~x67 && x66 && ~x68 && x61 && x60 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && ~x67 && x66 && ~x68 && x61 && ~x60 && x62 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x67 && x66 && ~x68 && x61 && ~x60 && ~x62 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s118;
						end
					else if( x65 && ~x67 && x66 && ~x68 && ~x61 && x60 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s118;
						end
					else if( x65 && ~x67 && x66 && ~x68 && ~x61 && ~x60 )
						nx_state = s40;
					else if( x65 && ~x67 && ~x66 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x65 && ~x67 && ~x66 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x67 && ~x66 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x67 && ~x66 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x66 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x66 && ~x21 && x23 && x22 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( x65 && ~x67 && ~x66 && ~x21 && x23 && x22 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x67 && ~x66 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x67 && ~x66 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x66 && ~x21 && x23 && x22 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x66 && ~x21 && x23 && ~x22 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x67 && ~x66 && ~x21 && x23 && ~x22 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x67 && ~x66 && ~x21 && x23 && ~x22 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x66 && ~x21 && x23 && ~x22 && ~x20 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x66 && ~x21 && ~x23 && x18 && x14 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x67 && ~x66 && ~x21 && ~x23 && x18 && x14 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x67 && ~x66 && ~x21 && ~x23 && x18 && ~x14 && x13 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x67 && ~x66 && ~x21 && ~x23 && x18 && ~x14 && x13 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x67 && ~x66 && ~x21 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x66 && ~x21 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x68 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && x68 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && x68 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && x68 && x21 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x68 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x65 && x68 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x65 && x68 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && x68 && ~x21 && ~x20 )
						nx_state = s1;
					else if( ~x65 && ~x68 && x62 )
						nx_state = s1;
					else if( ~x65 && ~x68 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && ~x68 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x68 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x68 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x68 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x68 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x68 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else nx_state = s4;
				s5 : if( x65 && x22 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x65 && ~x22 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s121;
						end
					else if( ~x65 && x21 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && ~x21 && x23 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x65 && ~x21 && ~x23 && x22 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x21 && ~x23 && ~x22 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else nx_state = s5;
				s6 : if( x22 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	
							nx_state = s111;
						end
					else if( ~x22 )
						nx_state = s1;
					else nx_state = s6;
				s7 : if( x65 && x67 && x66 && x22 )
						nx_state = s1;
					else if( x65 && x67 && x66 && ~x22 && x23 && x19 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x65 && x67 && x66 && ~x22 && x23 && x19 && x15 && ~x8 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x65 && x67 && x66 && ~x22 && x23 && x19 && ~x15 && x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x67 && x66 && ~x22 && x23 && x19 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s122;
						end
					else if( x65 && x67 && x66 && ~x22 && x23 && ~x19 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x67 && x66 && ~x22 && ~x23 )
						nx_state = s1;
					else if( x65 && x67 && ~x66 && x21 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x65 && x67 && ~x66 && ~x21 )
						nx_state = s1;
					else if( x65 && ~x67 && x66 && x68 && x20 )
						nx_state = s1;
					else if( x65 && ~x67 && x66 && x68 && ~x20 && x21 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && ~x67 && x66 && x68 && ~x20 && x21 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && ~x67 && x66 && x68 && ~x20 && x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && x66 && x68 && ~x20 && x21 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x67 && x66 && x68 && ~x20 && ~x21 )
						nx_state = s1;
					else if( x65 && ~x67 && x66 && ~x68 && x60 && x61 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x67 && x66 && ~x68 && x60 && x61 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x67 && x66 && ~x68 && x60 && x61 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && ~x67 && x66 && ~x68 && x60 && x61 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && ~x67 && x66 && ~x68 && x60 && ~x61 )
						nx_state = s39;
					else if( x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && x62 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && ~x62 )
						nx_state = s39;
					else if( x65 && ~x67 && x66 && ~x68 && ~x60 && ~x61 )
						nx_state = s40;
					else if( x65 && ~x67 && ~x66 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x65 && ~x67 && ~x66 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x67 && ~x66 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x67 && ~x66 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x66 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x66 && ~x21 && x23 && x22 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( x65 && ~x67 && ~x66 && ~x21 && x23 && x22 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x67 && ~x66 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x67 && ~x66 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x66 && ~x21 && x23 && x22 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x66 && ~x21 && x23 && ~x22 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x67 && ~x66 && ~x21 && x23 && ~x22 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x67 && ~x66 && ~x21 && x23 && ~x22 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x66 && ~x21 && x23 && ~x22 && ~x20 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x66 && ~x21 && ~x23 && x18 && x14 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x67 && ~x66 && ~x21 && ~x23 && x18 && x14 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x67 && ~x66 && ~x21 && ~x23 && x18 && ~x14 && x13 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x67 && ~x66 && ~x21 && ~x23 && x18 && ~x14 && x13 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x67 && ~x66 && ~x21 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x66 && ~x21 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x66 && x68 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && x66 && x68 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && x66 && x68 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && x66 && x68 && x21 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && x68 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x65 && x66 && x68 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x65 && x66 && x68 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && x66 && x68 && ~x21 && ~x20 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x68 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x21 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x21 && x22 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x65 && ~x66 && ~x21 && ~x22 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s123;
						end
					else nx_state = s7;
				s8 : if( x65 && x23 )
						begin
							y2 = 1'b1;	y16 = 1'b1;	y24 = 1'b1;	
							nx_state = s124;
						end
					else if( x65 && ~x23 && x18 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && ~x23 && x18 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && ~x23 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && ~x9 )
						nx_state = s1;
					else nx_state = s8;
				s9 : if( x22 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s125;
						end
					else if( ~x22 && x23 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( ~x22 && x23 && x15 && ~x8 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x22 && x23 && ~x15 && x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x22 && x23 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s122;
						end
					else if( ~x22 && ~x23 )
						begin
							y2 = 1'b1;	y16 = 1'b1;	y24 = 1'b1;	
							nx_state = s124;
						end
					else nx_state = s9;
				s10 : if( x65 && x66 && x67 && x22 && x16 && x15 && x8 && x14 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && x66 && x67 && x22 && x16 && x15 && x8 && ~x14 && x7 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s126;
						end
					else if( x65 && x66 && x67 && x22 && x16 && x15 && x8 && ~x14 && ~x7 && x12 )
						begin
							y2 = 1'b1;	
							nx_state = s85;
						end
					else if( x65 && x66 && x67 && x22 && x16 && x15 && x8 && ~x14 && ~x7 && ~x12 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && x67 && x22 && x16 && x15 && x8 && ~x14 && ~x7 && ~x12 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && x67 && x22 && x16 && x15 && x8 && ~x14 && ~x7 && ~x12 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && x66 && x67 && x22 && x16 && x15 && x8 && ~x14 && ~x7 && ~x12 && ~x17 )
						nx_state = s1;
					else if( x65 && x66 && x67 && x22 && x16 && x15 && ~x8 && x14 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( x65 && x66 && x67 && x22 && x16 && x15 && ~x8 && ~x14 && x7 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s127;
						end
					else if( x65 && x66 && x67 && x22 && x16 && x15 && ~x8 && ~x14 && ~x7 && x13 )
						begin
							y2 = 1'b1;	
							nx_state = s85;
						end
					else if( x65 && x66 && x67 && x22 && x16 && x15 && ~x8 && ~x14 && ~x7 && ~x13 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && x67 && x22 && x16 && x15 && ~x8 && ~x14 && ~x7 && ~x13 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && x67 && x22 && x16 && x15 && ~x8 && ~x14 && ~x7 && ~x13 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && x66 && x67 && x22 && x16 && x15 && ~x8 && ~x14 && ~x7 && ~x13 && ~x17 )
						nx_state = s1;
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && x8 && x9 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && x8 && x9 && ~x2 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && x8 && x9 && ~x2 && ~x4 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s111;
						end
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && x8 && ~x9 && x7 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && x8 && ~x9 && x7 && ~x2 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && x8 && ~x9 && x7 && ~x2 && ~x4 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s111;
						end
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && x8 && ~x9 && ~x7 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && x8 && ~x9 && ~x7 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && x8 && ~x9 && ~x7 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && x8 && ~x9 && ~x7 && ~x17 )
						nx_state = s1;
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && x7 && x11 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && x7 && x11 && ~x2 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && x7 && x11 && ~x2 && ~x4 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s111;
						end
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && x7 && ~x11 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && x7 && ~x11 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && x7 && ~x11 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && x7 && ~x11 && ~x17 )
						nx_state = s1;
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && ~x7 && x10 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && ~x7 && x10 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && ~x7 && x10 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && ~x7 && x10 && ~x17 )
						nx_state = s1;
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x2 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x65 && x66 && x67 && x22 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x2 && ~x4 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s111;
						end
					else if( x65 && x66 && x67 && x22 && ~x16 && x15 && x7 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x65 && x66 && x67 && x22 && ~x16 && x15 && ~x7 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( x65 && x66 && x67 && x22 && ~x16 && x15 && ~x7 && ~x2 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x65 && x66 && x67 && x22 && ~x16 && x15 && ~x7 && ~x2 && ~x4 && x8 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y28 = 1'b1;	
							nx_state = s129;
						end
					else if( x65 && x66 && x67 && x22 && ~x16 && x15 && ~x7 && ~x2 && ~x4 && ~x8 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s111;
						end
					else if( x65 && x66 && x67 && x22 && ~x16 && ~x15 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( x65 && x66 && x67 && x22 && ~x16 && ~x15 && ~x2 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x65 && x66 && x67 && x22 && ~x16 && ~x15 && ~x2 && ~x4 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( x65 && x66 && x67 && ~x22 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( x65 && x66 && ~x67 && x21 && x20 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s131;
						end
					else if( x65 && x66 && ~x67 && x21 && ~x20 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s132;
						end
					else if( x65 && x66 && ~x67 && ~x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s132;
						end
					else if( x65 && ~x66 && x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s32;
						end
					else if( x65 && ~x66 && ~x21 && x23 && x22 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x23 && ~x22 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s31;
						end
					else if( x65 && ~x66 && ~x21 && ~x23 && x22 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s32;
						end
					else if( x65 && ~x66 && ~x21 && ~x23 && ~x22 )
						nx_state = s1;
					else if( ~x65 && x20 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x20 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else nx_state = s10;
				s11 : if( x65 && x66 && x60 && x61 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x66 && x60 && x61 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x66 && x60 && x61 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x66 && x60 && x61 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x66 && x60 && ~x61 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && x60 && ~x61 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && x60 && ~x61 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x65 && x66 && x60 && ~x61 && ~x18 )
						nx_state = s39;
					else if( x65 && x66 && ~x60 && x61 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x66 && ~x60 && x61 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x66 && ~x60 && x61 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x65 && x66 && ~x60 && x61 && x62 && ~x18 )
						nx_state = s1;
					else if( x65 && x66 && ~x60 && x61 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && ~x60 && x61 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && ~x60 && x61 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x65 && x66 && ~x60 && x61 && ~x62 && ~x18 )
						nx_state = s39;
					else if( x65 && x66 && ~x60 && ~x61 )
						nx_state = s40;
					else if( x65 && ~x66 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x65 && ~x66 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x23 && x22 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( x65 && ~x66 && ~x21 && x23 && x22 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x66 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x66 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x23 && x22 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x23 && ~x22 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x66 && ~x21 && x23 && ~x22 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x66 && ~x21 && x23 && ~x22 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x23 && ~x22 && ~x20 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x23 && x18 && x14 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x21 && ~x23 && x18 && x14 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x66 && ~x21 && ~x23 && x18 && ~x14 && x13 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x21 && ~x23 && x18 && ~x14 && x13 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x66 && ~x21 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x68 && x5 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && x68 && x5 && ~x18 && x21 && x6 )
						nx_state = s11;
					else if( ~x65 && x68 && x5 && ~x18 && x21 && ~x6 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x65 && x68 && x5 && ~x18 && ~x21 && x4 )
						nx_state = s11;
					else if( ~x65 && x68 && x5 && ~x18 && ~x21 && ~x4 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x65 && x68 && ~x5 && x21 && x4 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x65 && x68 && ~x5 && x21 && ~x4 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s15;
						end
					else if( ~x65 && x68 && ~x5 && ~x21 && x6 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x65 && x68 && ~x5 && ~x21 && ~x6 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s15;
						end
					else if( ~x65 && ~x68 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && ~x68 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && ~x68 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x68 && x62 && ~x61 )
						nx_state = s1;
					else if( ~x65 && ~x68 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && ~x68 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x68 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x68 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x68 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x68 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x68 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else nx_state = s11;
				s12 : if( x65 && x67 && x66 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && x66 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && x66 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && x67 && x66 && x22 && ~x17 )
						nx_state = s1;
					else if( x65 && x67 && x66 && ~x22 && x3 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && x66 && ~x22 && ~x3 && x19 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x65 && x67 && x66 && ~x22 && ~x3 && x19 && x15 && ~x8 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x65 && x67 && x66 && ~x22 && ~x3 && x19 && ~x15 && x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x67 && x66 && ~x22 && ~x3 && x19 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s122;
						end
					else if( x65 && x67 && x66 && ~x22 && ~x3 && ~x19 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x67 && ~x66 )
						nx_state = s1;
					else if( x65 && ~x67 && x66 && x68 && x20 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x67 && x66 && x68 && x20 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x67 && x66 && x68 && x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && x66 && x68 && x20 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x67 && x66 && x68 && ~x20 && x21 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x65 && ~x67 && x66 && x68 && ~x20 && ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x67 && x66 && x68 && ~x20 && ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x67 && x66 && x68 && ~x20 && ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && x66 && x68 && ~x20 && ~x21 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x67 && x66 && ~x68 && x60 && x61 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x67 && x66 && ~x68 && x60 && x61 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x67 && x66 && ~x68 && x60 && x61 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && ~x67 && x66 && ~x68 && x60 && x61 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && ~x67 && x66 && ~x68 && x60 && ~x61 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x67 && x66 && ~x68 && x60 && ~x61 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x67 && x66 && ~x68 && x60 && ~x61 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x65 && ~x67 && x66 && ~x68 && x60 && ~x61 && ~x18 )
						nx_state = s39;
					else if( x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && x62 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x65 && ~x67 && x66 && ~x68 && ~x60 && x61 && ~x62 && ~x18 )
						nx_state = s39;
					else if( x65 && ~x67 && x66 && ~x68 && ~x60 && ~x61 )
						nx_state = s40;
					else if( x65 && ~x67 && ~x66 && x21 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x66 && ~x21 && x19 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x67 && ~x66 && ~x21 && x19 && ~x18 )
						nx_state = s12;
					else if( x65 && ~x67 && ~x66 && ~x21 && ~x19 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							nx_state = s97;
						end
					else if( ~x65 && x68 && x21 && x6 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && x68 && x21 && x6 && ~x18 )
						nx_state = s12;
					else if( ~x65 && x68 && x21 && ~x6 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x65 && x68 && ~x21 && x4 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && x68 && ~x21 && x4 && ~x18 )
						nx_state = s12;
					else if( ~x65 && x68 && ~x21 && ~x4 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x65 && ~x68 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && ~x68 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && ~x68 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x68 && x62 && ~x61 )
						nx_state = s1;
					else if( ~x65 && ~x68 && ~x62 && x63 )
						nx_state = s1;
					else if( ~x65 && ~x68 && ~x62 && ~x63 && x64 && x16 && x8 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && ~x68 && ~x62 && ~x63 && x64 && x16 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x68 && ~x62 && ~x63 && x64 && ~x16 && x4 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x65 && ~x68 && ~x62 && ~x63 && x64 && ~x16 && ~x4 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x65 && ~x68 && ~x62 && ~x63 && ~x64 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else nx_state = s12;
				s13 : if( x65 && x67 && x21 && x68 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x65 && x67 && x21 && x68 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x65 && x67 && x21 && x68 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x65 && x67 && x21 && x68 && ~x8 )
						nx_state = s1;
					else if( x65 && x67 && x21 && ~x68 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x67 && x21 && ~x68 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x67 && x21 && ~x68 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && x67 && x21 && ~x68 && ~x4 )
						nx_state = s1;
					else if( x65 && x67 && ~x21 && x68 && x23 && x22 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x21 && x68 && x23 && x22 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x21 && x68 && x23 && x22 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && x67 && ~x21 && x68 && x23 && x22 && ~x8 )
						nx_state = s1;
					else if( x65 && x67 && ~x21 && x68 && x23 && ~x22 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x21 && x68 && x23 && ~x22 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x21 && x68 && x23 && ~x22 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && x67 && ~x21 && x68 && x23 && ~x22 && ~x9 )
						nx_state = s1;
					else if( x65 && x67 && ~x21 && x68 && ~x23 && x8 && x22 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x21 && x68 && ~x23 && x8 && x22 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x21 && x68 && ~x23 && x8 && x22 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x65 && x67 && ~x21 && x68 && ~x23 && x8 && ~x22 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x21 && x68 && ~x23 && x8 && ~x22 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x21 && x68 && ~x23 && x8 && ~x22 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && x67 && ~x21 && x68 && ~x23 && ~x8 )
						nx_state = s1;
					else if( x65 && x67 && ~x21 && ~x68 && x22 && x19 && x18 && x11 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && x67 && ~x21 && ~x68 && x22 && x19 && x18 && ~x11 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x67 && ~x21 && ~x68 && x22 && x19 && x18 && ~x11 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x67 && ~x21 && ~x68 && x22 && x19 && x18 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && x67 && ~x21 && ~x68 && x22 && x19 && x18 && ~x11 && ~x4 )
						nx_state = s1;
					else if( x65 && x67 && ~x21 && ~x68 && x22 && x19 && ~x18 )
						nx_state = s1;
					else if( x65 && x67 && ~x21 && ~x68 && x22 && ~x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x67 && ~x21 && ~x68 && x22 && ~x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x67 && ~x21 && ~x68 && x22 && ~x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && x67 && ~x21 && ~x68 && x22 && ~x19 && ~x4 )
						nx_state = s1;
					else if( x65 && x67 && ~x21 && ~x68 && ~x22 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x67 && ~x21 && ~x68 && ~x22 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x67 && ~x21 && ~x68 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && x67 && ~x21 && ~x68 && ~x22 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x67 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x65 && ~x67 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x67 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x67 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x21 && x23 && x22 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( x65 && ~x67 && ~x21 && x23 && x22 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x67 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x67 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x21 && x23 && x22 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x21 && x23 && ~x22 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x67 && ~x21 && x23 && ~x22 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x67 && ~x21 && x23 && ~x22 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x21 && x23 && ~x22 && ~x20 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x21 && ~x23 && x18 && x14 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x67 && ~x21 && ~x23 && x18 && x14 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x67 && ~x21 && ~x23 && x18 && ~x14 && x13 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x67 && ~x21 && ~x23 && x18 && ~x14 && x13 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x67 && ~x21 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x21 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && x68 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x68 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && x66 && x67 && ~x68 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && x66 && x67 && ~x68 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x68 && x62 && ~x61 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && x21 && x17 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x66 && ~x67 && x21 && x17 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x66 && ~x67 && x21 && x17 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && x21 && ~x17 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && ~x21 && ~x22 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x22 && x21 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x22 && ~x21 && x16 && x12 && x19 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x22 && ~x21 && x16 && x12 && ~x19 && x18 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x65 && ~x66 && x22 && ~x21 && x16 && x12 && ~x19 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x22 && ~x21 && x16 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x22 && ~x21 && ~x16 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x22 )
						nx_state = s1;
					else nx_state = s13;
				s14 : if( x21 )
						begin
							y10 = 1'b1;	
							nx_state = s139;
						end
					else if( ~x21 && x19 && x16 && x10 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s67;
						end
					else if( ~x21 && x19 && x16 && ~x10 )
						begin
							y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s113;
						end
					else if( ~x21 && x19 && ~x16 && x17 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x21 && x19 && ~x16 && ~x17 )
						begin
							y5 = 1'b1;	y17 = 1'b1;	
							nx_state = s115;
						end
					else if( ~x21 && ~x19 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	
							nx_state = s141;
						end
					else nx_state = s14;
				s15 : if( x65 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( ~x65 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	
							nx_state = s142;
						end
					else nx_state = s15;
				s16 : if( x66 && x67 && x65 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && x67 && x65 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && x67 && x65 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x66 && x67 && x65 && x22 && ~x17 )
						nx_state = s1;
					else if( x66 && x67 && x65 && ~x22 && x18 && x13 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x66 && x67 && x65 && ~x22 && x18 && x13 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x67 && x65 && ~x22 && x18 && ~x13 && x12 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x66 && x67 && x65 && ~x22 && x18 && ~x13 && x12 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x67 && x65 && ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x66 && x67 && x65 && ~x22 && ~x18 )
						nx_state = s1;
					else if( x66 && x67 && ~x65 && x68 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && x67 && ~x65 && x68 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && x67 && ~x65 && x68 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x66 && x67 && ~x65 && x68 && x21 && ~x19 )
						nx_state = s1;
					else if( x66 && x67 && ~x65 && x68 && ~x21 )
						begin
							y10 = 1'b1;	
							nx_state = s139;
						end
					else if( x66 && x67 && ~x65 && ~x68 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x66 && x67 && ~x65 && ~x68 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x66 && x67 && ~x65 && ~x68 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x66 && x67 && ~x65 && ~x68 && x62 && ~x61 )
						nx_state = s1;
					else if( x66 && x67 && ~x65 && ~x68 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && x67 && ~x65 && ~x68 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( x66 && x67 && ~x65 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && x67 && ~x65 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( x66 && x67 && ~x65 && ~x68 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x66 && x67 && ~x65 && ~x68 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( x66 && x67 && ~x65 && ~x68 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x66 && x67 && ~x65 && ~x68 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x66 && x67 && ~x65 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x66 && x67 && ~x65 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x66 && x67 && ~x65 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x66 && x67 && ~x65 && ~x68 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else if( x66 && ~x67 && x65 && x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && ~x67 && x65 && x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && ~x67 && x65 && x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && ~x67 && x65 && x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x66 && ~x67 && x65 && x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && ~x67 && x65 && x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && ~x67 && x65 && x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && ~x67 && x65 && x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( x66 && ~x67 && x65 && ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && ~x67 && x65 && ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && ~x67 && x65 && ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && ~x67 && x65 && ~x21 && ~x19 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && x21 && x68 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x66 && ~x67 && ~x65 && x21 && x68 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x66 && ~x67 && ~x65 && x21 && x68 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && x21 && x68 && ~x9 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && x21 && ~x68 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s143;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x68 && x22 && x9 && x7 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x68 && x22 && x9 && ~x7 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && x68 && x22 && ~x9 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && x68 && ~x22 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x68 && ~x22 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x68 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && x68 && ~x22 && ~x4 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x68 && x23 && x22 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x68 && x23 && ~x22 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x68 && x23 && ~x22 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x68 && x23 && ~x22 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x68 && x23 && ~x22 && ~x19 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x68 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x66 && x65 && x21 && x67 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && x21 && x67 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && x21 && x67 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x66 && x65 && x21 && x67 && ~x4 )
						nx_state = s1;
					else if( ~x66 && x65 && x21 && ~x67 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x66 && x65 && x21 && ~x67 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && x21 && ~x67 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && x21 && ~x67 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && x21 && ~x67 && ~x18 && ~x19 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && x67 && x22 && x18 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && ~x21 && x67 && x22 && x18 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && ~x21 && x67 && x22 && x18 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && x67 && x22 && x18 && ~x4 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && x67 && x22 && ~x18 && x10 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x66 && x65 && ~x21 && x67 && x22 && ~x18 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && ~x21 && x67 && x22 && ~x18 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && ~x21 && x67 && x22 && ~x18 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && x67 && x22 && ~x18 && ~x10 && ~x4 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && x67 && ~x22 && x19 && x10 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x66 && x65 && ~x21 && x67 && ~x22 && x19 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && ~x21 && x67 && ~x22 && x19 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && ~x21 && x67 && ~x22 && x19 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && x67 && ~x22 && x19 && ~x10 && ~x4 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && x67 && ~x22 && ~x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && ~x21 && x67 && ~x22 && ~x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && ~x21 && x67 && ~x22 && ~x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && x67 && ~x22 && ~x19 && ~x4 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x67 && x23 && x22 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( ~x66 && x65 && ~x21 && ~x67 && x23 && x22 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( ~x66 && x65 && ~x21 && ~x67 && x23 && x22 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( ~x66 && x65 && ~x21 && ~x67 && x23 && x22 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x67 && x23 && x22 && ~x19 && ~x17 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x67 && x23 && ~x22 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x66 && x65 && ~x21 && ~x67 && ~x23 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x66 && ~x65 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x66 && ~x65 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x66 && ~x65 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x20 && ~x18 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x66 && ~x65 && ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x66 && ~x65 && ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x66 && ~x65 && ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x66 && ~x65 && ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else nx_state = s16;
				s17 : if( x66 && x67 )
						nx_state = s1;
					else if( x66 && ~x67 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x67 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x67 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x4 )
						nx_state = s1;
					else if( ~x66 && x24 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && ~x24 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s150;
						end
					else nx_state = s17;
				s18 : if( x63 && x62 )
						begin
							y34 = 1'b1;	
							nx_state = s21;
						end
					else if( x63 && ~x62 && x15 && x8 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x63 && ~x62 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x63 && ~x62 && ~x15 && x16 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( x63 && ~x62 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x63 )
						begin
							y34 = 1'b1;	
							nx_state = s21;
						end
					else nx_state = s18;
				s19 : if( x66 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( ~x66 && x26 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x66 && ~x26 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else nx_state = s19;
				s20 : if( x64 )
						nx_state = s1;
					else if( ~x64 && x63 && x18 && x15 && x8 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x64 && x63 && x18 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x64 && x63 && x18 && ~x15 && x16 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x64 && x63 && x18 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x64 && x63 && ~x18 )
						begin
							y31 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x64 && ~x63 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else nx_state = s20;
				s21 : if( x63 )
						begin
							y35 = 1'b1;	
							nx_state = s26;
						end
					else if( ~x63 && x62 )
						begin
							y35 = 1'b1;	
							nx_state = s26;
						end
					else if( ~x63 && ~x62 && x64 && x16 && x8 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x63 && ~x62 && x64 && x16 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x63 && ~x62 && x64 && ~x16 && x4 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x63 && ~x62 && x64 && ~x16 && ~x4 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x63 && ~x62 && ~x64 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x63 && ~x62 && ~x64 && x15 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x63 && ~x62 && ~x64 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s151;
						end
					else if( ~x63 && ~x62 && ~x64 && ~x15 && ~x16 && x14 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x63 && ~x62 && ~x64 && ~x15 && ~x16 && ~x14 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s152;
						end
					else nx_state = s21;
				s22 : if( x65 && x21 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( x65 && ~x21 && x22 && x23 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x21 && x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && ~x21 && ~x22 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x67 && x64 && x63 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && x67 && x64 && ~x63 )
						nx_state = s1;
					else if( ~x65 && x67 && ~x64 && x63 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x67 && ~x64 && ~x63 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x65 && ~x67 && x21 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && x23 && x22 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x67 && ~x21 && x23 && x22 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x67 && ~x21 && x23 && x22 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && x23 && x22 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && x23 && ~x22 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && ~x23 )
						nx_state = s1;
					else nx_state = s22;
				s23 : if( x65 && x16 && x11 && x12 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x65 && x16 && x11 && ~x12 && x13 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x65 && x16 && x11 && ~x12 && ~x13 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s154;
						end
					else if( x65 && x16 && ~x11 && x13 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s63;
						end
					else if( x65 && x16 && ~x11 && ~x13 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( x65 && ~x16 && x17 && x11 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x65 && ~x16 && x17 && x11 && ~x13 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( x65 && ~x16 && x17 && ~x11 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x65 && ~x16 && ~x17 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x65 && x66 && x62 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && x66 && ~x62 && x63 && x64 && x17 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && x66 && ~x62 && x63 && x64 && x17 && ~x13 && x12 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && x66 && ~x62 && x63 && x64 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x62 && x63 && x64 && ~x17 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x62 && x63 && ~x64 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && x64 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s152;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && x14 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && x14 && ~x8 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && ~x14 && x7 && x8 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && ~x14 && x7 && ~x8 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && ~x14 && ~x7 && x8 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s65;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && x19 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && x19 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && ~x14 && ~x7 && ~x8 && x13 )
						begin
							y3 = 1'b1;	
							nx_state = s65;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && x19 && x12 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && x19 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && x7 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && x7 && ~x3 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && x7 && ~x3 && ~x4 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && ~x7 && x9 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && ~x7 && x9 && ~x3 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && ~x7 && x9 && ~x3 && ~x4 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && ~x7 && ~x9 && x3 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && ~x7 && ~x9 && ~x3 && x19 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && ~x7 && ~x9 && ~x3 && x19 && ~x13 && x12 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && ~x7 && ~x9 && ~x3 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && x8 && ~x7 && ~x9 && ~x3 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && x7 && x11 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && x7 && x11 && ~x3 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && x7 && x11 && ~x3 && ~x4 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && x7 && ~x11 && x3 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && x7 && ~x11 && ~x3 && x19 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && x7 && ~x11 && ~x3 && x19 && ~x13 && x12 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && x7 && ~x11 && ~x3 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && x7 && ~x11 && ~x3 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && ~x7 && x10 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && ~x7 && x10 && ~x3 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && ~x7 && x10 && ~x3 && ~x4 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && x3 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x3 && x19 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x3 && x19 && ~x13 && x12 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x3 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x3 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && ~x16 && x15 && x7 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s159;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && ~x16 && x15 && ~x7 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && ~x16 && x15 && ~x7 && ~x3 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && ~x16 && x15 && ~x7 && ~x3 && ~x4 && x8 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && ~x16 && x15 && ~x7 && ~x3 && ~x4 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && ~x16 && ~x15 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && ~x16 && ~x15 && ~x3 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && ~x16 && ~x15 && ~x3 && ~x4 && x14 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y28 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x64 && ~x16 && ~x15 && ~x3 && ~x4 && ~x14 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && x26 && x17 && x11 && x13 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && x26 && x17 && x11 && ~x13 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && x26 && x17 && ~x11 && x12 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && x26 && x17 && ~x11 && x12 && ~x13 )
						begin
							y14 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && x26 && x17 && ~x11 && ~x12 && x13 && x14 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s161;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && x26 && x17 && ~x11 && ~x12 && x13 && ~x14 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && x26 && x17 && ~x11 && ~x12 && x13 && ~x14 && x18 && ~x15 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && x16 && x26 && x17 && ~x11 && ~x12 && x13 && ~x14 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && x16 && x26 && x17 && ~x11 && ~x12 && ~x13 && x15 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s161;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && x26 && x17 && ~x11 && ~x12 && ~x13 && ~x15 && x18 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && x26 && x17 && ~x11 && ~x12 && ~x13 && ~x15 && x18 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && x16 && x26 && x17 && ~x11 && ~x12 && ~x13 && ~x15 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && x16 && x26 && ~x17 && x13 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && x26 && ~x17 && ~x13 && x12 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && x26 && ~x17 && ~x13 && ~x12 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && x26 && ~x17 && ~x13 && ~x12 && ~x2 && x11 && x4 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && x26 && ~x17 && ~x13 && ~x12 && ~x2 && x11 && ~x4 )
						begin
							y8 = 1'b1;	y17 = 1'b1;	y23 = 1'b1;	
							nx_state = s164;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && x26 && ~x17 && ~x13 && ~x12 && ~x2 && ~x11 && x4 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && x26 && ~x17 && ~x13 && ~x12 && ~x2 && ~x11 && ~x4 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s165;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && x11 && x13 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && x11 && ~x13 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && ~x11 && x12 && x13 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && ~x11 && x12 && ~x13 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && ~x11 && ~x12 && x13 && x14 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s167;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && ~x11 && ~x12 && x13 && ~x14 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && ~x11 && ~x12 && x13 && ~x14 && x20 && ~x15 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && ~x11 && ~x12 && x13 && ~x14 && ~x20 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && ~x11 && ~x12 && ~x13 && x15 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s167;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && ~x11 && ~x12 && ~x13 && ~x15 && x20 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && ~x11 && ~x12 && ~x13 && ~x15 && x20 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && x17 && ~x11 && ~x12 && ~x13 && ~x15 && ~x20 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && x11 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && x11 && ~x3 && x12 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && x11 && ~x3 && x12 && ~x4 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s169;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && x11 && ~x3 && ~x12 && x13 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && x11 && ~x3 && ~x12 && x13 && ~x4 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s170;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && x11 && ~x3 && ~x12 && ~x13 && x4 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s165;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && x11 && ~x3 && ~x12 && ~x13 && ~x4 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && ~x11 && x13 && x12 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && ~x11 && x13 && ~x12 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s170;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && ~x11 && ~x13 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && ~x11 && ~x13 && ~x12 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && ~x11 && ~x13 && ~x12 && ~x3 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x66 && x67 && x24 && x16 && ~x26 && ~x17 && ~x11 && ~x13 && ~x12 && ~x3 && ~x4 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s171;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && x11 && x9 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && x11 && x9 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && x11 && x9 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && x11 && x9 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && x11 && ~x9 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && x11 && ~x9 && ~x2 && x4 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && x11 && ~x9 && ~x2 && ~x4 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s165;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && ~x11 && x12 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && ~x11 && x12 && ~x2 && x4 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && ~x11 && x12 && ~x2 && ~x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && ~x11 && ~x12 && x8 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && ~x11 && ~x12 && x8 && ~x2 && x4 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && ~x11 && ~x12 && x8 && ~x2 && ~x4 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s165;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && ~x11 && ~x12 && ~x8 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && ~x11 && ~x12 && ~x8 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && ~x11 && ~x12 && ~x8 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && x13 && ~x11 && ~x12 && ~x8 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && x11 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && x11 && ~x2 && x4 )
						begin
							y6 = 1'b1;	
							nx_state = s172;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && x11 && ~x2 && ~x4 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && x12 && x10 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && x12 && x10 && ~x2 && x4 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && x12 && x10 && ~x2 && ~x4 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s165;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && x12 && ~x10 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && x12 && ~x10 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && x12 && ~x10 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && x12 && ~x10 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && ~x12 && x9 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && ~x12 && x9 && ~x2 && x4 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && ~x12 && x9 && ~x2 && ~x4 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s165;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && ~x12 && ~x9 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && ~x12 && ~x9 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && ~x12 && ~x9 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && x17 && ~x13 && ~x11 && ~x12 && ~x9 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && ~x17 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && ~x17 && ~x2 && x4 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && x26 && ~x17 && ~x2 && ~x4 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && x11 && x9 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && x11 && x9 && ~x4 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && x11 && ~x9 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && x11 && ~x9 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && x11 && ~x9 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && x11 && ~x9 && ~x20 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && ~x11 && x12 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && ~x11 && x12 && ~x4 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && ~x11 && ~x12 && x7 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && ~x11 && ~x12 && x7 && ~x4 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && ~x11 && ~x12 && ~x7 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && ~x11 && ~x12 && ~x7 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && ~x11 && ~x12 && ~x7 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && x13 && ~x11 && ~x12 && ~x7 && ~x20 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && x11 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s173;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && x11 && ~x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && x12 && x10 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && x12 && x10 && ~x4 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && x12 && ~x10 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && x12 && ~x10 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && x12 && ~x10 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && x12 && ~x10 && ~x20 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && x8 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && x8 && ~x4 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && ~x8 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && ~x8 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && ~x8 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && ~x8 && ~x20 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && ~x17 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x66 && x67 && x24 && ~x16 && ~x26 && ~x3 && ~x17 && ~x4 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s174;
						end
					else if( ~x65 && ~x66 && x67 && ~x24 && x25 && x26 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x66 && x67 && ~x24 && x25 && ~x26 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && x67 && ~x24 && x25 && ~x26 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && x67 && ~x24 && x25 && ~x26 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && ~x24 && x25 && ~x26 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && ~x24 && ~x25 && x26 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x65 && ~x66 && x67 && ~x24 && ~x25 && x26 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x65 && ~x66 && x67 && ~x24 && ~x25 && x26 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && ~x24 && ~x25 && ~x26 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && x68 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && x21 && x10 && x11 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && x21 && x10 && ~x11 )
						nx_state = s23;
					else if( ~x65 && ~x66 && ~x67 && ~x68 && x21 && ~x10 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s104;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s176;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && x19 && x15 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y17 = 1'b1;	
							nx_state = s177;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && x19 && ~x15 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && x15 && x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && x15 && ~x14 && x16 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && x15 && ~x14 && ~x16 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && x15 && ~x14 && ~x16 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && x15 && ~x14 && ~x16 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && x15 && ~x14 && ~x16 && ~x5 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && ~x15 && x14 && x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && ~x15 && x14 && ~x18 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && ~x15 && x14 && ~x18 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && ~x15 && x14 && ~x18 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && ~x15 && x14 && ~x18 && ~x5 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && ~x15 && ~x14 && x17 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && ~x5 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && x10 && ~x19 && ~x20 )
						begin
							y21 = 1'b1;	
							nx_state = s151;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x22 && ~x8 && ~x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x22 && x10 && x19 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x22 && x10 && x19 && ~x15 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x22 && x10 && ~x19 && x20 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x22 && x10 && ~x19 && ~x20 )
						begin
							y21 = 1'b1;	
							nx_state = s151;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x22 && ~x10 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s104;
						end
					else nx_state = s23;
				s24 : if( x65 && x21 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x21 && x22 && x23 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( x65 && ~x21 && x22 && ~x23 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x65 && ~x21 && ~x22 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x66 && x67 && x64 && x63 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && x66 && x67 && x64 && ~x63 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x64 && x63 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x66 && x67 && ~x64 && ~x63 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( ~x65 && x66 && ~x67 && x21 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s180;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x24 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && x10 && x26 && x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && x10 && x26 && ~x12 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && x10 && ~x26 && x12 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s165;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && x10 && ~x26 && ~x12 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && x11 && x26 && x12 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s165;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && x11 && x26 && ~x12 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && x11 && ~x26 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && x11 && ~x26 && ~x12 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && x12 && x13 && x26 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && x12 && x13 && ~x26 )
						begin
							y8 = 1'b1;	
							nx_state = s181;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && x12 && ~x13 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && x12 && ~x13 && x19 && ~x14 && x26 )
						nx_state = s24;
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && x12 && ~x13 && x19 && ~x14 && ~x26 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && x12 && ~x13 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && ~x12 && x14 && x26 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && ~x12 && x14 && ~x26 )
						begin
							y8 = 1'b1;	
							nx_state = s181;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && ~x12 && ~x14 && x19 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && ~x12 && ~x14 && x19 && ~x13 && x26 )
						nx_state = s24;
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && ~x12 && ~x14 && x19 && ~x13 && ~x26 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && x16 && ~x10 && ~x11 && ~x12 && ~x14 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && x10 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && x10 && ~x3 && x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && x10 && ~x3 && ~x1 && x11 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s171;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && x10 && ~x3 && ~x1 && ~x11 && x12 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s183;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && x10 && ~x3 && ~x1 && ~x11 && ~x12 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && ~x10 && x11 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && ~x10 && x11 && ~x12 )
						begin
							y6 = 1'b1;	
							nx_state = s172;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && ~x10 && ~x11 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && ~x10 && ~x11 && ~x3 && x12 && x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && ~x10 && ~x11 && ~x3 && x12 && ~x1 )
						begin
							y6 = 1'b1;	
							nx_state = s184;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && ~x10 && ~x11 && ~x3 && ~x12 && x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && x26 && ~x10 && ~x11 && ~x3 && ~x12 && ~x1 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && x10 && x5 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && x10 && ~x5 && x2 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s174;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && x10 && ~x5 && ~x2 && x11 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s187;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && x10 && ~x5 && ~x2 && ~x11 && x12 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s187;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && x10 && ~x5 && ~x2 && ~x11 && ~x12 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s171;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && ~x10 && x11 && x12 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && ~x10 && x11 && ~x12 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s187;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && ~x10 && ~x11 && x5 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && ~x10 && ~x11 && ~x5 && x2 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s174;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && ~x10 && ~x11 && ~x5 && ~x2 && x12 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s187;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x15 && ~x16 && ~x26 && ~x10 && ~x11 && ~x5 && ~x2 && ~x12 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && x10 && x12 && x8 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && x10 && x12 && ~x8 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && x10 && x12 && ~x8 && ~x3 && x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && x10 && x12 && ~x8 && ~x3 && ~x1 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && x10 && ~x12 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && x12 && x7 && x11 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && x12 && x7 && x11 && ~x3 && x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && x12 && x7 && x11 && ~x3 && ~x1 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && x12 && x7 && ~x11 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && x12 && ~x7 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && x12 && ~x7 && ~x3 && x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && x12 && ~x7 && ~x3 && ~x1 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && ~x12 && x11 && x9 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && ~x12 && x11 && ~x9 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && ~x12 && x11 && ~x9 && ~x3 && x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && ~x12 && x11 && ~x9 && ~x3 && ~x1 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && ~x12 && ~x11 && x8 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && ~x12 && ~x11 && x8 && ~x3 && x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && ~x12 && ~x11 && x8 && ~x3 && ~x1 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && x16 && ~x10 && ~x12 && ~x11 && ~x8 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && ~x16 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && ~x16 && ~x3 && x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && x26 && ~x16 && ~x3 && ~x1 )
						begin
							y6 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && x5 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && x10 && x8 && x2 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s174;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && x10 && x8 && ~x2 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && x10 && ~x8 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && x10 && ~x8 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && x10 && ~x8 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && x10 && ~x8 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && ~x10 && x11 && x2 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s174;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && ~x10 && x11 && ~x2 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && ~x10 && ~x11 && x7 && x2 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s174;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && ~x10 && ~x11 && x7 && ~x2 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && ~x10 && ~x11 && ~x7 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && ~x10 && ~x11 && ~x7 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && ~x10 && ~x11 && ~x7 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && x12 && ~x10 && ~x11 && ~x7 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && x10 && x2 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && x10 && ~x2 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s174;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && x11 && x9 && x2 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s174;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && x11 && x9 && ~x2 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && x11 && ~x9 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && x11 && ~x9 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && x11 && ~x9 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && x11 && ~x9 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && ~x11 && x8 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && ~x11 && x8 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && ~x11 && x8 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && ~x11 && x8 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && ~x11 && ~x8 && x2 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s174;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && x16 && ~x12 && ~x10 && ~x11 && ~x8 && ~x2 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && ~x16 && x2 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s174;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x15 && ~x26 && ~x5 && ~x16 && ~x2 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s19;
						end
					else if( ~x65 && ~x66 && ~x24 && ~x25 && x26 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x65 && ~x66 && ~x24 && ~x25 && ~x26 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s190;
						end
					else nx_state = s24;
				s25 : if( x66 && x65 && x15 && x16 && x12 && x10 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x66 && x65 && x15 && x16 && x12 && ~x10 && x20 && x13 && x11 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s126;
						end
					else if( x66 && x65 && x15 && x16 && x12 && ~x10 && x20 && x13 && ~x11 )
						begin
							y4 = 1'b1;	
							nx_state = s191;
						end
					else if( x66 && x65 && x15 && x16 && x12 && ~x10 && x20 && ~x13 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && x65 && x15 && x16 && x12 && ~x10 && x20 && ~x13 && x19 && ~x14 )
						nx_state = s1;
					else if( x66 && x65 && x15 && x16 && x12 && ~x10 && x20 && ~x13 && ~x19 )
						nx_state = s1;
					else if( x66 && x65 && x15 && x16 && x12 && ~x10 && ~x20 && x21 && x11 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s126;
						end
					else if( x66 && x65 && x15 && x16 && x12 && ~x10 && ~x20 && x21 && ~x11 && x13 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s125;
						end
					else if( x66 && x65 && x15 && x16 && x12 && ~x10 && ~x20 && x21 && ~x11 && ~x13 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && x15 && x16 && x12 && ~x10 && ~x20 && x21 && ~x11 && ~x13 && x19 && ~x14 )
						nx_state = s1;
					else if( x66 && x65 && x15 && x16 && x12 && ~x10 && ~x20 && x21 && ~x11 && ~x13 && ~x19 )
						nx_state = s1;
					else if( x66 && x65 && x15 && x16 && x12 && ~x10 && ~x20 && ~x21 && x13 && x11 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s126;
						end
					else if( x66 && x65 && x15 && x16 && x12 && ~x10 && ~x20 && ~x21 && x13 && ~x11 )
						begin
							y4 = 1'b1;	
							nx_state = s191;
						end
					else if( x66 && x65 && x15 && x16 && x12 && ~x10 && ~x20 && ~x21 && ~x13 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && x65 && x15 && x16 && x12 && ~x10 && ~x20 && ~x21 && ~x13 && x19 && ~x14 )
						nx_state = s1;
					else if( x66 && x65 && x15 && x16 && x12 && ~x10 && ~x20 && ~x21 && ~x13 && ~x19 )
						nx_state = s1;
					else if( x66 && x65 && x15 && x16 && ~x12 && x10 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( x66 && x65 && x15 && x16 && ~x12 && ~x10 && x11 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s192;
						end
					else if( x66 && x65 && x15 && x16 && ~x12 && ~x10 && ~x11 && x14 && x20 )
						begin
							y4 = 1'b1;	
							nx_state = s191;
						end
					else if( x66 && x65 && x15 && x16 && ~x12 && ~x10 && ~x11 && x14 && ~x20 && x21 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s125;
						end
					else if( x66 && x65 && x15 && x16 && ~x12 && ~x10 && ~x11 && x14 && ~x20 && ~x21 )
						begin
							y4 = 1'b1;	
							nx_state = s191;
						end
					else if( x66 && x65 && x15 && x16 && ~x12 && ~x10 && ~x11 && ~x14 && x19 && x13 && x20 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && x65 && x15 && x16 && ~x12 && ~x10 && ~x11 && ~x14 && x19 && x13 && ~x20 && x21 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && x15 && x16 && ~x12 && ~x10 && ~x11 && ~x14 && x19 && x13 && ~x20 && ~x21 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && x65 && x15 && x16 && ~x12 && ~x10 && ~x11 && ~x14 && x19 && ~x13 )
						nx_state = s1;
					else if( x66 && x65 && x15 && x16 && ~x12 && ~x10 && ~x11 && ~x14 && ~x19 )
						nx_state = s1;
					else if( x66 && x65 && x15 && ~x16 && x10 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x66 && x65 && x15 && ~x16 && x10 && ~x2 && x20 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x66 && x65 && x15 && ~x16 && x10 && ~x2 && x20 && ~x4 && x11 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x66 && x65 && x15 && ~x16 && x10 && ~x2 && x20 && ~x4 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s193;
						end
					else if( x66 && x65 && x15 && ~x16 && x10 && ~x2 && x20 && ~x4 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s194;
						end
					else if( x66 && x65 && x15 && ~x16 && x10 && ~x2 && ~x20 && x21 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( x66 && x65 && x15 && ~x16 && x10 && ~x2 && ~x20 && x21 && ~x3 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x66 && x65 && x15 && ~x16 && x10 && ~x2 && ~x20 && x21 && ~x3 && ~x11 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s193;
						end
					else if( x66 && x65 && x15 && ~x16 && x10 && ~x2 && ~x20 && x21 && ~x3 && ~x11 && ~x12 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s195;
						end
					else if( x66 && x65 && x15 && ~x16 && x10 && ~x2 && ~x20 && ~x21 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x66 && x65 && x15 && ~x16 && x10 && ~x2 && ~x20 && ~x21 && ~x4 && x11 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x66 && x65 && x15 && ~x16 && x10 && ~x2 && ~x20 && ~x21 && ~x4 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s193;
						end
					else if( x66 && x65 && x15 && ~x16 && x10 && ~x2 && ~x20 && ~x21 && ~x4 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s194;
						end
					else if( x66 && x65 && x15 && ~x16 && ~x10 && x11 && x20 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x66 && x65 && x15 && ~x16 && ~x10 && x11 && ~x20 && x21 && x12 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && x65 && x15 && ~x16 && ~x10 && x11 && ~x20 && x21 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s194;
						end
					else if( x66 && x65 && x15 && ~x16 && ~x10 && x11 && ~x20 && ~x21 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x66 && x65 && x15 && ~x16 && ~x10 && ~x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x66 && x65 && x15 && ~x16 && ~x10 && ~x11 && ~x2 && x20 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x66 && x65 && x15 && ~x16 && ~x10 && ~x11 && ~x2 && x20 && ~x4 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s196;
						end
					else if( x66 && x65 && x15 && ~x16 && ~x10 && ~x11 && ~x2 && x20 && ~x4 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s192;
						end
					else if( x66 && x65 && x15 && ~x16 && ~x10 && ~x11 && ~x2 && ~x20 && x21 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( x66 && x65 && x15 && ~x16 && ~x10 && ~x11 && ~x2 && ~x20 && x21 && ~x3 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( x66 && x65 && x15 && ~x16 && ~x10 && ~x11 && ~x2 && ~x20 && x21 && ~x3 && ~x12 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s198;
						end
					else if( x66 && x65 && x15 && ~x16 && ~x10 && ~x11 && ~x2 && ~x20 && ~x21 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x66 && x65 && x15 && ~x16 && ~x10 && ~x11 && ~x2 && ~x20 && ~x21 && ~x4 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s196;
						end
					else if( x66 && x65 && x15 && ~x16 && ~x10 && ~x11 && ~x2 && ~x20 && ~x21 && ~x4 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s192;
						end
					else if( x66 && x65 && ~x15 && x20 && x16 && x10 && x12 && x8 )
						nx_state = s1;
					else if( x66 && x65 && ~x15 && x20 && x16 && x10 && x12 && ~x8 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x66 && x65 && ~x15 && x20 && x16 && x10 && x12 && ~x8 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x66 && x65 && ~x15 && x20 && x16 && x10 && x12 && ~x8 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s199;
						end
					else if( x66 && x65 && ~x15 && x20 && x16 && x10 && ~x12 && x9 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x66 && x65 && ~x15 && x20 && x16 && x10 && ~x12 && x9 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s200;
						end
					else if( x66 && x65 && ~x15 && x20 && x16 && x10 && ~x12 && x9 && ~x2 && ~x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x66 && x65 && ~x15 && x20 && x16 && x10 && ~x12 && ~x9 )
						nx_state = s1;
					else if( x66 && x65 && ~x15 && x20 && x16 && ~x10 && x12 && x7 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x66 && x65 && ~x15 && x20 && x16 && ~x10 && x12 && x7 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x66 && x65 && ~x15 && x20 && x16 && ~x10 && x12 && x7 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s199;
						end
					else if( x66 && x65 && ~x15 && x20 && x16 && ~x10 && x12 && ~x7 && x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x66 && x65 && ~x15 && x20 && x16 && ~x10 && x12 && ~x7 && x11 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x66 && x65 && ~x15 && x20 && x16 && ~x10 && x12 && ~x7 && x11 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s199;
						end
					else if( x66 && x65 && ~x15 && x20 && x16 && ~x10 && x12 && ~x7 && ~x11 )
						nx_state = s1;
					else if( x66 && x65 && ~x15 && x20 && x16 && ~x10 && ~x12 && x11 && x9 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x66 && x65 && ~x15 && x20 && x16 && ~x10 && ~x12 && x11 && x9 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x66 && x65 && ~x15 && x20 && x16 && ~x10 && ~x12 && x11 && x9 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s199;
						end
					else if( x66 && x65 && ~x15 && x20 && x16 && ~x10 && ~x12 && x11 && ~x9 )
						nx_state = s1;
					else if( x66 && x65 && ~x15 && x20 && x16 && ~x10 && ~x12 && ~x11 && x8 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x66 && x65 && ~x15 && x20 && x16 && ~x10 && ~x12 && ~x11 && x8 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x66 && x65 && ~x15 && x20 && x16 && ~x10 && ~x12 && ~x11 && x8 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s199;
						end
					else if( x66 && x65 && ~x15 && x20 && x16 && ~x10 && ~x12 && ~x11 && ~x8 )
						nx_state = s1;
					else if( x66 && x65 && ~x15 && x20 && ~x16 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x66 && x65 && ~x15 && x20 && ~x16 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x66 && x65 && ~x15 && x20 && ~x16 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s201;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && x10 && x8 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s202;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && x10 && x8 && ~x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && x10 && ~x8 && x12 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && x10 && ~x8 && x12 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && x10 && ~x8 && x12 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && x10 && ~x8 && x12 && ~x19 )
						nx_state = s1;
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && x10 && ~x8 && ~x12 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s202;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && x10 && ~x8 && ~x12 && ~x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && x12 && x11 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && x12 && x11 && ~x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y11 = 1'b1;	
							nx_state = s192;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && x12 && ~x11 && x7 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s202;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && x12 && ~x11 && x7 && ~x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && x12 && ~x11 && ~x7 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && x12 && ~x11 && ~x7 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && x12 && ~x11 && ~x7 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && x12 && ~x11 && ~x7 && ~x19 )
						nx_state = s1;
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && x11 && x9 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s202;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && x11 && x9 && ~x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && x11 && ~x9 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && x11 && ~x9 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && x11 && ~x9 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && x11 && ~x9 && ~x19 )
						nx_state = s1;
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && ~x11 && x8 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && ~x11 && x8 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && ~x11 && x8 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && ~x11 && x8 && ~x19 )
						nx_state = s1;
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && ~x11 && ~x8 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s202;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && x16 && ~x10 && ~x12 && ~x11 && ~x8 && ~x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && ~x16 && x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( x66 && x65 && ~x15 && ~x20 && x21 && ~x2 && ~x16 && ~x3 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && x10 && x12 && x8 )
						nx_state = s1;
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && x10 && x12 && ~x8 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && x10 && x12 && ~x8 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && x10 && x12 && ~x8 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s199;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && x10 && ~x12 && x9 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && x10 && ~x12 && x9 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s200;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && x10 && ~x12 && x9 && ~x2 && ~x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && x10 && ~x12 && ~x9 )
						nx_state = s1;
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && x12 && x7 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && x12 && x7 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && x12 && x7 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s199;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && x12 && ~x7 && x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && x12 && ~x7 && x11 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && x12 && ~x7 && x11 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s199;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && x12 && ~x7 && ~x11 )
						nx_state = s1;
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && ~x12 && x11 && x9 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && ~x12 && x11 && x9 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && ~x12 && x11 && x9 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s199;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && ~x12 && x11 && ~x9 )
						nx_state = s1;
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && ~x12 && ~x11 && x8 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && ~x12 && ~x11 && x8 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && ~x12 && ~x11 && x8 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s199;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && x16 && ~x10 && ~x12 && ~x11 && ~x8 )
						nx_state = s1;
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && ~x16 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && ~x16 && ~x2 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x66 && x65 && ~x15 && ~x20 && ~x21 && ~x16 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s201;
						end
					else if( x66 && ~x65 && x62 && x16 && x15 && x14 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && ~x65 && x62 && x16 && x15 && x14 && ~x9 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && ~x65 && x62 && x16 && x15 && ~x14 && x7 && x9 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s157;
						end
					else if( x66 && ~x65 && x62 && x16 && x15 && ~x14 && x7 && ~x9 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s158;
						end
					else if( x66 && ~x65 && x62 && x16 && x15 && ~x14 && ~x7 && x9 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s65;
						end
					else if( x66 && ~x65 && x62 && x16 && x15 && ~x14 && ~x7 && x9 && ~x12 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x66 && ~x65 && x62 && x16 && x15 && ~x14 && ~x7 && x9 && ~x12 && x61 && ~x13 )
						nx_state = s1;
					else if( x66 && ~x65 && x62 && x16 && x15 && ~x14 && ~x7 && x9 && ~x12 && ~x61 )
						nx_state = s1;
					else if( x66 && ~x65 && x62 && x16 && x15 && ~x14 && ~x7 && ~x9 && x13 )
						begin
							y3 = 1'b1;	
							nx_state = s65;
						end
					else if( x66 && ~x65 && x62 && x16 && x15 && ~x14 && ~x7 && ~x9 && ~x13 && x61 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x66 && ~x65 && x62 && x16 && x15 && ~x14 && ~x7 && ~x9 && ~x13 && x61 && ~x12 )
						nx_state = s1;
					else if( x66 && ~x65 && x62 && x16 && x15 && ~x14 && ~x7 && ~x9 && ~x13 && ~x61 )
						nx_state = s1;
					else if( x66 && ~x65 && x62 && x16 && ~x15 && x9 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( x66 && ~x65 && x62 && x16 && ~x15 && x9 && ~x3 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x66 && ~x65 && x62 && x16 && ~x15 && x9 && ~x3 && ~x4 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && x7 && x11 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && x7 && x11 && ~x3 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && x7 && x11 && ~x3 && ~x4 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && x7 && ~x11 && x3 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && x7 && ~x11 && ~x3 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && x7 && ~x11 && ~x3 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && x7 && ~x11 && ~x3 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && x7 && ~x11 && ~x3 && ~x61 )
						nx_state = s1;
					else if( x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && ~x7 && x10 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && ~x7 && x10 && ~x3 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && ~x7 && x10 && ~x3 && ~x4 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && ~x7 && ~x10 && x3 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && ~x7 && ~x10 && ~x3 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && ~x7 && ~x10 && ~x3 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && ~x7 && ~x10 && ~x3 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x66 && ~x65 && x62 && x16 && ~x15 && ~x9 && ~x7 && ~x10 && ~x3 && ~x61 )
						nx_state = s1;
					else if( x66 && ~x65 && x62 && ~x16 && x15 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( x66 && ~x65 && x62 && ~x16 && x15 && ~x7 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( x66 && ~x65 && x62 && ~x16 && x15 && ~x7 && ~x3 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x66 && ~x65 && x62 && ~x16 && x15 && ~x7 && ~x3 && ~x4 && x8 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x66 && ~x65 && x62 && ~x16 && x15 && ~x7 && ~x3 && ~x4 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( x66 && ~x65 && x62 && ~x16 && ~x15 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( x66 && ~x65 && x62 && ~x16 && ~x15 && ~x3 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x66 && ~x65 && x62 && ~x16 && ~x15 && ~x3 && ~x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( x66 && ~x65 && ~x62 && x63 && x64 && x17 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && ~x65 && ~x62 && x63 && x64 && x17 && ~x13 && x12 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && ~x65 && ~x62 && x63 && x64 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x62 && x63 && x64 && ~x17 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x62 && x63 && ~x64 && x15 && x8 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x66 && ~x65 && ~x62 && x63 && ~x64 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x66 && ~x65 && ~x62 && x63 && ~x64 && ~x15 && x16 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x66 && ~x65 && ~x62 && x63 && ~x64 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s135;
						end
					else if( x66 && ~x65 && ~x62 && ~x63 && x64 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x66 && ~x65 && ~x62 && ~x63 && ~x64 && x6 && x15 && x8 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && ~x65 && ~x62 && ~x63 && ~x64 && x6 && x15 && ~x8 )
						begin
							y18 = 1'b1;	
							nx_state = s203;
						end
					else if( x66 && ~x65 && ~x62 && ~x63 && ~x64 && x6 && ~x15 && x16 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && ~x65 && ~x62 && ~x63 && ~x64 && x6 && ~x15 && ~x16 && x14 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s204;
						end
					else if( x66 && ~x65 && ~x62 && ~x63 && ~x64 && x6 && ~x15 && ~x16 && ~x14 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s20;
						end
					else if( x66 && ~x65 && ~x62 && ~x63 && ~x64 && ~x6 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x66 && x65 && x21 && x15 && x9 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x66 && x65 && x21 && x15 && ~x9 && x6 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x66 && x65 && x21 && x15 && ~x9 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x66 && x65 && x21 && ~x15 && x16 && x9 && x8 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x66 && x65 && x21 && ~x15 && x16 && x9 && ~x8 && x10 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x66 && x65 && x21 && ~x15 && x16 && x9 && ~x8 && ~x10 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x66 && x65 && x21 && ~x15 && x16 && x9 && ~x8 && ~x10 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && x21 && ~x15 && x16 && x9 && ~x8 && ~x10 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && x21 && ~x15 && x16 && x9 && ~x8 && ~x10 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && x21 && ~x15 && x16 && x9 && ~x8 && ~x10 && ~x18 && ~x19 )
						nx_state = s1;
					else if( ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && x8 && x12 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && x8 && ~x12 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && x8 && ~x12 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && x8 && ~x12 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && x8 && ~x12 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && x8 && ~x12 && ~x18 && ~x19 )
						nx_state = s1;
					else if( ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && ~x8 && x11 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && ~x8 && ~x11 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && ~x8 && ~x11 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && ~x8 && ~x11 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && ~x8 && ~x11 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && x21 && ~x15 && x16 && ~x9 && ~x8 && ~x11 && ~x18 && ~x19 )
						nx_state = s1;
					else if( ~x66 && x65 && x21 && ~x15 && ~x16 && x6 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x66 && x65 && x21 && ~x15 && ~x16 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x66 && x65 && ~x21 && x22 && x18 && x14 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( ~x66 && x65 && ~x21 && x22 && x18 && ~x14 && x13 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( ~x66 && x65 && ~x21 && x22 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && x22 && ~x18 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && x23 && x15 && x9 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && x23 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && x23 && ~x15 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x23 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && ~x65 && x68 && x20 && x15 && x8 )
						begin
							y2 = 1'b1;	y13 = 1'b1;	
							nx_state = s206;
						end
					else if( ~x66 && ~x65 && x68 && x20 && x15 && ~x8 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x66 && ~x65 && x68 && x20 && x15 && ~x8 && ~x6 )
						begin
							y2 = 1'b1;	y13 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x66 && ~x65 && x68 && x20 && ~x15 && x16 && x7 && x8 )
						begin
							y2 = 1'b1;	y13 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x66 && ~x65 && x68 && x20 && ~x15 && x16 && x7 && ~x8 )
						begin
							y2 = 1'b1;	y13 = 1'b1;	
							nx_state = s206;
						end
					else if( ~x66 && ~x65 && x68 && x20 && ~x15 && x16 && ~x7 )
						begin
							y2 = 1'b1;	y13 = 1'b1;	
							nx_state = s206;
						end
					else if( ~x66 && ~x65 && x68 && x20 && ~x15 && ~x16 && x6 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s209;
						end
					else if( ~x66 && ~x65 && x68 && x20 && ~x15 && ~x16 && ~x6 )
						begin
							y2 = 1'b1;	y13 = 1'b1;	
							nx_state = s208;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && x21 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && x14 && x8 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && x14 && ~x8 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s126;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && ~x14 && x7 && x8 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	y20 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && ~x14 && x7 && ~x8 )
						begin
							y12 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && ~x14 && ~x7 && x8 && x12 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && x17 && ~x13 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && ~x17 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && ~x14 && ~x7 && ~x8 && x13 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && x17 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && x17 && ~x12 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && ~x17 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && x7 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && x7 && ~x2 && x3 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && x7 && ~x2 && ~x3 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && ~x7 && x9 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && ~x7 && x9 && ~x2 && x3 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && ~x7 && x9 && ~x2 && ~x3 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && ~x7 && ~x9 && x2 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && ~x7 && ~x9 && ~x2 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && ~x7 && ~x9 && ~x2 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && ~x7 && ~x9 && ~x2 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && x8 && ~x7 && ~x9 && ~x2 && ~x17 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && x7 && x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && x7 && x11 && ~x2 && x3 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && x7 && x11 && ~x2 && ~x3 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && x7 && ~x11 && x2 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && x7 && ~x11 && ~x2 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && x7 && ~x11 && ~x2 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && x7 && ~x11 && ~x2 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && x7 && ~x11 && ~x2 && ~x17 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && ~x7 && x10 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && ~x7 && x10 && ~x2 && x3 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && ~x7 && x10 && ~x2 && ~x3 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && x2 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x2 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x2 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x2 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x2 && ~x17 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x16 && x15 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x16 && x15 && ~x7 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x16 && x15 && ~x7 && ~x2 && x3 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x16 && x15 && ~x7 && ~x2 && ~x3 && x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x16 && x15 && ~x7 && ~x2 && ~x3 && ~x8 )
						begin
							y2 = 1'b1;	y13 = 1'b1;	
							nx_state = s206;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x16 && ~x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x16 && ~x15 && ~x2 && x3 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x66 && ~x65 && x68 && ~x20 && ~x21 && ~x16 && ~x15 && ~x2 && ~x3 )
						begin
							y7 = 1'b1;	y12 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x66 && ~x65 && ~x68 && x24 && x26 && x11 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x66 && ~x65 && ~x68 && x24 && x26 && ~x11 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x66 && ~x65 && ~x68 && x24 && x26 && ~x11 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x66 && ~x65 && ~x68 && x24 && x26 && ~x11 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x68 && x24 && x26 && ~x11 && ~x18 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x68 && x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x66 && ~x65 && ~x68 && x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x66 && ~x65 && ~x68 && x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x68 && x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x68 && ~x24 && x25 && x26 && x15 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x68 && ~x24 && x25 && x26 && ~x15 && x3 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x66 && ~x65 && ~x68 && ~x24 && x25 && x26 && ~x15 && ~x3 && x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x66 && ~x65 && ~x68 && ~x24 && x25 && x26 && ~x15 && ~x3 && ~x1 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x18 && x15 && x10 && x11 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s187;
						end
					else if( ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x18 && x15 && x10 && ~x11 && x12 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x18 && x15 && x10 && ~x11 && ~x12 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x18 && x15 && ~x10 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x18 && ~x15 && x16 && x10 && x12 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x18 && ~x15 && x16 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x18 && ~x15 && x16 && ~x10 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && x18 && ~x15 && ~x16 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x66 && ~x65 && ~x68 && ~x24 && x25 && ~x26 && ~x18 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && x10 && x12 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && x10 && x12 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && x10 && x12 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && x10 && x12 && ~x18 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && x10 && ~x12 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s165;
						end
					else if( ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && ~x10 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && ~x10 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && ~x10 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && x26 && ~x10 && ~x18 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x68 && ~x24 && ~x25 && ~x26 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else nx_state = s25;
				s26 : if( x65 && x21 && x15 && x9 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( x65 && x21 && x15 && ~x9 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( x65 && x21 && ~x15 && x16 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x65 && x21 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s212;
						end
					else if( x65 && ~x21 && x23 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x23 && x22 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x21 && ~x23 && ~x22 && x17 && x15 && x9 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( x65 && ~x21 && ~x23 && ~x22 && x17 && x15 && ~x9 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( x65 && ~x21 && ~x23 && ~x22 && x17 && ~x15 && x16 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( x65 && ~x21 && ~x23 && ~x22 && x17 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s205;
						end
					else if( x65 && ~x21 && ~x23 && ~x22 && ~x17 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( ~x65 && x62 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( ~x65 && ~x62 && x63 )
						begin
							y19 = 1'b1;	
							nx_state = s213;
						end
					else if( ~x65 && ~x62 && ~x63 )
						nx_state = s1;
					else nx_state = s26;
				s27 : if( x66 && x65 && x67 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && x65 && x67 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && x65 && x67 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x66 && x65 && x67 && x22 && ~x17 )
						nx_state = s1;
					else if( x66 && x65 && x67 && ~x22 && x18 && x13 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x66 && x65 && x67 && ~x22 && x18 && x13 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && x67 && ~x22 && x18 && ~x13 && x12 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x66 && x65 && x67 && ~x22 && x18 && ~x13 && x12 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && x67 && ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x66 && x65 && x67 && ~x22 && ~x18 )
						nx_state = s1;
					else if( x66 && x65 && ~x67 && x21 && x20 && x12 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && x65 && ~x67 && x21 && x20 && x12 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && x65 && ~x67 && x21 && x20 && x12 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && x65 && ~x67 && x21 && x20 && x12 && ~x17 )
						nx_state = s1;
					else if( x66 && x65 && ~x67 && x21 && x20 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( x66 && x65 && ~x67 && x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && ~x67 && x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && ~x67 && x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( x66 && x65 && ~x67 && ~x21 && x12 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && x65 && ~x67 && ~x21 && x12 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && x65 && ~x67 && ~x21 && x12 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && x65 && ~x67 && ~x21 && x12 && ~x19 )
						nx_state = s1;
					else if( x66 && x65 && ~x67 && ~x21 && ~x12 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x66 && ~x65 && x67 && x62 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x66 && ~x65 && x67 && x62 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x66 && ~x65 && x67 && x62 && ~x15 && x16 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x66 && ~x65 && x67 && x62 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y28 = 1'b1;	
							nx_state = s135;
						end
					else if( x66 && ~x65 && x67 && ~x62 && x63 && x6 && x15 && x8 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && ~x65 && x67 && ~x62 && x63 && x6 && x15 && ~x8 )
						begin
							y18 = 1'b1;	
							nx_state = s203;
						end
					else if( x66 && ~x65 && x67 && ~x62 && x63 && x6 && ~x15 && x16 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && ~x65 && x67 && ~x62 && x63 && x6 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s204;
						end
					else if( x66 && ~x65 && x67 && ~x62 && x63 && ~x6 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && ~x65 && x67 && ~x62 && ~x63 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && x21 && x16 && x15 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s214;
						end
					else if( x66 && ~x65 && ~x67 && x21 && x16 && x15 && ~x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s215;
						end
					else if( x66 && ~x65 && ~x67 && x21 && x16 && ~x15 && x10 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x66 && ~x65 && ~x67 && x21 && x16 && ~x15 && ~x10 )
						begin
							y14 = 1'b1;	y16 = 1'b1;	
							nx_state = s216;
						end
					else if( x66 && ~x65 && ~x67 && x21 && ~x16 && x17 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s215;
						end
					else if( x66 && ~x65 && ~x67 && x21 && ~x16 && x17 && ~x10 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	
							nx_state = s217;
						end
					else if( x66 && ~x65 && ~x67 && x21 && ~x16 && ~x17 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s215;
						end
					else if( x66 && ~x65 && ~x67 && x21 && ~x16 && ~x17 && ~x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s218;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && x10 && x22 && x4 && x17 && x15 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s219;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && x10 && x22 && x4 && x17 && ~x15 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && x10 && x22 && x4 && ~x17 && x18 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s219;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && x10 && x22 && x4 && ~x17 && ~x18 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s219;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && x10 && x22 && ~x4 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && x10 && ~x22 && x7 && x16 && x15 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s219;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && x10 && ~x22 && x7 && x16 && ~x15 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s220;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && x10 && ~x22 && x7 && ~x16 && x17 && x15 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s219;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && x10 && ~x22 && x7 && ~x16 && x17 && ~x15 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s220;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && x10 && ~x22 && x7 && ~x16 && ~x17 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s219;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && x10 && ~x22 && ~x7 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s220;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && x17 && x4 && x15 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s219;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && x17 && x4 && ~x15 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	
							nx_state = s221;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && x17 && ~x4 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && x15 && x12 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && x15 && ~x12 && x14 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && x15 && ~x12 && ~x14 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && x15 && ~x12 && ~x14 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && x15 && ~x12 && ~x14 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && x15 && ~x12 && ~x14 && ~x7 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && ~x15 && x14 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && ~x15 && x14 && ~x13 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && ~x15 && x14 && ~x13 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && ~x15 && x14 && ~x13 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && ~x15 && x14 && ~x13 && ~x7 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && ~x15 && ~x14 && x11 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && ~x15 && ~x14 && ~x11 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && ~x15 && ~x14 && ~x11 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && ~x15 && ~x14 && ~x11 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && x18 && ~x15 && ~x14 && ~x11 && ~x7 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && ~x18 && x4 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s220;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && x22 && ~x17 && ~x18 && ~x4 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && x16 && x7 && x15 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s222;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && x16 && x7 && ~x15 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && x16 && ~x7 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s220;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && x14 && x13 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s220;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && x14 && ~x13 && x15 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s220;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && x14 && ~x13 && ~x15 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && x14 && ~x13 && ~x15 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && x14 && ~x13 && ~x15 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && x14 && ~x13 && ~x15 && ~x4 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && ~x14 && x15 && x12 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s220;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && ~x14 && x15 && ~x12 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && ~x14 && x15 && ~x12 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && ~x14 && x15 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && ~x14 && x15 && ~x12 && ~x4 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && ~x14 && ~x15 && x11 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s220;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && ~x14 && ~x15 && ~x11 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && ~x14 && ~x15 && ~x11 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && ~x14 && ~x15 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && x17 && ~x14 && ~x15 && ~x11 && ~x4 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && ~x17 && x7 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x10 && ~x22 && ~x16 && ~x17 && ~x7 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s220;
						end
					else if( ~x66 && x65 && x21 && x67 )
						nx_state = s1;
					else if( ~x66 && x65 && x21 && ~x67 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && x21 && ~x67 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && x21 && ~x67 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && x21 && ~x67 && ~x19 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && x22 && x67 && x23 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x66 && x65 && ~x21 && x22 && x67 && x23 && ~x18 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x66 && x65 && ~x21 && x22 && x67 && x23 && ~x18 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x66 && x65 && ~x21 && x22 && x67 && x23 && ~x18 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && x22 && x67 && x23 && ~x18 && ~x8 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && x22 && x67 && ~x23 )
						begin
							y6 = 1'b1;	y19 = 1'b1;	
							nx_state = s223;
						end
					else if( ~x66 && x65 && ~x21 && x22 && ~x67 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( ~x66 && x65 && ~x21 && x22 && ~x67 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( ~x66 && x65 && ~x21 && x22 && ~x67 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( ~x66 && x65 && ~x21 && x22 && ~x67 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && x22 && ~x67 && ~x19 && ~x17 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && x67 && x23 )
						begin
							y6 = 1'b1;	y19 = 1'b1;	
							nx_state = s223;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && x67 && ~x23 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && x67 && ~x23 && ~x19 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && x67 && ~x23 && ~x19 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && x67 && ~x23 && ~x19 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && x67 && ~x23 && ~x19 && ~x8 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && x7 && x23 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && x7 && x23 && ~x9 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && x7 && ~x23 && x9 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && x7 && ~x23 && ~x9 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && x8 && x23 && x9 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && x8 && x23 && ~x9 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && x8 && ~x23 && x9 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && x8 && ~x23 && ~x9 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && x23 && x13 && x9 )
						begin
							y4 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && x23 && x13 && ~x9 && x14 )
						begin
							y4 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && x23 && x13 && ~x9 && ~x14 && x20 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && x23 && x13 && ~x9 && ~x14 && ~x20 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && x23 && ~x13 && x14 && x9 && x20 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && x23 && ~x13 && x14 && x9 && ~x20 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && x23 && ~x13 && x14 && ~x9 )
						begin
							y4 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && x23 && ~x13 && ~x14 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && ~x23 && x13 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s224;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && ~x23 && x13 && ~x9 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s224;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && ~x23 && x13 && ~x9 && ~x14 && x18 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && ~x23 && x13 && ~x9 && ~x14 && ~x18 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && ~x23 && ~x13 && x14 && x9 && x18 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && ~x23 && ~x13 && x14 && x9 && ~x18 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && ~x23 && ~x13 && x14 && ~x9 )
						begin
							y22 = 1'b1;	
							nx_state = s224;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && x16 && ~x7 && ~x8 && ~x23 && ~x13 && ~x14 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && ~x16 && x7 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && ~x16 && ~x7 && x8 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && ~x16 && ~x7 && ~x8 && x5 )
						begin
							y1 = 1'b1;	
							nx_state = s22;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && ~x16 && ~x7 && ~x8 && ~x5 && x2 && x23 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && ~x16 && ~x7 && ~x8 && ~x5 && x2 && ~x23 && x9 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && ~x16 && ~x7 && ~x8 && ~x5 && x2 && ~x23 && ~x9 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && ~x16 && ~x7 && ~x8 && ~x5 && ~x2 && x9 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && ~x16 && ~x7 && ~x8 && ~x5 && ~x2 && ~x9 && x23 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && x15 && ~x16 && ~x7 && ~x8 && ~x5 && ~x2 && ~x9 && ~x23 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && x5 )
						begin
							y1 = 1'b1;	
							nx_state = s22;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && x9 && x10 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && x9 && ~x10 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && x9 && ~x10 && ~x8 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && x9 && ~x10 && ~x8 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && x9 && ~x10 && ~x8 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && x9 && ~x10 && ~x8 && ~x20 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && ~x9 && x8 && x12 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && ~x9 && x8 && ~x12 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && ~x9 && x8 && ~x12 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && ~x9 && x8 && ~x12 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && ~x9 && x8 && ~x12 && ~x20 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && ~x9 && ~x8 && x11 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && ~x9 && ~x8 && ~x11 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && ~x9 && ~x8 && ~x11 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && ~x9 && ~x8 && ~x11 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && x16 && ~x9 && ~x8 && ~x11 && ~x20 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && ~x16 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && x23 && ~x16 && ~x2 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && x9 && ~x10 && x8 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && x9 && ~x10 && ~x8 && x18 && x14 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && x9 && ~x10 && ~x8 && x18 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && x9 && ~x10 && ~x8 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && x9 && ~x10 && ~x8 && ~x18 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && ~x9 && x8 && x12 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && ~x9 && x8 && ~x12 && x18 && x14 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && ~x9 && x8 && ~x12 && x18 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && ~x9 && x8 && ~x12 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && ~x9 && x8 && ~x12 && ~x18 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && ~x9 && ~x8 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && ~x9 && ~x8 && ~x11 && x18 && x14 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && ~x9 && ~x8 && ~x11 && x18 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && ~x9 && ~x8 && ~x11 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && x16 && ~x9 && ~x8 && ~x11 && ~x18 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && ~x16 && x2 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x66 && x65 && ~x21 && ~x22 && ~x67 && ~x15 && ~x5 && ~x23 && ~x16 && ~x2 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x66 && ~x65 && x67 && x20 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x66 && ~x65 && x67 && ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x66 && ~x65 && x67 && ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x66 && ~x65 && x67 && ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x66 && ~x65 && x67 && ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x67 && x21 && x9 && x3 )
						nx_state = s40;
					else if( ~x66 && ~x65 && ~x67 && x21 && x9 && ~x3 && x4 )
						nx_state = s40;
					else if( ~x66 && ~x65 && ~x67 && x21 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x67 && x21 && ~x9 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && x12 && x19 && x15 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && x12 && x19 && ~x15 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && x12 && ~x19 && x20 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && x12 && ~x19 && ~x20 )
						begin
							y6 = 1'b1;	y21 = 1'b1;	
							nx_state = s225;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s27;
				s28 : if( x21 && x65 )
						nx_state = s1;
					else if( x21 && ~x65 && x16 && x6 && x15 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s214;
						end
					else if( x21 && ~x65 && x16 && x6 && x15 && ~x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s215;
						end
					else if( x21 && ~x65 && x16 && x6 && ~x15 && x10 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x21 && ~x65 && x16 && x6 && ~x15 && ~x10 )
						begin
							y14 = 1'b1;	y16 = 1'b1;	
							nx_state = s216;
						end
					else if( x21 && ~x65 && x16 && ~x6 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s220;
						end
					else if( x21 && ~x65 && ~x16 && x17 && x10 && x6 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s215;
						end
					else if( x21 && ~x65 && ~x16 && x17 && x10 && ~x6 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s220;
						end
					else if( x21 && ~x65 && ~x16 && x17 && ~x10 && x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x21 && ~x65 && ~x16 && x17 && ~x10 && ~x6 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s226;
						end
					else if( x21 && ~x65 && ~x16 && ~x17 && x6 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s215;
						end
					else if( x21 && ~x65 && ~x16 && ~x17 && x6 && ~x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s218;
						end
					else if( x21 && ~x65 && ~x16 && ~x17 && ~x6 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s220;
						end
					else if( ~x21 && x22 && x65 && x23 && x5 && x18 && x15 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && x22 && x65 && x23 && x5 && x18 && ~x15 )
						begin
							y15 = 1'b1;	y20 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x21 && x22 && x65 && x23 && x5 && ~x18 && x19 && x15 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s228;
						end
					else if( ~x21 && x22 && x65 && x23 && x5 && ~x18 && x19 && ~x15 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && x22 && x65 && x23 && x5 && ~x18 && ~x19 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x21 && x22 && x65 && x23 && ~x5 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && x22 && x65 && ~x23 )
						begin
							y12 = 1'b1;	y19 = 1'b1;	
							nx_state = s230;
						end
					else if( ~x21 && x22 && ~x65 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && ~x22 && x65 && x23 && x19 && x6 && x16 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( ~x21 && ~x22 && x65 && x23 && x19 && x6 && ~x16 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x21 && ~x22 && x65 && x23 && x19 && ~x6 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && x20 && x16 && x6 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s228;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && x20 && x16 && ~x6 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && x20 && ~x16 && x17 && x18 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && x20 && ~x16 && x17 && x18 && ~x6 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && x20 && ~x16 && x17 && ~x18 && x14 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && x20 && ~x16 && x17 && ~x18 && ~x14 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && x20 && ~x16 && ~x17 && x18 && x14 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && x20 && ~x16 && ~x17 && x18 && ~x14 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && x20 && ~x16 && ~x17 && ~x18 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && x20 && ~x16 && ~x17 && ~x18 && ~x6 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && ~x20 && x6 )
						begin
							y12 = 1'b1;	
							nx_state = s231;
						end
					else if( ~x21 && ~x22 && x65 && x23 && ~x19 && ~x20 && ~x6 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x65 && ~x23 && x5 && x18 && x15 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x65 && ~x23 && x5 && x18 && ~x15 )
						begin
							y15 = 1'b1;	y20 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x21 && ~x22 && x65 && ~x23 && x5 && ~x18 && x19 && x15 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s228;
						end
					else if( ~x21 && ~x22 && x65 && ~x23 && x5 && ~x18 && x19 && ~x15 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x65 && ~x23 && x5 && ~x18 && ~x19 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x21 && ~x22 && x65 && ~x23 && ~x5 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && ~x65 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s232;
						end
					else nx_state = s28;
				s29 : if( x65 && x21 )
						nx_state = s1;
					else if( x65 && ~x21 && x22 && x23 && x18 && x19 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && ~x21 && x22 && x23 && x18 && x19 && x15 && ~x17 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x21 && x22 && x23 && x18 && x19 && ~x15 && x16 && x17 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s157;
						end
					else if( x65 && ~x21 && x22 && x23 && x18 && x19 && ~x15 && x16 && ~x17 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y20 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s227;
						end
					else if( x65 && ~x21 && x22 && x23 && x18 && x19 && ~x15 && ~x16 && x8 && x10 && x17 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && x22 && x23 && x18 && x19 && ~x15 && ~x16 && x8 && x10 && ~x17 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x65 && ~x21 && x22 && x23 && x18 && x19 && ~x15 && ~x16 && x8 && ~x10 && x11 && x17 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x65 && ~x21 && x22 && x23 && x18 && x19 && ~x15 && ~x16 && x8 && ~x10 && x11 && ~x17 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && x22 && x23 && x18 && x19 && ~x15 && ~x16 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && ~x21 && x22 && x23 && x18 && x19 && ~x15 && ~x16 && ~x8 )
						nx_state = s1;
					else if( x65 && ~x21 && x22 && x23 && x18 && ~x19 && x16 && x15 )
						begin
							y18 = 1'b1;	
							nx_state = s203;
						end
					else if( x65 && ~x21 && x22 && x23 && x18 && ~x19 && x16 && ~x15 && x17 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x65 && ~x21 && x22 && x23 && x18 && ~x19 && x16 && ~x15 && ~x17 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s233;
						end
					else if( x65 && ~x21 && x22 && x23 && x18 && ~x19 && ~x16 && x17 && x15 )
						begin
							y18 = 1'b1;	
							nx_state = s234;
						end
					else if( x65 && ~x21 && x22 && x23 && x18 && ~x19 && ~x16 && x17 && ~x15 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s235;
						end
					else if( x65 && ~x21 && x22 && x23 && x18 && ~x19 && ~x16 && ~x17 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s236;
						end
					else if( x65 && ~x21 && x22 && x23 && x18 && ~x19 && ~x16 && ~x17 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x65 && ~x21 && x22 && x23 && x18 && ~x19 && ~x16 && ~x17 && ~x4 && ~x6 && x15 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s227;
						end
					else if( x65 && ~x21 && x22 && x23 && x18 && ~x19 && ~x16 && ~x17 && ~x4 && ~x6 && ~x15 )
						begin
							y16 = 1'b1;	y20 = 1'b1;	
							nx_state = s227;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x18 && x19 && x15 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s236;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x18 && x19 && x15 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x18 && x19 && x15 && ~x4 && ~x6 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s117;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && x17 && x13 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s236;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && x17 && x13 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && x17 && x13 && ~x4 && ~x6 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s227;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && x17 && ~x13 && x16 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s236;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && x17 && ~x13 && x16 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && x17 && ~x13 && x16 && ~x4 && ~x6 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s227;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && x17 && ~x13 && ~x16 )
						nx_state = s1;
					else if( x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && ~x17 && x16 && x14 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s236;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && ~x17 && x16 && x14 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && ~x17 && x16 && x14 && ~x4 && ~x6 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s227;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && ~x17 && x16 && ~x14 )
						nx_state = s1;
					else if( x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && x12 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s236;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && x12 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && x12 && ~x4 && ~x6 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s227;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && ~x12 )
						nx_state = s1;
					else if( x65 && ~x21 && x22 && x23 && ~x18 && ~x19 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s236;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x18 && ~x19 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x18 && ~x19 && ~x4 && ~x6 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x65 && ~x21 && x22 && ~x23 && x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( x65 && ~x21 && x22 && ~x23 && ~x15 && x19 && x18 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( x65 && ~x21 && x22 && ~x23 && ~x15 && x19 && ~x18 && x8 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && x22 && ~x23 && ~x15 && x19 && ~x18 && x8 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && x22 && ~x23 && ~x15 && x19 && ~x18 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x65 && ~x21 && x22 && ~x23 && ~x15 && x19 && ~x18 && ~x8 )
						nx_state = s1;
					else if( x65 && ~x21 && x22 && ~x23 && ~x15 && ~x19 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( x65 && ~x21 && ~x22 && x23 && x5 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s28;
						end
					else if( x65 && ~x21 && ~x22 && x23 && ~x5 && x19 && x6 && x16 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( x65 && ~x21 && ~x22 && x23 && ~x5 && x19 && x6 && ~x16 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x65 && ~x21 && ~x22 && x23 && ~x5 && x19 && ~x6 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && x20 && x16 && x6 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s228;
						end
					else if( x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && x20 && x16 && ~x6 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && x20 && ~x16 && x17 && x18 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && x20 && ~x16 && x17 && x18 && ~x6 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && x20 && ~x16 && x17 && ~x18 && x14 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && x20 && ~x16 && x17 && ~x18 && ~x14 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && x20 && ~x16 && ~x17 && x18 && x14 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && x20 && ~x16 && ~x17 && x18 && ~x14 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && x20 && ~x16 && ~x17 && ~x18 && x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && x20 && ~x16 && ~x17 && ~x18 && ~x6 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && ~x20 && x6 )
						begin
							y12 = 1'b1;	
							nx_state = s231;
						end
					else if( x65 && ~x21 && ~x22 && x23 && ~x5 && ~x19 && ~x20 && ~x6 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && x19 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && x19 && x15 && ~x17 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && x19 && ~x15 && x16 && x17 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s157;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && x19 && ~x15 && x16 && ~x17 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y20 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s227;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && x8 && x10 && x17 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && x8 && x10 && ~x17 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && x8 && ~x10 && x11 && x17 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && x8 && ~x10 && x11 && ~x17 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && ~x8 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && ~x19 && x16 && x15 )
						begin
							y18 = 1'b1;	
							nx_state = s203;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && ~x19 && x16 && ~x15 && x17 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && ~x19 && x16 && ~x15 && ~x17 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s233;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && ~x19 && ~x16 && x17 && x15 )
						begin
							y18 = 1'b1;	
							nx_state = s234;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && ~x19 && ~x16 && x17 && ~x15 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s235;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && ~x19 && ~x16 && ~x17 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s236;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && ~x19 && ~x16 && ~x17 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && ~x19 && ~x16 && ~x17 && ~x4 && ~x6 && x15 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s227;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && ~x19 && ~x16 && ~x17 && ~x4 && ~x6 && ~x15 )
						begin
							y16 = 1'b1;	y20 = 1'b1;	
							nx_state = s227;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && x15 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s236;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && x15 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && x15 && ~x4 && ~x6 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s117;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && x17 && x13 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s236;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && x17 && x13 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && x17 && x13 && ~x4 && ~x6 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s227;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && x17 && ~x13 && x16 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s236;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && x17 && ~x13 && x16 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && x17 && ~x13 && x16 && ~x4 && ~x6 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s227;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && x17 && ~x13 && ~x16 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && ~x17 && x16 && x14 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s236;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && ~x17 && x16 && x14 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && ~x17 && x16 && x14 && ~x4 && ~x6 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s227;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && ~x17 && x16 && ~x14 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && x12 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s236;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && x12 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && x12 && ~x4 && ~x6 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s227;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && ~x12 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && ~x19 && x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s236;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && ~x19 && ~x4 && x6 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 && ~x19 && ~x4 && ~x6 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( ~x65 && x66 && x21 && x4 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s28;
						end
					else if( ~x65 && x66 && x21 && ~x4 && x16 && x6 && x15 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s214;
						end
					else if( ~x65 && x66 && x21 && ~x4 && x16 && x6 && x15 && ~x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s215;
						end
					else if( ~x65 && x66 && x21 && ~x4 && x16 && x6 && ~x15 && x10 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && x66 && x21 && ~x4 && x16 && x6 && ~x15 && ~x10 )
						begin
							y14 = 1'b1;	y16 = 1'b1;	
							nx_state = s216;
						end
					else if( ~x65 && x66 && x21 && ~x4 && x16 && ~x6 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s220;
						end
					else if( ~x65 && x66 && x21 && ~x4 && ~x16 && x17 && x10 && x6 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s215;
						end
					else if( ~x65 && x66 && x21 && ~x4 && ~x16 && x17 && x10 && ~x6 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s220;
						end
					else if( ~x65 && x66 && x21 && ~x4 && ~x16 && x17 && ~x10 && x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( ~x65 && x66 && x21 && ~x4 && ~x16 && x17 && ~x10 && ~x6 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s226;
						end
					else if( ~x65 && x66 && x21 && ~x4 && ~x16 && ~x17 && x6 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s215;
						end
					else if( ~x65 && x66 && x21 && ~x4 && ~x16 && ~x17 && x6 && ~x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s218;
						end
					else if( ~x65 && x66 && x21 && ~x4 && ~x16 && ~x17 && ~x6 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	
							nx_state = s220;
						end
					else if( ~x65 && x66 && ~x21 && x22 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s218;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x24 && x26 && x16 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x66 && x24 && x26 && x16 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x66 && x24 && x26 && x16 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x24 && x26 && x16 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x24 && x26 && ~x16 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s165;
						end
					else if( ~x65 && ~x66 && x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && ~x66 && x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && ~x66 && x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x24 && x25 && x26 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x26 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x26 && x19 && ~x14 && ~x13 )
						nx_state = s29;
					else if( ~x65 && ~x66 && ~x24 && x25 && x26 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x26 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x65 && ~x66 && ~x24 && ~x25 && x26 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x65 && ~x66 && ~x24 && ~x25 && ~x26 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s239;
						end
					else nx_state = s29;
				s30 : if( x65 && x66 && x67 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && x67 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && x67 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && x66 && x67 && x22 && ~x17 )
						nx_state = s1;
					else if( x65 && x66 && x67 && ~x22 && x18 && x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && x66 && x67 && ~x22 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && x66 && x67 && ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && x66 && x67 && ~x22 && ~x18 )
						nx_state = s1;
					else if( x65 && x66 && ~x67 && x60 && x61 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x66 && ~x67 && x60 && x61 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x66 && ~x67 && x60 && x61 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x66 && ~x67 && x60 && x61 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x66 && ~x67 && x60 && ~x61 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && ~x67 && x60 && ~x61 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && ~x67 && x60 && ~x61 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x65 && x66 && ~x67 && x60 && ~x61 && ~x18 )
						nx_state = s39;
					else if( x65 && x66 && ~x67 && ~x60 && x61 && x62 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( x65 && x66 && ~x67 && ~x60 && x61 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && ~x67 && ~x60 && x61 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && ~x67 && ~x60 && x61 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x65 && x66 && ~x67 && ~x60 && x61 && ~x62 && ~x18 )
						nx_state = s39;
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 )
						nx_state = s40;
					else if( x65 && ~x66 && x67 && x21 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x65 && ~x66 && x67 && x21 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x65 && ~x66 && x67 && x21 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && x21 && ~x8 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && ~x21 && x23 && x22 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( x65 && ~x66 && x67 && ~x21 && x23 && ~x22 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s240;
						end
					else if( x65 && ~x66 && x67 && ~x21 && ~x23 && x22 && x3 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s240;
						end
					else if( x65 && ~x66 && x67 && ~x21 && ~x23 && x22 && ~x3 && x6 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( x65 && ~x66 && x67 && ~x21 && ~x23 && x22 && ~x3 && x6 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x65 && ~x66 && x67 && ~x21 && ~x23 && x22 && ~x3 && x6 && ~x18 && x19 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x65 && ~x66 && x67 && ~x21 && ~x23 && x22 && ~x3 && x6 && ~x18 && x19 && ~x15 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x65 && ~x66 && x67 && ~x21 && ~x23 && x22 && ~x3 && x6 && ~x18 && ~x19 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( x65 && ~x66 && x67 && ~x21 && ~x23 && x22 && ~x3 && ~x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s28;
						end
					else if( x65 && ~x66 && x67 && ~x21 && ~x23 && ~x22 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( x65 && ~x66 && ~x67 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	y25 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x65 )
						begin
							y6 = 1'b1;	y21 = 1'b1;	y26 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s30;
				s31 : if( x21 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s241;
						end
					else if( ~x21 && x23 && x22 )
						nx_state = s1;
					else if( ~x21 && x23 && ~x22 && x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x21 && x23 && ~x22 && ~x16 && x20 && x19 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x21 && x23 && ~x22 && ~x16 && x20 && ~x19 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x21 && x23 && ~x22 && ~x16 && ~x20 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x21 && ~x23 && x22 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x21 && ~x23 && ~x22 )
						nx_state = s1;
					else nx_state = s31;
				s32 : if( x21 && x18 && x19 && x15 && x17 )
						begin
							y15 = 1'b1;	y20 = 1'b1;	
							nx_state = s227;
						end
					else if( x21 && x18 && x19 && x15 && ~x17 )
						begin
							y16 = 1'b1;	y20 = 1'b1;	
							nx_state = s227;
						end
					else if( x21 && x18 && x19 && ~x15 && x16 && x17 )
						begin
							y18 = 1'b1;	
							nx_state = s203;
						end
					else if( x21 && x18 && x19 && ~x15 && x16 && ~x17 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s233;
						end
					else if( x21 && x18 && x19 && ~x15 && ~x16 && x17 && x10 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x21 && x18 && x19 && ~x15 && ~x16 && x17 && ~x10 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && x18 && x19 && ~x15 && ~x16 && x17 && ~x10 && x8 && ~x9 )
						nx_state = s1;
					else if( x21 && x18 && x19 && ~x15 && ~x16 && x17 && ~x10 && ~x8 )
						nx_state = s1;
					else if( x21 && x18 && x19 && ~x15 && ~x16 && ~x17 && x9 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x21 && x18 && x19 && ~x15 && ~x16 && ~x17 && ~x9 && x8 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && x18 && x19 && ~x15 && ~x16 && ~x17 && ~x9 && x8 && ~x10 )
						nx_state = s1;
					else if( x21 && x18 && x19 && ~x15 && ~x16 && ~x17 && ~x9 && ~x8 )
						nx_state = s1;
					else if( x21 && x18 && ~x19 && x16 && x15 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s243;
						end
					else if( x21 && x18 && ~x19 && x16 && ~x15 && x17 && x14 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s227;
						end
					else if( x21 && x18 && ~x19 && x16 && ~x15 && x17 && ~x14 )
						begin
							y12 = 1'b1;	y19 = 1'b1;	
							nx_state = s230;
						end
					else if( x21 && x18 && ~x19 && x16 && ~x15 && ~x17 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( x21 && x18 && ~x19 && ~x16 && x17 && x15 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s44;
						end
					else if( x21 && x18 && ~x19 && ~x16 && x17 && x15 && ~x3 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x21 && x18 && ~x19 && ~x16 && x17 && x15 && ~x3 && ~x5 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s228;
						end
					else if( x21 && x18 && ~x19 && ~x16 && x17 && ~x15 )
						begin
							y6 = 1'b1;	y19 = 1'b1;	
							nx_state = s223;
						end
					else if( x21 && x18 && ~x19 && ~x16 && ~x17 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s44;
						end
					else if( x21 && x18 && ~x19 && ~x16 && ~x17 && ~x3 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x21 && x18 && ~x19 && ~x16 && ~x17 && ~x3 && ~x5 && x15 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y28 = 1'b1;	
							nx_state = s244;
						end
					else if( x21 && x18 && ~x19 && ~x16 && ~x17 && ~x3 && ~x5 && ~x15 )
						begin
							y18 = 1'b1;	
							nx_state = s234;
						end
					else if( x21 && ~x18 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s44;
						end
					else if( x21 && ~x18 && ~x3 && x19 && x15 && x17 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x21 && ~x18 && ~x3 && x19 && x15 && x17 && ~x5 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s228;
						end
					else if( x21 && ~x18 && ~x3 && x19 && x15 && ~x17 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s245;
						end
					else if( x21 && ~x18 && ~x3 && x19 && x15 && ~x17 && ~x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && x16 && x17 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && x16 && x17 && ~x5 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y20 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s227;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && x16 && ~x17 && x14 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && x16 && ~x17 && x14 && ~x5 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y20 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s227;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && x16 && ~x17 && ~x14 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && x16 && ~x17 && ~x14 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && x16 && ~x17 && ~x14 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && x16 && ~x17 && ~x14 && ~x8 )
						nx_state = s1;
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && x17 && x12 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && x17 && x12 && ~x5 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y20 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s227;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && x17 && ~x12 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && x17 && ~x12 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && x17 && ~x12 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && x17 && ~x12 && ~x8 )
						nx_state = s1;
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && ~x17 && x13 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && ~x17 && x13 && ~x5 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y20 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s227;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && ~x17 && ~x13 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && ~x17 && ~x13 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && ~x17 && ~x13 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x18 && ~x3 && x19 && ~x15 && ~x16 && ~x17 && ~x13 && ~x8 )
						nx_state = s1;
					else if( x21 && ~x18 && ~x3 && ~x19 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( x21 && ~x18 && ~x3 && ~x19 && ~x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x21 && x22 && x23 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x21 && x22 && ~x23 && x15 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x21 && x22 && ~x23 && ~x15 && x19 && x18 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x21 && x22 && ~x23 && ~x15 && x19 && ~x18 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x21 && x22 && ~x23 && ~x15 && ~x19 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x21 && ~x22 && x23 && x4 && x19 && x16 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x21 && ~x22 && x23 && x4 && x19 && ~x16 )
						begin
							y15 = 1'b1;	y20 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x21 && ~x22 && x23 && x4 && ~x19 && x20 && x16 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s117;
						end
					else if( ~x21 && ~x22 && x23 && x4 && ~x19 && x20 && ~x16 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x21 && ~x22 && x23 && x4 && ~x19 && ~x20 )
						begin
							y3 = 1'b1;	y12 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x21 && ~x22 && x23 && ~x4 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x21 && ~x22 && ~x23 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else nx_state = s32;
				s33 : if( x21 && x18 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && x18 && x15 && ~x17 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	
							nx_state = s244;
						end
					else if( x21 && x18 && ~x15 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x21 && ~x18 && x19 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x18 && x19 && x15 && ~x17 )
						begin
							y8 = 1'b1;	
							nx_state = s246;
						end
					else if( x21 && ~x18 && x19 && ~x15 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s227;
						end
					else if( x21 && ~x18 && ~x19 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s31;
						end
					else if( ~x21 && x22 && x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s161;
						end
					else nx_state = s33;
				s34 : if( x21 && x6 && x18 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && x6 && x18 && x15 && ~x17 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	
							nx_state = s244;
						end
					else if( x21 && x6 && x18 && ~x15 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x21 && x6 && ~x18 && x19 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && x6 && ~x18 && x19 && x15 && ~x17 )
						begin
							y8 = 1'b1;	
							nx_state = s246;
						end
					else if( x21 && x6 && ~x18 && x19 && ~x15 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s227;
						end
					else if( x21 && x6 && ~x18 && ~x19 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s31;
						end
					else if( x21 && ~x6 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x21 && x23 && x22 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( ~x21 && x23 && x22 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x21 && x23 && x22 && ~x18 && x19 && x15 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x21 && x23 && x22 && ~x18 && x19 && ~x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( ~x21 && x23 && x22 && ~x18 && ~x19 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s33;
						end
					else if( ~x21 && x23 && ~x22 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s161;
						end
					else if( ~x21 && ~x23 && x22 )
						nx_state = s1;
					else if( ~x21 && ~x23 && ~x22 )
						begin
							y12 = 1'b1;	y19 = 1'b1;	
							nx_state = s230;
						end
					else nx_state = s34;
				s35 : if( 1'b1 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else nx_state = s35;
				s36 : if( x21 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s240;
						end
					else if( ~x21 && x22 && x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( ~x21 && x22 && ~x23 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && ~x19 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x23 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s161;
						end
					else nx_state = s36;
				s37 : if( x13 && x17 && x21 && x16 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s249;
						end
					else if( x13 && x17 && x21 && ~x16 && x18 && x15 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s249;
						end
					else if( x13 && x17 && x21 && ~x16 && x18 && ~x15 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else if( x13 && x17 && x21 && ~x16 && ~x18 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s249;
						end
					else if( x13 && x17 && ~x21 && x22 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s249;
						end
					else if( x13 && x17 && ~x21 && ~x22 && x15 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s249;
						end
					else if( x13 && x17 && ~x21 && ~x22 && ~x15 && x19 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s249;
						end
					else if( x13 && x17 && ~x21 && ~x22 && ~x15 && ~x19 && x20 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s249;
						end
					else if( x13 && x17 && ~x21 && ~x22 && ~x15 && ~x19 && ~x20 && x16 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s249;
						end
					else if( x13 && x17 && ~x21 && ~x22 && ~x15 && ~x19 && ~x20 && ~x16 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else if( x13 && ~x17 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s249;
						end
					else nx_state = s37;
				s38 : if( x66 && x15 && x12 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x66 && x15 && x12 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s250;
						end
					else if( x66 && x15 && ~x12 && x7 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x15 && ~x12 && ~x7 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( x66 && ~x15 && x16 && x7 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s251;
						end
					else if( x66 && ~x15 && x16 && x7 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( x66 && ~x15 && x16 && ~x7 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s252;
						end
					else if( x66 && ~x15 && ~x16 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s253;
						end
					else if( x66 && ~x15 && ~x16 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x66 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else nx_state = s38;
				s39 : if( x65 )
						nx_state = s1;
					else if( ~x65 && x20 )
						nx_state = s1;
					else if( ~x65 && ~x20 && x21 && x15 && x8 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x65 && ~x20 && x21 && x15 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x16 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s209;
						end
					else if( ~x65 && ~x20 && ~x21 )
						begin
							y3 = 1'b1;	y20 = 1'b1;	
							nx_state = s42;
						end
					else nx_state = s39;
				s40 : if( x66 && x65 && x60 && x61 && x15 && x2 && x12 && x7 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s67;
						end
					else if( x66 && x65 && x60 && x61 && x15 && x2 && x12 && ~x7 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s131;
						end
					else if( x66 && x65 && x60 && x61 && x15 && x2 && ~x12 && x7 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s255;
						end
					else if( x66 && x65 && x60 && x61 && x15 && x2 && ~x12 && ~x7 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s254;
						end
					else if( x66 && x65 && x60 && x61 && x15 && ~x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s255;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && x16 && x7 && x12 && x2 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s256;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && x16 && x7 && x12 && ~x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s255;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && x16 && x7 && ~x12 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s255;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && x12 && x9 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s255;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && x12 && ~x9 && x11 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s255;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && x12 && ~x9 && ~x11 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && x12 && ~x9 && ~x11 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && x12 && ~x9 && ~x11 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && x12 && ~x9 && ~x11 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && ~x12 && x11 && x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s255;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && ~x12 && x11 && ~x10 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && ~x12 && x11 && ~x10 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && ~x12 && x11 && ~x10 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && ~x12 && x11 && ~x10 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && ~x12 && ~x11 && x8 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s255;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && ~x12 && ~x11 && ~x8 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && ~x12 && ~x11 && ~x8 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && ~x12 && ~x11 && ~x8 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && x16 && ~x7 && ~x12 && ~x11 && ~x8 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && ~x16 && x2 && x7 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s257;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && ~x16 && x2 && ~x7 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( x66 && x65 && x60 && x61 && ~x15 && ~x16 && ~x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s255;
						end
					else if( x66 && x65 && x60 && ~x61 && x11 )
						nx_state = s1;
					else if( x66 && x65 && x60 && ~x61 && ~x11 && x7 )
						nx_state = s1;
					else if( x66 && x65 && x60 && ~x61 && ~x11 && ~x7 && x16 && x15 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && x65 && x60 && ~x61 && ~x11 && ~x7 && x16 && x15 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && x65 && x60 && ~x61 && ~x11 && ~x7 && x16 && x15 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x66 && x65 && x60 && ~x61 && ~x11 && ~x7 && x16 && x15 && ~x18 )
						nx_state = s39;
					else if( x66 && x65 && x60 && ~x61 && ~x11 && ~x7 && x16 && ~x15 )
						nx_state = s1;
					else if( x66 && x65 && x60 && ~x61 && ~x11 && ~x7 && ~x16 )
						nx_state = s1;
					else if( x66 && x65 && ~x60 && x61 && x62 && x16 && x11 && x12 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x66 && x65 && ~x60 && x61 && x62 && x16 && x11 && ~x12 && x13 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x66 && x65 && ~x60 && x61 && x62 && x16 && x11 && ~x12 && ~x13 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s154;
						end
					else if( x66 && x65 && ~x60 && x61 && x62 && x16 && ~x11 && x13 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s63;
						end
					else if( x66 && x65 && ~x60 && x61 && x62 && x16 && ~x11 && ~x13 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( x66 && x65 && ~x60 && x61 && x62 && ~x16 && x17 && x11 && x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s258;
						end
					else if( x66 && x65 && ~x60 && x61 && x62 && ~x16 && x17 && x11 && ~x13 && x2 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x66 && x65 && ~x60 && x61 && x62 && ~x16 && x17 && x11 && ~x13 && ~x2 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( x66 && x65 && ~x60 && x61 && x62 && ~x16 && x17 && ~x11 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s258;
						end
					else if( x66 && x65 && ~x60 && x61 && x62 && ~x16 && ~x17 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( x66 && x65 && ~x60 && x61 && ~x62 && x11 )
						nx_state = s1;
					else if( x66 && x65 && ~x60 && x61 && ~x62 && ~x11 && x7 )
						nx_state = s1;
					else if( x66 && x65 && ~x60 && x61 && ~x62 && ~x11 && ~x7 && x16 && x15 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && x65 && ~x60 && x61 && ~x62 && ~x11 && ~x7 && x16 && x15 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && x65 && ~x60 && x61 && ~x62 && ~x11 && ~x7 && x16 && x15 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x66 && x65 && ~x60 && x61 && ~x62 && ~x11 && ~x7 && x16 && x15 && ~x18 )
						nx_state = s39;
					else if( x66 && x65 && ~x60 && x61 && ~x62 && ~x11 && ~x7 && x16 && ~x15 )
						nx_state = s1;
					else if( x66 && x65 && ~x60 && x61 && ~x62 && ~x11 && ~x7 && ~x16 )
						nx_state = s1;
					else if( x66 && x65 && ~x60 && ~x61 && x62 && x18 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && x65 && ~x60 && ~x61 && x62 && x18 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && x65 && ~x60 && ~x61 && x62 && x18 && ~x13 && ~x14 )
						nx_state = s1;
					else if( x66 && x65 && ~x60 && ~x61 && x62 && ~x18 )
						nx_state = s1;
					else if( x66 && x65 && ~x60 && ~x61 && ~x62 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && x65 && ~x60 && ~x61 && ~x62 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && x65 && ~x60 && ~x61 && ~x62 && x19 && ~x13 && ~x14 )
						nx_state = s1;
					else if( x66 && x65 && ~x60 && ~x61 && ~x62 && ~x19 )
						nx_state = s1;
					else if( x66 && ~x65 && x21 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x21 && x22 && x23 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x66 && ~x65 && ~x21 && x22 && ~x23 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x21 && ~x22 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( x66 && ~x65 && ~x21 && ~x22 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( x66 && ~x65 && ~x21 && ~x22 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x21 && ~x22 && x23 && ~x19 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x21 && ~x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x66 && x65 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x4 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && x20 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && ~x20 && x21 )
						nx_state = s39;
					else if( ~x66 && ~x65 && x67 && ~x20 && ~x21 && x18 && x15 && x8 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x66 && ~x65 && x67 && ~x20 && ~x21 && x18 && x15 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x66 && ~x65 && x67 && ~x20 && ~x21 && x18 && ~x15 && x16 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && ~x65 && x67 && ~x20 && ~x21 && x18 && ~x15 && ~x16 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s209;
						end
					else if( ~x66 && ~x65 && x67 && ~x20 && ~x21 && ~x18 )
						nx_state = s39;
					else if( ~x66 && ~x65 && ~x67 && x21 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && x3 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y9 = 1'b1;	
							nx_state = s107;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && x3 && ~x2 )
						nx_state = s40;
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x3 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && x2 && x11 )
						nx_state = s40;
					else if( ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && x2 && ~x11 )
						nx_state = s40;
					else if( ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else nx_state = s40;
				s41 : if( x20 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x20 && x21 && x15 && x8 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x20 && x21 && x15 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x20 && x21 && ~x15 && x16 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x20 && x21 && ~x15 && ~x16 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s209;
						end
					else if( ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else nx_state = s41;
				s42 : if( x21 )
						nx_state = s1;
					else if( ~x21 && x15 && x8 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x21 && x15 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x21 && ~x15 && x16 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x21 && ~x15 && ~x16 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s209;
						end
					else nx_state = s42;
				s43 : if( x65 && x66 && x68 && x21 && x20 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s259;
						end
					else if( x65 && x66 && x68 && x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x66 && x68 && x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x66 && x68 && x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x66 && x68 && x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( x65 && x66 && x68 && ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x66 && x68 && ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x66 && x68 && ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x66 && x68 && ~x21 && ~x19 )
						nx_state = s1;
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && x7 && x12 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && x7 && ~x12 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s260;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && ~x7 && x12 && x14 && x11 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s261;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && ~x7 && x12 && x14 && ~x11 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && ~x7 && x12 && ~x14 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && ~x7 && x12 && ~x14 && x19 && ~x13 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && ~x7 && x12 && ~x14 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && ~x7 && ~x12 && x13 && x11 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s262;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && ~x7 && ~x12 && x13 && ~x11 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && ~x7 && ~x12 && ~x13 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && ~x7 && ~x12 && ~x13 && x19 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && x16 && ~x7 && ~x12 && ~x13 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && x11 && x7 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && x11 && ~x7 && x12 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && x11 && ~x7 && ~x12 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s257;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && ~x11 && x1 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && ~x11 && ~x1 && x12 && x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s74;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && ~x11 && ~x1 && x12 && ~x3 && x7 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s69;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && ~x11 && ~x1 && x12 && ~x3 && ~x7 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s257;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && ~x11 && ~x1 && ~x12 && x7 && x3 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s263;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && ~x11 && ~x1 && ~x12 && x7 && ~x3 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && ~x11 && ~x1 && ~x12 && ~x7 && x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s74;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && x15 && ~x16 && ~x11 && ~x1 && ~x12 && ~x7 && ~x3 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && x1 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && x7 && x12 && x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s74;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && x7 && x12 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s257;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && x7 && ~x12 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s74;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && x12 && x11 && x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s74;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && x12 && x11 && ~x3 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && x12 && ~x11 && x9 && x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s74;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && x12 && ~x11 && x9 && ~x3 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && x12 && ~x11 && ~x9 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && x12 && ~x11 && ~x9 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && x12 && ~x11 && ~x9 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && x12 && ~x11 && ~x9 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && x11 && x10 && x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s74;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && x11 && x10 && ~x3 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && x11 && ~x10 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && x11 && ~x10 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && x11 && ~x10 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && x11 && ~x10 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && ~x11 && x8 && x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s74;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && ~x11 && x8 && ~x3 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && ~x11 && ~x8 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && ~x11 && ~x8 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && ~x11 && ~x8 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && x16 && ~x7 && ~x12 && ~x11 && ~x8 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && ~x16 && x3 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s74;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && ~x16 && ~x3 && x7 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s257;
						end
					else if( x65 && x66 && ~x68 && x61 && x60 && ~x15 && ~x1 && ~x16 && ~x3 && ~x7 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s264;
						end
					else if( x65 && x66 && ~x68 && x61 && ~x60 && x62 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && x66 && ~x68 && x61 && ~x60 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && ~x68 && x61 && ~x60 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && ~x68 && x61 && ~x60 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x65 && x66 && ~x68 && x61 && ~x60 && ~x62 && ~x18 )
						nx_state = s39;
					else if( x65 && x66 && ~x68 && ~x61 && x60 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && ~x68 && ~x61 && x60 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && ~x68 && ~x61 && x60 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x65 && x66 && ~x68 && ~x61 && x60 && ~x18 )
						nx_state = s39;
					else if( x65 && x66 && ~x68 && ~x61 && ~x60 && x62 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( x65 && x66 && ~x68 && ~x61 && ~x60 && ~x62 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && ~x66 && x68 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && x68 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && x68 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x66 && x68 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x68 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x65 && ~x66 && ~x68 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x68 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x68 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x68 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x68 && ~x21 && x23 && x22 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x23 && x22 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x68 && ~x21 && x23 && x22 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x68 && ~x21 && x23 && ~x22 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x23 && ~x22 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x23 && ~x22 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x68 && ~x21 && x23 && ~x22 && ~x20 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x68 && ~x21 && ~x23 && x18 && x14 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && ~x23 && x18 && x14 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && ~x23 && x18 && ~x14 && x13 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && ~x23 && x18 && ~x14 && x13 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x68 && ~x21 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x67 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x67 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x67 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x67 && x20 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x67 && ~x20 )
						nx_state = s1;
					else if( ~x65 && ~x67 && x21 && x68 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x65 && ~x67 && x21 && x68 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x65 && ~x67 && x21 && x68 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x65 && ~x67 && x21 && x68 && ~x3 )
						nx_state = s1;
					else if( ~x65 && ~x67 && x21 && ~x68 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && x12 && x17 )
						begin
							y8 = 1'b1;	
							nx_state = s246;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && x12 && ~x17 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && ~x12 && x17 && x8 && x16 )
						begin
							y8 = 1'b1;	y22 = 1'b1;	
							nx_state = s267;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && ~x12 && x17 && x8 && ~x16 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s268;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && ~x12 && x17 && ~x8 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && ~x12 && x17 && ~x8 && x6 && ~x7 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && ~x12 && x17 && ~x8 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && ~x12 && ~x17 && x7 && x16 )
						begin
							y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s269;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && ~x12 && ~x17 && x7 && ~x16 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s268;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && ~x12 && ~x17 && ~x7 && x6 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && ~x12 && ~x17 && ~x7 && x6 && ~x8 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && x19 && ~x12 && ~x17 && ~x7 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && ~x19 && x16 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s270;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && ~x19 && x16 && ~x12 && x17 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && ~x19 && x16 && ~x12 && ~x17 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && ~x19 && ~x16 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && ~x19 && ~x16 && ~x2 && x3 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && ~x19 && ~x16 && ~x2 && ~x3 && x17 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s272;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && ~x19 && ~x16 && ~x2 && ~x3 && x17 && ~x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s272;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && ~x19 && ~x16 && ~x2 && ~x3 && ~x17 && x12 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && x18 && ~x19 && ~x16 && ~x2 && ~x3 && ~x17 && ~x12 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && x12 && x3 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && x12 && ~x3 && x17 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && x12 && ~x3 && ~x17 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && x16 && x17 && x3 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && x16 && x17 && ~x3 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && x16 && ~x17 && x15 && x3 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && x16 && ~x17 && x15 && ~x3 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && x16 && ~x17 && ~x15 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && x16 && ~x17 && ~x15 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && x16 && ~x17 && ~x15 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && x16 && ~x17 && ~x15 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && x17 && x14 && x3 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && x17 && x14 && ~x3 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && x17 && ~x14 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && x17 && ~x14 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && x17 && ~x14 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && x17 && ~x14 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && ~x17 && x13 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && ~x17 && x13 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && ~x17 && x13 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && ~x17 && x13 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && ~x17 && ~x13 && x3 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && x19 && ~x12 && ~x16 && ~x17 && ~x13 && ~x3 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && ~x19 && x3 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && ~x19 && ~x3 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x68 && ~x18 && ~x2 && ~x19 && ~x3 && ~x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s272;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && ~x68 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s126;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && x15 && x17 )
						begin
							y8 = 1'b1;	
							nx_state = s246;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && x15 && ~x17 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && ~x15 && x16 && x17 )
						begin
							y8 = 1'b1;	y22 = 1'b1;	
							nx_state = s267;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && ~x15 && x16 && ~x17 )
						begin
							y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s269;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && ~x15 && ~x16 && x17 && x10 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && ~x15 && ~x16 && x17 && ~x10 && x9 && x8 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && ~x15 && ~x16 && x17 && ~x10 && x9 && ~x8 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && ~x15 && ~x16 && x17 && ~x10 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && ~x15 && ~x16 && ~x17 && x9 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && ~x15 && ~x16 && ~x17 && ~x9 && x8 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && ~x15 && ~x16 && ~x17 && ~x9 && x8 && ~x10 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && x19 && ~x15 && ~x16 && ~x17 && ~x9 && ~x8 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && ~x19 && x16 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s274;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && ~x19 && ~x16 && x2 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s173;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && ~x19 && ~x16 && ~x2 && x5 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s275;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && ~x19 && ~x16 && ~x2 && ~x5 && x15 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && x18 && ~x19 && ~x16 && ~x2 && ~x5 && ~x15 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && x2 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s173;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && x15 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s275;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && x16 && x17 && x5 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s275;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && x16 && x17 && ~x5 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && x16 && ~x17 && x14 && x5 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s275;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && x16 && ~x17 && x14 && ~x5 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && x16 && ~x17 && ~x14 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && x16 && ~x17 && ~x14 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && x16 && ~x17 && ~x14 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && x16 && ~x17 && ~x14 && ~x8 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && x17 && x13 && x5 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s275;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && x17 && x13 && ~x5 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && x17 && ~x13 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && x17 && ~x13 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && x17 && ~x13 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && x17 && ~x13 && ~x8 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && ~x17 && x12 && x5 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s275;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && ~x17 && x12 && ~x5 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && ~x17 && ~x12 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && ~x17 && ~x12 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && ~x17 && ~x12 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && x19 && ~x15 && ~x16 && ~x17 && ~x12 && ~x8 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && ~x19 && x5 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s275;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x18 && ~x2 && ~x19 && ~x5 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s274;
						end
					else if( ~x65 && ~x67 && ~x21 && ~x22 && ~x68 )
						nx_state = s1;
					else nx_state = s43;
				s44 : if( x65 && x66 && x67 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x65 && x66 && ~x67 && x21 && x20 )
						begin
							y9 = 1'b1;	y24 = 1'b1;	
							nx_state = s276;
						end
					else if( x65 && x66 && ~x67 && x21 && ~x20 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( x65 && x66 && ~x67 && ~x21 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( x65 && ~x66 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x65 && x20 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( ~x65 && ~x20 && x21 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y21 = 1'b1;	
							nx_state = s45;
						end
					else if( ~x65 && ~x20 && ~x21 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else nx_state = s44;
				s45 : if( x20 )
						nx_state = s1;
					else if( ~x20 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	
							nx_state = s277;
						end
					else nx_state = s45;
				s46 : if( x24 && x26 && x19 )
						nx_state = s46;
					else if( x24 && x26 && ~x19 )
						nx_state = s1;
					else if( x24 && ~x26 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else if( ~x24 && x25 && x26 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x26 && x15 && x6 && x10 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x24 && x25 && ~x26 && x15 && x6 && x10 && ~x11 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s172;
						end
					else if( ~x24 && x25 && ~x26 && x15 && x6 && x10 && ~x11 && ~x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x24 && x25 && ~x26 && x15 && x6 && ~x10 )
						begin
							y8 = 1'b1;	y17 = 1'b1;	y23 = 1'b1;	
							nx_state = s164;
						end
					else if( ~x24 && x25 && ~x26 && x15 && ~x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && x10 && x8 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && x10 && ~x8 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && x10 && ~x8 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && x10 && ~x8 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && x10 && ~x8 && ~x19 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && ~x10 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && ~x10 && ~x7 && x11 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && ~x10 && ~x7 && ~x11 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && ~x10 && ~x7 && ~x11 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && ~x10 && ~x7 && ~x11 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && x12 && ~x10 && ~x7 && ~x11 && ~x19 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && ~x10 && x11 && x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && ~x10 && x11 && ~x9 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && ~x10 && x11 && ~x9 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && ~x10 && x11 && ~x9 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && ~x10 && x11 && ~x9 && ~x19 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && ~x10 && ~x11 && x8 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && ~x10 && ~x11 && x8 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && ~x10 && ~x11 && x8 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && ~x10 && ~x11 && x8 && ~x19 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x26 && ~x15 && x16 && ~x12 && ~x10 && ~x11 && ~x8 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && ~x16 && x6 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x24 && x25 && ~x26 && ~x15 && ~x16 && ~x6 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x24 && ~x25 && x26 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else if( ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else nx_state = s46;
				s47 : if( x68 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x68 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x68 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x68 && x20 && ~x18 )
						nx_state = s1;
					else if( x68 && ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( x68 && ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( x68 && ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x68 && ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( x68 && ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( x68 && ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( x68 && ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x68 && ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else if( ~x68 && x24 && x26 )
						begin
							y17 = 1'b1;	
							nx_state = s279;
						end
					else if( ~x68 && x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x68 && x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x68 && x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x68 && x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x68 && ~x24 && x25 && x26 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x68 && ~x24 && x25 && ~x26 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 )
						nx_state = s1;
					else if( ~x68 && ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x68 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x68 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x68 && ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else nx_state = s47;
				s48 : if( x66 && x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x66 && x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x66 && x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && x21 && ~x18 )
						nx_state = s1;
					else if( x66 && ~x21 && x22 && x23 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x66 && ~x21 && x22 && ~x23 && x18 && x14 )
						nx_state = s40;
					else if( x66 && ~x21 && x22 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s40;
					else if( x66 && ~x21 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && ~x21 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( x66 && ~x21 && ~x22 && x23 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( x66 && ~x21 && ~x22 && ~x23 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s180;
						end
					else if( ~x66 && x24 && x26 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x66 && x24 && x26 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x66 && x24 && x26 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x66 && x24 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x66 && x24 && ~x26 )
						nx_state = s1;
					else if( ~x66 && ~x24 && x25 && x26 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x66 && ~x24 && x25 && x26 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x66 && ~x24 && x25 && x26 && x19 && ~x14 && ~x13 )
						nx_state = s48;
					else if( ~x66 && ~x24 && x25 && x26 && ~x19 )
						nx_state = s1;
					else if( ~x66 && ~x24 && x25 && ~x26 )
						nx_state = s1;
					else if( ~x66 && ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x66 && ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x66 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x66 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else nx_state = s48;
				s49 : if( x24 && x26 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( x24 && x26 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( x24 && x26 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x24 && x26 && ~x18 )
						nx_state = s1;
					else if( x24 && ~x26 )
						nx_state = s1;
					else if( ~x24 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x25 && x19 && ~x14 && ~x13 && x26 )
						nx_state = s49;
					else if( ~x24 && x25 && x19 && ~x14 && ~x13 && ~x26 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else nx_state = s49;
				s50 : if( x65 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && x22 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x22 && x18 && x13 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && ~x22 && x18 && x13 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && ~x22 && x18 && ~x13 && x12 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && ~x22 && x18 && ~x13 && x12 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && ~x22 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x26 && x24 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x65 && x26 && ~x24 && x25 )
						nx_state = s1;
					else if( ~x65 && x26 && ~x24 && ~x25 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x65 && x26 && ~x24 && ~x25 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x65 && x26 && ~x24 && ~x25 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x26 && ~x24 && ~x25 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x26 && x24 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s280;
						end
					else if( ~x65 && ~x26 && ~x24 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x26 && ~x24 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x26 && ~x24 && x25 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x26 && ~x24 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x26 && ~x24 && ~x25 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x65 && ~x26 && ~x24 && ~x25 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x65 && ~x26 && ~x24 && ~x25 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x26 && ~x24 && ~x25 && ~x17 )
						nx_state = s1;
					else nx_state = s50;
				s51 : if( x65 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x4 )
						nx_state = s1;
					else if( ~x65 && x24 && x26 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x65 && ~x24 && x25 && x26 )
						begin
							y11 = 1'b1;	y16 = 1'b1;	y25 = 1'b1;	
							nx_state = s281;
						end
					else if( ~x65 && ~x24 && x25 && ~x26 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && ~x24 && ~x25 && x26 && x3 && x16 && x11 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s46;
						end
					else if( ~x65 && ~x24 && ~x25 && x26 && x3 && x16 && ~x11 && x12 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s46;
						end
					else if( ~x65 && ~x24 && ~x25 && x26 && x3 && x16 && ~x11 && ~x12 && x10 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x24 && ~x25 && x26 && x3 && x16 && ~x11 && ~x12 && ~x10 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && ~x24 && ~x25 && x26 && x3 && ~x16 && x17 && x10 && x12 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( ~x65 && ~x24 && ~x25 && x26 && x3 && ~x16 && x17 && x10 && ~x12 )
						begin
							y17 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x65 && ~x24 && ~x25 && x26 && x3 && ~x16 && x17 && ~x10 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( ~x65 && ~x24 && ~x25 && x26 && x3 && ~x16 && ~x17 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s46;
						end
					else if( ~x65 && ~x24 && ~x25 && x26 && ~x3 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x24 && ~x25 && ~x26 && x4 && x15 && x11 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else if( ~x65 && ~x24 && ~x25 && ~x26 && x4 && x15 && ~x11 && x12 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else if( ~x65 && ~x24 && ~x25 && ~x26 && x4 && x15 && ~x11 && ~x12 && x10 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x65 && ~x24 && ~x25 && ~x26 && x4 && x15 && ~x11 && ~x12 && ~x10 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && ~x24 && ~x25 && ~x26 && x4 && ~x15 && x16 && x10 && x12 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x65 && ~x24 && ~x25 && ~x26 && x4 && ~x15 && x16 && x10 && ~x12 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s239;
						end
					else if( ~x65 && ~x24 && ~x25 && ~x26 && x4 && ~x15 && x16 && ~x10 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x65 && ~x24 && ~x25 && ~x26 && x4 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else if( ~x65 && ~x24 && ~x25 && ~x26 && ~x4 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s165;
						end
					else nx_state = s51;
				s52 : if( x66 && x21 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( x66 && ~x21 && x22 && x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s219;
						end
					else if( x66 && ~x21 && x22 && ~x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s28;
						end
					else if( x66 && ~x21 && ~x22 )
						begin
							y8 = 1'b1;	y18 = 1'b1;	
							nx_state = s82;
						end
					else if( ~x66 && x24 && x11 && x26 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && x24 && x11 && ~x26 && x13 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x66 && x24 && x11 && ~x26 && x13 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x66 && x24 && x11 && ~x26 && x13 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x66 && x24 && x11 && ~x26 && x13 && ~x20 )
						nx_state = s1;
					else if( ~x66 && x24 && x11 && ~x26 && ~x13 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s282;
						end
					else if( ~x66 && x24 && ~x11 && x26 && x12 && x13 && x16 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x66 && x24 && ~x11 && x26 && x12 && x13 && x16 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x66 && x24 && ~x11 && x26 && x12 && x13 && x16 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x66 && x24 && ~x11 && x26 && x12 && x13 && x16 && ~x18 )
						nx_state = s1;
					else if( ~x66 && x24 && ~x11 && x26 && x12 && x13 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && x24 && ~x11 && x26 && x12 && ~x13 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && x24 && ~x11 && x26 && ~x12 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && x24 && ~x11 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x66 && x24 && ~x11 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x66 && x24 && ~x11 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x66 && x24 && ~x11 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x66 && ~x24 && x25 && x26 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && ~x24 && x25 && ~x26 )
						nx_state = s1;
					else if( ~x66 && ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x66 && ~x24 && ~x25 && ~x26 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else nx_state = s52;
				s53 : if( x66 && x67 && x65 && x22 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	
							nx_state = s111;
						end
					else if( x66 && x67 && x65 && ~x22 && x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x66 && x67 && x65 && ~x22 && ~x23 && x18 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x67 && x65 && ~x22 && ~x23 && x18 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x67 && x65 && ~x22 && ~x23 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x66 && x67 && x65 && ~x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( x66 && x67 && ~x65 && x63 && x15 && x64 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( x66 && x67 && ~x65 && x63 && x15 && x64 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x66 && x67 && ~x65 && x63 && x15 && ~x64 && x16 && x8 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x67 && ~x65 && x63 && x15 && ~x64 && x16 && x8 && ~x14 && x7 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s157;
						end
					else if( x66 && x67 && ~x65 && x63 && x15 && ~x64 && x16 && x8 && ~x14 && ~x7 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s65;
						end
					else if( x66 && x67 && ~x65 && x63 && x15 && ~x64 && x16 && x8 && ~x14 && ~x7 && ~x12 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( x66 && x67 && ~x65 && x63 && x15 && ~x64 && x16 && ~x8 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && x67 && ~x65 && x63 && x15 && ~x64 && x16 && ~x8 && ~x14 && x7 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s158;
						end
					else if( x66 && x67 && ~x65 && x63 && x15 && ~x64 && x16 && ~x8 && ~x14 && ~x7 && x13 )
						begin
							y3 = 1'b1;	
							nx_state = s65;
						end
					else if( x66 && x67 && ~x65 && x63 && x15 && ~x64 && x16 && ~x8 && ~x14 && ~x7 && ~x13 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( x66 && x67 && ~x65 && x63 && x15 && ~x64 && ~x16 && x7 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s159;
						end
					else if( x66 && x67 && ~x65 && x63 && x15 && ~x64 && ~x16 && ~x7 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( x66 && x67 && ~x65 && x63 && x15 && ~x64 && ~x16 && ~x7 && ~x3 && x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( x66 && x67 && ~x65 && x63 && x15 && ~x64 && ~x16 && ~x7 && ~x3 && ~x5 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x66 && x67 && ~x65 && x63 && x15 && ~x64 && ~x16 && ~x7 && ~x3 && ~x5 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && x16 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s151;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && x8 && x7 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && x8 && x7 && ~x3 && x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && x8 && x7 && ~x3 && ~x5 )
						begin
							y21 = 1'b1;	
							nx_state = s151;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && x8 && ~x7 && x9 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && x8 && ~x7 && x9 && ~x3 && x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && x8 && ~x7 && x9 && ~x3 && ~x5 )
						begin
							y21 = 1'b1;	
							nx_state = s151;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && x8 && ~x7 && ~x9 && x3 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && x8 && ~x7 && ~x9 && ~x3 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && ~x8 && x7 && x11 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && ~x8 && x7 && x11 && ~x3 && x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && ~x8 && x7 && x11 && ~x3 && ~x5 )
						begin
							y21 = 1'b1;	
							nx_state = s151;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && ~x8 && x7 && ~x11 && x3 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && ~x8 && x7 && ~x11 && ~x3 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && ~x8 && ~x7 && x10 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && ~x8 && ~x7 && x10 && ~x3 && x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && ~x8 && ~x7 && x10 && ~x3 && ~x5 )
						begin
							y21 = 1'b1;	
							nx_state = s151;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && ~x8 && ~x7 && ~x10 && x3 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && x16 && ~x64 && ~x8 && ~x7 && ~x10 && ~x3 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && ~x16 && x64 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s135;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && ~x16 && ~x64 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && ~x16 && ~x64 && ~x3 && x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( x66 && x67 && ~x65 && x63 && ~x15 && ~x16 && ~x64 && ~x3 && ~x5 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y28 = 1'b1;	
							nx_state = s135;
						end
					else if( x66 && x67 && ~x65 && ~x63 && x64 && x19 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x66 && x67 && ~x65 && ~x63 && x64 && x19 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x66 && x67 && ~x65 && ~x63 && x64 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x66 && x67 && ~x65 && ~x63 && x64 && ~x19 )
						nx_state = s1;
					else if( x66 && x67 && ~x65 && ~x63 && ~x64 )
						nx_state = s1;
					else if( x66 && ~x67 && x65 && x61 && x60 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && ~x67 && x65 && x61 && x60 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && ~x67 && x65 && x61 && x60 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x66 && ~x67 && x65 && x61 && x60 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x66 && ~x67 && x65 && x61 && ~x60 && x62 && x11 && x13 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x66 && ~x67 && x65 && x61 && ~x60 && x62 && x11 && x13 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x66 && ~x67 && x65 && x61 && ~x60 && x62 && x11 && x13 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x66 && ~x67 && x65 && x61 && ~x60 && x62 && x11 && x13 && ~x18 )
						nx_state = s1;
					else if( x66 && ~x67 && x65 && x61 && ~x60 && x62 && x11 && ~x13 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( x66 && ~x67 && x65 && x61 && ~x60 && x62 && ~x11 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x66 && ~x67 && x65 && x61 && ~x60 && x62 && ~x11 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x66 && ~x67 && x65 && x61 && ~x60 && x62 && ~x11 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x66 && ~x67 && x65 && x61 && ~x60 && x62 && ~x11 && ~x18 )
						nx_state = s1;
					else if( x66 && ~x67 && x65 && x61 && ~x60 && ~x62 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x66 && ~x67 && x65 && x61 && ~x60 && ~x62 && ~x7 )
						nx_state = s39;
					else if( x66 && ~x67 && x65 && ~x61 && x60 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x66 && ~x67 && x65 && ~x61 && x60 && ~x7 )
						nx_state = s39;
					else if( x66 && ~x67 && x65 && ~x61 && ~x60 && x62 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( x66 && ~x67 && x65 && ~x61 && ~x60 && ~x62 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s258;
						end
					else if( x66 && ~x67 && ~x65 && x21 && x68 && x9 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x66 && ~x67 && ~x65 && x21 && x68 && x9 && ~x8 && x7 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x66 && ~x67 && ~x65 && x21 && x68 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && x21 && x68 && ~x9 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && x21 && ~x68 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x66 && ~x67 && ~x65 && x21 && ~x68 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x66 && ~x67 && ~x65 && x21 && ~x68 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && x21 && ~x68 && ~x18 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && x5 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && x17 && x10 && x15 && x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s283;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && x17 && x10 && x15 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && x17 && x10 && ~x15 && x16 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && x17 && x10 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && x17 && ~x10 && x6 )
						begin
							y13 = 1'b1;	y16 = 1'b1;	
							nx_state = s284;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && x17 && ~x10 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && ~x17 && x18 && x6 && x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s219;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && ~x17 && x18 && x6 && ~x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && ~x17 && x18 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && ~x17 && ~x18 && x6 && x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s219;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && ~x17 && ~x18 && x6 && ~x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s28;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && x68 && ~x5 && ~x17 && ~x18 && ~x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && x23 && x18 && x15 && x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && x23 && x18 && x15 && ~x10 && x12 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && x23 && x18 && x15 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s285;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && x23 && x18 && ~x15 && x16 && x10 && x12 )
						begin
							y14 = 1'b1;	
							nx_state = s286;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && x23 && x18 && ~x15 && x16 && x10 && ~x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && x23 && x18 && ~x15 && x16 && ~x10 )
						begin
							y14 = 1'b1;	
							nx_state = s286;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && x23 && x18 && ~x15 && ~x16 )
						nx_state = s40;
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && x23 && ~x18 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && ~x23 && x18 && x14 )
						nx_state = s40;
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s40;
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && x22 && ~x68 && ~x23 && ~x18 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && x10 && x15 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && x10 && ~x15 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && ~x10 && x15 && x6 && x14 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && ~x10 && x15 && x6 && ~x14 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s287;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && ~x10 && x15 && ~x6 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && ~x10 && x15 && ~x6 && x4 && ~x5 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && ~x10 && x15 && ~x6 && ~x4 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && ~x10 && ~x15 && x5 && x14 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s288;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && ~x10 && ~x15 && x5 && ~x14 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s287;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && ~x10 && ~x15 && ~x5 && x4 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && ~x10 && ~x15 && ~x5 && x4 && ~x6 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && x17 && ~x10 && ~x15 && ~x5 && ~x4 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && x14 && x10 )
						begin
							y13 = 1'b1;	y16 = 1'b1;	
							nx_state = s289;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && x14 && ~x10 && x15 )
						begin
							y13 = 1'b1;	y16 = 1'b1;	
							nx_state = s284;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && x14 && ~x10 && ~x15 )
						begin
							y12 = 1'b1;	
							nx_state = s290;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && ~x14 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && ~x14 && ~x2 && x15 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && ~x14 && ~x2 && x15 && ~x3 && x10 )
						begin
							y12 = 1'b1;	
							nx_state = s291;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && ~x14 && ~x2 && x15 && ~x3 && ~x10 )
						begin
							y12 = 1'b1;	
							nx_state = s292;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && ~x14 && ~x2 && ~x15 && x10 && x3 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	
							nx_state = s221;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && ~x14 && ~x2 && ~x15 && x10 && ~x3 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && ~x14 && ~x2 && ~x15 && ~x10 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && x16 && ~x17 && ~x14 && ~x2 && ~x15 && ~x10 && ~x3 )
						begin
							y14 = 1'b1;	y16 = 1'b1;	
							nx_state = s216;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && x10 && x15 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && x10 && x15 && ~x3 )
						begin
							y12 = 1'b1;	
							nx_state = s290;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && x10 && ~x15 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && x15 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && x15 && ~x3 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && x13 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && x13 && ~x3 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && ~x13 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && ~x13 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && ~x13 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && ~x13 && ~x4 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && x12 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && x12 && ~x3 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && ~x12 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && ~x12 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && ~x12 && ~x4 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && x11 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && x11 && ~x3 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && ~x11 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && ~x11 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && ~x11 && ~x4 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && ~x17 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && ~x17 && ~x3 && x10 )
						begin
							y12 = 1'b1;	
							nx_state = s293;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && x68 && ~x16 && ~x2 && ~x17 && ~x3 && ~x10 )
						begin
							y12 = 1'b1;	
							nx_state = s231;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && ~x68 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && ~x68 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && ~x68 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && ~x68 && x23 && ~x19 )
						nx_state = s1;
					else if( x66 && ~x67 && ~x65 && ~x21 && ~x22 && ~x68 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x66 && x65 && x15 && x9 && x21 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x66 && x65 && x15 && x9 && ~x21 && x23 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x66 && x65 && x15 && x9 && ~x21 && ~x23 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s294;
						end
					else if( ~x66 && x65 && x15 && ~x9 && x21 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x66 && x65 && x15 && ~x9 && ~x21 && x23 && x6 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x66 && x65 && x15 && ~x9 && ~x21 && x23 && ~x6 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x66 && x65 && x15 && ~x9 && ~x21 && ~x23 && x6 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x66 && x65 && x15 && ~x9 && ~x21 && ~x23 && ~x6 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s294;
						end
					else if( ~x66 && x65 && ~x15 && x21 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && x23 && x9 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && x23 && ~x9 && x12 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && x23 && ~x9 && ~x12 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && x23 && ~x9 && ~x12 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && x23 && ~x9 && ~x12 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && x23 && ~x9 && ~x12 && ~x20 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && ~x23 && x9 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s294;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && ~x23 && ~x9 && x12 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s294;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && ~x23 && ~x9 && ~x12 && x18 && x14 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && ~x23 && ~x9 && ~x12 && x18 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && ~x23 && ~x9 && ~x12 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && x8 && ~x23 && ~x9 && ~x12 && ~x18 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && x23 && x9 && x10 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && x23 && x9 && ~x10 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && x23 && x9 && ~x10 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && x23 && x9 && ~x10 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && x23 && x9 && ~x10 && ~x20 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && x23 && ~x9 && x11 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && x23 && ~x9 && ~x11 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && x23 && ~x9 && ~x11 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && x23 && ~x9 && ~x11 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && x23 && ~x9 && ~x11 && ~x20 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && ~x23 && x9 && x10 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s294;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && ~x23 && x9 && ~x10 && x18 && x14 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && ~x23 && x9 && ~x10 && x18 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && ~x23 && x9 && ~x10 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && ~x23 && x9 && ~x10 && ~x18 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && ~x23 && ~x9 && x11 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s294;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && ~x23 && ~x9 && ~x11 && x18 && x14 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && ~x23 && ~x9 && ~x11 && x18 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && ~x23 && ~x9 && ~x11 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x15 && ~x21 && x16 && ~x8 && ~x23 && ~x9 && ~x11 && ~x18 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x15 && ~x21 && ~x16 && x23 && x6 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && ~x16 && x23 && ~x6 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && ~x16 && ~x23 && x6 )
						begin
							y31 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x66 && x65 && ~x15 && ~x21 && ~x16 && ~x23 && ~x6 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s294;
						end
					else if( ~x66 && ~x65 && x24 && x26 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x66 && ~x65 && x24 && x26 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x66 && ~x65 && x24 && x26 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x24 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x24 && ~x26 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x66 && ~x65 && ~x24 && x25 && x26 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x66 && ~x65 && ~x24 && x25 && x26 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x66 && ~x65 && ~x24 && x25 && x26 && x19 && ~x14 && ~x13 )
						nx_state = s53;
					else if( ~x66 && ~x65 && ~x24 && x25 && x26 && ~x19 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x24 && x25 && ~x26 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s189;
						end
					else if( ~x66 && ~x65 && ~x24 && ~x25 && x26 && x16 && x10 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && ~x65 && ~x24 && ~x25 && x26 && x16 && ~x10 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && ~x65 && ~x24 && ~x25 && x26 && x16 && ~x10 && ~x11 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && ~x65 && ~x24 && ~x25 && x26 && x16 && ~x10 && ~x11 && ~x12 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x66 && ~x65 && ~x24 && ~x25 && x26 && ~x16 && x17 && x10 && x12 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s282;
						end
					else if( ~x66 && ~x65 && ~x24 && ~x25 && x26 && ~x16 && x17 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x66 && ~x65 && ~x24 && ~x25 && x26 && ~x16 && x17 && ~x10 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s282;
						end
					else if( ~x66 && ~x65 && ~x24 && ~x25 && x26 && ~x16 && ~x17 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && ~x65 && ~x24 && ~x25 && ~x26 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else nx_state = s53;
				s54 : if( x65 && x21 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s139;
						end
					else if( x65 && ~x21 && x22 && x23 && x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x15 && x19 && x18 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x15 && x19 && ~x18 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s295;
						end
					else if( x65 && ~x21 && x22 && x23 && ~x15 && ~x19 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( x65 && ~x21 && x22 && ~x23 && x11 && x18 && x15 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x65 && ~x21 && x22 && ~x23 && x11 && x18 && ~x15 )
						begin
							y15 = 1'b1;	y20 = 1'b1;	
							nx_state = s227;
						end
					else if( x65 && ~x21 && x22 && ~x23 && x11 && ~x18 && x19 && x15 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s247;
						end
					else if( x65 && ~x21 && x22 && ~x23 && x11 && ~x18 && x19 && ~x15 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x65 && ~x21 && x22 && ~x23 && x11 && ~x18 && ~x19 )
						begin
							y12 = 1'b1;	
							nx_state = s231;
						end
					else if( x65 && ~x21 && x22 && ~x23 && ~x11 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x65 && ~x21 && ~x22 && x23 && x16 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( x65 && ~x21 && ~x22 && x23 && ~x16 && x20 && x19 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( x65 && ~x21 && ~x22 && x23 && ~x16 && x20 && ~x19 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && ~x22 && x23 && ~x16 && x20 && ~x19 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && ~x22 && x23 && ~x16 && x20 && ~x19 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x22 && x23 && ~x16 && x20 && ~x19 && ~x9 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x22 && x23 && ~x16 && ~x20 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x15 && x19 && x18 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x15 && x19 && ~x18 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s295;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x15 && ~x19 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( ~x65 && x24 && x16 && x26 && x11 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s171;
						end
					else if( ~x65 && x24 && x16 && x26 && ~x11 && x7 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && x24 && x16 && x26 && ~x11 && ~x7 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s171;
						end
					else if( ~x65 && x24 && x16 && ~x26 && x6 && x11 && x12 )
						begin
							y11 = 1'b1;	
							nx_state = s296;
						end
					else if( ~x65 && x24 && x16 && ~x26 && x6 && x11 && ~x12 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s297;
						end
					else if( ~x65 && x24 && x16 && ~x26 && x6 && x11 && ~x12 && ~x13 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x65 && x24 && x16 && ~x26 && x6 && ~x11 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && x24 && x16 && ~x26 && ~x6 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x65 && x24 && ~x16 && x26 && x7 && x17 && x13 && x11 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && x24 && ~x16 && x26 && x7 && x17 && x13 && ~x11 && x12 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( ~x65 && x24 && ~x16 && x26 && x7 && x17 && x13 && ~x11 && ~x12 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && x24 && ~x16 && x26 && x7 && x17 && ~x13 && x11 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s183;
						end
					else if( ~x65 && x24 && ~x16 && x26 && x7 && x17 && ~x13 && ~x11 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && x24 && ~x16 && x26 && x7 && ~x17 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x65 && x24 && ~x16 && x26 && ~x7 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s171;
						end
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && x11 && x9 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && x11 && ~x9 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && x11 && ~x9 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && x11 && ~x9 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && x11 && ~x9 && ~x20 )
						nx_state = s1;
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && ~x11 && x7 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && ~x11 && ~x7 && x12 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && ~x11 && ~x7 && ~x12 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && ~x11 && ~x7 && ~x12 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && ~x11 && ~x7 && ~x12 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && x13 && ~x11 && ~x7 && ~x12 && ~x20 )
						nx_state = s1;
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && x11 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && ~x11 && x12 && x10 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && ~x11 && x12 && ~x10 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && ~x11 && x12 && ~x10 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && ~x11 && x12 && ~x10 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && ~x11 && x12 && ~x10 && ~x20 )
						nx_state = s1;
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && ~x11 && ~x12 && x8 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && ~x11 && ~x12 && ~x8 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && ~x11 && ~x12 && ~x8 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && ~x11 && ~x12 && ~x8 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && x24 && ~x16 && ~x26 && x17 && ~x13 && ~x11 && ~x12 && ~x8 && ~x20 )
						nx_state = s1;
					else if( ~x65 && x24 && ~x16 && ~x26 && ~x17 && x6 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x24 && ~x16 && ~x26 && ~x17 && ~x6 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x65 && ~x24 && x25 && x26 && x1 )
						begin
							y8 = 1'b1;	y17 = 1'b1;	y23 = 1'b1;	
							nx_state = s164;
						end
					else if( ~x65 && ~x24 && x25 && x26 && ~x1 && x18 )
						nx_state = s1;
					else if( ~x65 && ~x24 && x25 && x26 && ~x1 && ~x18 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x65 && ~x24 && x25 && ~x26 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( ~x65 && ~x24 && x25 && ~x26 && ~x2 && x18 && x15 && x10 && x11 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s187;
						end
					else if( ~x65 && ~x24 && x25 && ~x26 && ~x2 && x18 && x15 && x10 && ~x11 && x12 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x65 && ~x24 && x25 && ~x26 && ~x2 && x18 && x15 && x10 && ~x11 && ~x12 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x65 && ~x24 && x25 && ~x26 && ~x2 && x18 && x15 && ~x10 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && ~x24 && x25 && ~x26 && ~x2 && x18 && ~x15 && x16 && x10 && x12 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x65 && ~x24 && x25 && ~x26 && ~x2 && x18 && ~x15 && x16 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && ~x24 && x25 && ~x26 && ~x2 && x18 && ~x15 && x16 && ~x10 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x65 && ~x24 && x25 && ~x26 && ~x2 && x18 && ~x15 && ~x16 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x65 && ~x24 && x25 && ~x26 && ~x2 && ~x18 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x65 && ~x24 && ~x25 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else nx_state = s54;
				s55 : if( x65 && x21 )
						nx_state = s1;
					else if( x65 && ~x21 && x22 && x23 )
						nx_state = s1;
					else if( x65 && ~x21 && x22 && ~x23 && x15 && x9 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x21 && x22 && ~x23 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x65 && ~x21 && x22 && ~x23 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && x22 && ~x23 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s205;
						end
					else if( x65 && ~x21 && ~x22 && x23 && x17 && x15 && x9 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( x65 && ~x21 && ~x22 && x23 && x17 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x65 && ~x21 && ~x22 && x23 && x17 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && ~x22 && x23 && x17 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s205;
						end
					else if( x65 && ~x21 && ~x22 && x23 && ~x17 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( ~x65 && x66 && x63 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x63 && x62 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x63 && ~x62 )
						begin
							y21 = 1'b1;	
							nx_state = s298;
						end
					else if( ~x65 && ~x66 && x25 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	y24 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x65 && ~x66 && ~x25 )
						nx_state = s1;
					else nx_state = s55;
				s56 : if( x66 && x65 && x67 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && x65 && x67 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && x65 && x67 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x66 && x65 && x67 && x22 && ~x17 )
						nx_state = s1;
					else if( x66 && x65 && x67 && ~x22 && x18 && x13 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x66 && x65 && x67 && ~x22 && x18 && x13 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && x67 && ~x22 && x18 && ~x13 && x12 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x66 && x65 && x67 && ~x22 && x18 && ~x13 && x12 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && x67 && ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x66 && x65 && x67 && ~x22 && ~x18 )
						nx_state = s1;
					else if( x66 && x65 && ~x67 && x21 && x20 )
						nx_state = s1;
					else if( x66 && x65 && ~x67 && x21 && ~x20 && x3 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && x18 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y21 = 1'b1;	
							nx_state = s299;
						end
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && x15 && x10 && x11 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s192;
						end
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s193;
						end
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && x15 && x10 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y13 = 1'b1;	
							nx_state = s192;
						end
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s300;
						end
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s192;
						end
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && x10 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && x10 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && x10 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && x10 && ~x19 )
						nx_state = s1;
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && ~x10 && x12 && x11 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s199;
						end
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && ~x10 && x12 && ~x11 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && ~x10 && x12 && ~x11 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && ~x10 && x12 && ~x11 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && ~x10 && x12 && ~x11 && ~x19 )
						nx_state = s1;
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && ~x10 && ~x12 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && ~x10 && ~x12 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && ~x10 && ~x12 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && x16 && ~x10 && ~x12 && ~x19 )
						nx_state = s1;
					else if( x66 && x65 && ~x67 && x21 && ~x20 && ~x3 && ~x18 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s201;
						end
					else if( x66 && x65 && ~x67 && ~x21 && x15 && x10 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x66 && x65 && ~x67 && ~x21 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s301;
						end
					else if( x66 && x65 && ~x67 && ~x21 && x15 && x10 && ~x11 && ~x12 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s195;
						end
					else if( x66 && x65 && ~x67 && ~x21 && x15 && ~x10 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( x66 && x65 && ~x67 && ~x21 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s192;
						end
					else if( x66 && x65 && ~x67 && ~x21 && ~x15 && x16 && x10 && x12 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s259;
						end
					else if( x66 && x65 && ~x67 && ~x21 && ~x15 && x16 && x10 && ~x12 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s302;
						end
					else if( x66 && x65 && ~x67 && ~x21 && ~x15 && x16 && ~x10 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s259;
						end
					else if( x66 && x65 && ~x67 && ~x21 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s303;
						end
					else if( x66 && ~x65 && x21 && x15 && x4 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x66 && ~x65 && x21 && x15 && x4 && ~x10 && x12 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x66 && ~x65 && x21 && x15 && x4 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( x66 && ~x65 && x21 && x15 && ~x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( x66 && ~x65 && x21 && ~x15 && x16 && x10 && x12 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( x66 && ~x65 && x21 && ~x15 && x16 && x10 && ~x12 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s304;
						end
					else if( x66 && ~x65 && x21 && ~x15 && x16 && ~x10 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( x66 && ~x65 && x21 && ~x15 && ~x16 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( x66 && ~x65 && x21 && ~x15 && ~x16 && ~x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( x66 && ~x65 && ~x21 && x22 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( x66 && ~x65 && ~x21 && ~x22 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s250;
						end
					else if( x66 && ~x65 && ~x21 && ~x22 && ~x23 )
						begin
							y2 = 1'b1;	
							nx_state = s85;
						end
					else if( ~x66 && x65 && x68 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x66 && x65 && x68 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x66 && x65 && x68 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x66 && x65 && x68 && ~x5 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x68 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x66 && x65 && ~x68 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && ~x68 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && ~x68 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x68 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && x7 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && x7 && ~x9 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && x8 && x9 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && x8 && ~x9 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && ~x8 && x9 && x13 )
						begin
							y4 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && ~x8 && x9 && ~x13 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && ~x8 && x9 && ~x13 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && ~x8 && x9 && ~x13 && ~x19 && x17 && ~x14 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && ~x8 && x9 && ~x13 && ~x19 && ~x17 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && ~x8 && ~x9 && x14 )
						begin
							y4 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && ~x8 && ~x9 && ~x14 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && ~x8 && ~x9 && ~x14 && ~x19 && x17 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && ~x8 && ~x9 && ~x14 && ~x19 && x17 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && x16 && ~x7 && ~x8 && ~x9 && ~x14 && ~x19 && ~x17 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && ~x16 && x7 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && ~x16 && ~x7 && x8 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && ~x16 && ~x7 && ~x8 && x4 )
						begin
							y1 = 1'b1;	
							nx_state = s22;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && ~x16 && ~x7 && ~x8 && ~x4 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && ~x16 && ~x7 && ~x8 && ~x4 && ~x5 && x9 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && x15 && ~x16 && ~x7 && ~x8 && ~x4 && ~x5 && ~x9 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && x4 )
						begin
							y1 = 1'b1;	
							nx_state = s22;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && x9 && ~x10 && x8 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && x9 && ~x10 && ~x8 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && x9 && ~x10 && ~x8 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && x9 && ~x10 && ~x8 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && x9 && ~x10 && ~x8 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && x9 && ~x10 && ~x8 && ~x19 && ~x17 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && x8 && x12 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && x8 && ~x12 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && x8 && ~x12 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && x8 && ~x12 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && x8 && ~x12 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && x8 && ~x12 && ~x19 && ~x17 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && ~x8 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && ~x8 && ~x11 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && ~x8 && ~x11 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && ~x8 && ~x11 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && ~x8 && ~x11 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && x16 && ~x9 && ~x8 && ~x11 && ~x19 && ~x17 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && ~x16 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && x22 && ~x15 && ~x4 && ~x16 && ~x5 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s212;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && ~x22 && x2 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x2 && x17 && x15 && x9 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x2 && x17 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x2 && x17 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x2 && x17 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x66 && x65 && ~x68 && ~x21 && ~x22 && ~x2 && ~x17 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( ~x66 && ~x65 && x20 && x15 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x66 && ~x65 && x20 && ~x15 )
						begin
							y7 = 1'b1;	y12 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x66 && ~x65 && ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x66 && ~x65 && ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x66 && ~x65 && ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x66 && ~x65 && ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x66 && ~x65 && ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else nx_state = s56;
				s57 : if( x21 )
						nx_state = s1;
					else if( ~x21 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else nx_state = s57;
				s58 : if( x68 && x21 && x20 )
						begin
							y4 = 1'b1;	
							nx_state = s191;
						end
					else if( x68 && x21 && ~x20 )
						nx_state = s1;
					else if( x68 && ~x21 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x68 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else nx_state = s58;
				s59 : if( x65 && x21 )
						nx_state = s1;
					else if( x65 && ~x21 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s60;
						end
					else if( ~x65 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x20 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x65 && ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x65 && ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else nx_state = s59;
				s60 : if( x21 && x20 && x2 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s306;
						end
					else if( x21 && x20 && ~x2 && x18 && x15 && x10 && x11 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s192;
						end
					else if( x21 && x20 && ~x2 && x18 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s193;
						end
					else if( x21 && x20 && ~x2 && x18 && x15 && x10 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s194;
						end
					else if( x21 && x20 && ~x2 && x18 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s300;
						end
					else if( x21 && x20 && ~x2 && x18 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s192;
						end
					else if( x21 && x20 && ~x2 && x18 && ~x15 && x16 && x10 && x12 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s259;
						end
					else if( x21 && x20 && ~x2 && x18 && ~x15 && x16 && x10 && ~x12 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( x21 && x20 && ~x2 && x18 && ~x15 && x16 && ~x10 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s259;
						end
					else if( x21 && x20 && ~x2 && x18 && ~x15 && ~x16 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x21 && x20 && ~x2 && ~x18 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	
							nx_state = s307;
						end
					else if( x21 && ~x20 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	
							nx_state = s307;
						end
					else if( ~x21 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	
							nx_state = s307;
						end
					else nx_state = s60;
				s61 : if( x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( ~x21 )
						nx_state = s1;
					else nx_state = s61;
				s62 : if( x65 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( ~x65 && x66 && x21 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s232;
						end
					else if( ~x65 && x66 && ~x21 && x22 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s262;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && x10 && x16 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s219;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && x10 && ~x16 && x17 && x15 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s219;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && x10 && ~x16 && x17 && ~x15 && x3 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s214;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && x10 && ~x16 && x17 && ~x15 && ~x3 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s308;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && x10 && ~x16 && ~x17 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s219;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && ~x10 && x16 && x15 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s309;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && ~x10 && x16 && ~x15 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s310;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && ~x10 && ~x16 && x17 && x15 && x14 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && ~x10 && ~x16 && x17 && x15 && ~x14 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s79;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && ~x10 && ~x16 && x17 && ~x15 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s79;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && ~x10 && ~x16 && ~x17 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s311;
						end
					else if( ~x65 && ~x66 && x68 && x21 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x66 && x68 && ~x21 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x65 && ~x66 && ~x68 && x22 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && ~x66 && ~x68 && ~x22 && x21 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && ~x66 && ~x68 && ~x22 && ~x21 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else nx_state = s62;
				s63 : if( x61 && x60 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x61 && ~x60 && x62 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x61 && ~x60 && ~x62 )
						nx_state = s40;
					else if( ~x61 && x60 )
						nx_state = s40;
					else if( ~x61 && ~x60 && x62 )
						nx_state = s40;
					else if( ~x61 && ~x60 && ~x62 )
						nx_state = s1;
					else nx_state = s63;
				s64 : if( x60 && x61 )
						begin
							y14 = 1'b1;	
							nx_state = s286;
						end
					else if( x60 && ~x61 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x60 && x62 && x61 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x60 && x62 && x61 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x60 && x62 && x61 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( ~x60 && x62 && x61 && ~x18 )
						nx_state = s1;
					else if( ~x60 && x62 && ~x61 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s312;
						end
					else if( ~x60 && ~x62 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s154;
						end
					else nx_state = s64;
				s65 : if( x65 && x66 && x61 && x60 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( x65 && x66 && x61 && ~x60 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s258;
						end
					else if( x65 && x66 && ~x61 && x60 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s258;
						end
					else if( x65 && x66 && ~x61 && ~x60 )
						nx_state = s40;
					else if( x65 && ~x66 )
						begin
							y15 = 1'b1;	y21 = 1'b1;	y28 = 1'b1;	
							nx_state = s313;
						end
					else if( ~x65 && x66 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && ~x66 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && x19 && ~x14 && ~x13 )
						nx_state = s65;
					else if( ~x65 && ~x66 && ~x19 )
						nx_state = s1;
					else nx_state = s65;
				s66 : if( x61 && x60 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s68;
						end
					else if( x61 && ~x60 && x62 )
						nx_state = s1;
					else if( x61 && ~x60 && ~x62 )
						nx_state = s39;
					else if( ~x61 && x60 )
						nx_state = s39;
					else if( ~x61 && ~x60 && x62 && x4 && x15 && x12 && x7 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s314;
						end
					else if( ~x61 && ~x60 && x62 && x4 && x15 && x12 && ~x7 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s315;
						end
					else if( ~x61 && ~x60 && x62 && x4 && x15 && ~x12 && x7 )
						nx_state = s316;
					else if( ~x61 && ~x60 && x62 && x4 && x15 && ~x12 && ~x7 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x61 && ~x60 && x62 && x4 && ~x15 && x16 && x7 && x12 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s315;
						end
					else if( ~x61 && ~x60 && x62 && x4 && ~x15 && x16 && x7 && ~x12 )
						nx_state = s316;
					else if( ~x61 && ~x60 && x62 && x4 && ~x15 && x16 && ~x7 )
						nx_state = s316;
					else if( ~x61 && ~x60 && x62 && x4 && ~x15 && ~x16 && x7 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x61 && ~x60 && x62 && x4 && ~x15 && ~x16 && ~x7 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x61 && ~x60 && x62 && ~x4 )
						nx_state = s316;
					else if( ~x61 && ~x60 && ~x62 && x15 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x61 && ~x60 && ~x62 && x15 && ~x7 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x61 && ~x60 && ~x62 && x15 && ~x7 && ~x11 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x61 && ~x60 && ~x62 && ~x15 && x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x61 && ~x60 && ~x62 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else nx_state = s66;
				s67 : if( x65 && x60 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s68;
						end
					else if( x65 && ~x60 && x61 )
						nx_state = s1;
					else if( x65 && ~x60 && ~x61 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s118;
						end
					else if( ~x65 && x21 && x3 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	
							nx_state = s141;
						end
					else if( ~x65 && x21 && ~x3 && x20 && x16 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s113;
						end
					else if( ~x65 && x21 && ~x3 && x20 && x16 && ~x10 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && x21 && ~x3 && x20 && ~x16 && x17 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x65 && x21 && ~x3 && x20 && ~x16 && ~x17 )
						begin
							y5 = 1'b1;	y17 = 1'b1;	
							nx_state = s115;
						end
					else if( ~x65 && x21 && ~x3 && ~x20 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s317;
						end
					else if( ~x65 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x65 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x65 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x21 && ~x20 )
						nx_state = s1;
					else nx_state = s67;
				s68 : if( x60 && x61 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x60 && x61 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x60 && x61 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x60 && x61 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x60 && ~x61 && x15 && x5 && x12 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s318;
						end
					else if( x60 && ~x61 && x15 && x5 && x12 && ~x7 )
						begin
							y4 = 1'b1;	
							nx_state = s318;
						end
					else if( x60 && ~x61 && x15 && x5 && ~x12 && x7 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( x60 && ~x61 && x15 && x5 && ~x12 && ~x7 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s254;
						end
					else if( x60 && ~x61 && x15 && ~x5 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( x60 && ~x61 && ~x15 && x16 && x7 && x12 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s75;
						end
					else if( x60 && ~x61 && ~x15 && x16 && x7 && x12 && ~x5 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( x60 && ~x61 && ~x15 && x16 && x7 && ~x12 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( x60 && ~x61 && ~x15 && x16 && ~x7 && x12 && x9 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( x60 && ~x61 && ~x15 && x16 && ~x7 && x12 && ~x9 && x11 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( x60 && ~x61 && ~x15 && x16 && ~x7 && x12 && ~x9 && ~x11 )
						nx_state = s1;
					else if( x60 && ~x61 && ~x15 && x16 && ~x7 && ~x12 && x11 && x10 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( x60 && ~x61 && ~x15 && x16 && ~x7 && ~x12 && x11 && ~x10 )
						nx_state = s1;
					else if( x60 && ~x61 && ~x15 && x16 && ~x7 && ~x12 && ~x11 && x8 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( x60 && ~x61 && ~x15 && x16 && ~x7 && ~x12 && ~x11 && ~x8 )
						nx_state = s1;
					else if( x60 && ~x61 && ~x15 && ~x16 && x5 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s253;
						end
					else if( x60 && ~x61 && ~x15 && ~x16 && x5 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x60 && ~x61 && ~x15 && ~x16 && ~x5 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( ~x60 && x61 && x62 )
						begin
							y14 = 1'b1;	
							nx_state = s286;
						end
					else if( ~x60 && x61 && ~x62 && x15 && x5 && x12 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s318;
						end
					else if( ~x60 && x61 && ~x62 && x15 && x5 && x12 && ~x7 )
						begin
							y4 = 1'b1;	
							nx_state = s318;
						end
					else if( ~x60 && x61 && ~x62 && x15 && x5 && ~x12 && x7 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( ~x60 && x61 && ~x62 && x15 && x5 && ~x12 && ~x7 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x60 && x61 && ~x62 && x15 && ~x5 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( ~x60 && x61 && ~x62 && ~x15 && x16 && x7 && x12 && x5 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x60 && x61 && ~x62 && ~x15 && x16 && x7 && x12 && ~x5 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( ~x60 && x61 && ~x62 && ~x15 && x16 && x7 && ~x12 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( ~x60 && x61 && ~x62 && ~x15 && x16 && ~x7 && x12 && x9 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( ~x60 && x61 && ~x62 && ~x15 && x16 && ~x7 && x12 && ~x9 && x11 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( ~x60 && x61 && ~x62 && ~x15 && x16 && ~x7 && x12 && ~x9 && ~x11 )
						nx_state = s1;
					else if( ~x60 && x61 && ~x62 && ~x15 && x16 && ~x7 && ~x12 && x11 && x10 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( ~x60 && x61 && ~x62 && ~x15 && x16 && ~x7 && ~x12 && x11 && ~x10 )
						nx_state = s1;
					else if( ~x60 && x61 && ~x62 && ~x15 && x16 && ~x7 && ~x12 && ~x11 && x8 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( ~x60 && x61 && ~x62 && ~x15 && x16 && ~x7 && ~x12 && ~x11 && ~x8 )
						nx_state = s1;
					else if( ~x60 && x61 && ~x62 && ~x15 && ~x16 && x5 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s253;
						end
					else if( ~x60 && x61 && ~x62 && ~x15 && ~x16 && x5 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x60 && x61 && ~x62 && ~x15 && ~x16 && ~x5 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( ~x60 && ~x61 && x62 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x60 && ~x61 && ~x62 )
						begin
							y3 = 1'b1;	
							nx_state = s320;
						end
					else nx_state = s68;
				s69 : if( x65 && x60 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s68;
						end
					else if( x65 && ~x60 && x61 )
						begin
							y2 = 1'b1;	y19 = 1'b1;	y24 = 1'b1;	
							nx_state = s321;
						end
					else if( x65 && ~x60 && ~x61 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( ~x65 )
						begin
							y14 = 1'b1;	
							nx_state = s286;
						end
					else nx_state = s69;
				s70 : if( x60 )
						nx_state = s316;
					else if( ~x60 && x61 )
						nx_state = s316;
					else if( ~x60 && ~x61 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else nx_state = s70;
				s71 : if( x60 )
						nx_state = s316;
					else if( ~x60 && x61 )
						nx_state = s316;
					else if( ~x60 && ~x61 && x17 && x62 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s255;
						end
					else if( ~x60 && ~x61 && x17 && ~x62 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x60 && ~x61 && ~x17 )
						nx_state = s39;
					else nx_state = s71;
				s72 : if( x65 && x66 && x61 && x60 )
						nx_state = s1;
					else if( x65 && x66 && x61 && ~x60 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x66 && x61 && ~x60 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x66 && x61 && ~x60 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x65 && x66 && x61 && ~x60 && x62 && ~x18 )
						nx_state = s1;
					else if( x65 && x66 && x61 && ~x60 && ~x62 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( x65 && x66 && ~x61 && x60 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( x65 && x66 && ~x61 && ~x60 && x62 && x7 && x15 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s292;
						end
					else if( x65 && x66 && ~x61 && ~x60 && x62 && x7 && x15 && ~x12 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s63;
						end
					else if( x65 && x66 && ~x61 && ~x60 && x62 && x7 && ~x15 && x16 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s290;
						end
					else if( x65 && x66 && ~x61 && ~x60 && x62 && x7 && ~x15 && x16 && ~x12 && x2 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s322;
						end
					else if( x65 && x66 && ~x61 && ~x60 && x62 && x7 && ~x15 && x16 && ~x12 && ~x2 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s262;
						end
					else if( x65 && x66 && ~x61 && ~x60 && x62 && x7 && ~x15 && ~x16 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && x66 && ~x61 && ~x60 && x62 && ~x7 && x15 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s290;
						end
					else if( x65 && x66 && ~x61 && ~x60 && x62 && ~x7 && x15 && ~x12 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s263;
						end
					else if( x65 && x66 && ~x61 && ~x60 && x62 && ~x7 && ~x15 && x16 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x65 && x66 && ~x61 && ~x60 && x62 && ~x7 && ~x15 && ~x16 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x66 && ~x61 && ~x60 && ~x62 && x4 && x15 && x7 )
						nx_state = s40;
					else if( x65 && x66 && ~x61 && ~x60 && ~x62 && x4 && x15 && ~x7 && x11 )
						nx_state = s40;
					else if( x65 && x66 && ~x61 && ~x60 && ~x62 && x4 && x15 && ~x7 && ~x11 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x66 && ~x61 && ~x60 && ~x62 && x4 && ~x15 && x16 )
						nx_state = s70;
					else if( x65 && x66 && ~x61 && ~x60 && ~x62 && x4 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( x65 && x66 && ~x61 && ~x60 && ~x62 && ~x4 )
						nx_state = s70;
					else if( x65 && ~x66 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( ~x65 && x21 && x66 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x21 && x66 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x21 && x66 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && x21 && x66 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x21 && ~x66 && x19 && x20 && x12 && x17 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	
							nx_state = s266;
						end
					else if( ~x65 && x21 && ~x66 && x19 && x20 && x12 && ~x17 )
						begin
							y8 = 1'b1;	y22 = 1'b1;	
							nx_state = s267;
						end
					else if( ~x65 && x21 && ~x66 && x19 && x20 && ~x12 && x16 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x65 && x21 && ~x66 && x19 && x20 && ~x12 && ~x16 && x17 && x5 )
						begin
							y8 = 1'b1;	
							nx_state = s181;
						end
					else if( ~x65 && x21 && ~x66 && x19 && x20 && ~x12 && ~x16 && x17 && ~x5 )
						begin
							y8 = 1'b1;	
							nx_state = s246;
						end
					else if( ~x65 && x21 && ~x66 && x19 && x20 && ~x12 && ~x16 && ~x17 && x4 )
						begin
							y8 = 1'b1;	
							nx_state = s181;
						end
					else if( ~x65 && x21 && ~x66 && x19 && x20 && ~x12 && ~x16 && ~x17 && ~x4 )
						begin
							y8 = 1'b1;	
							nx_state = s246;
						end
					else if( ~x65 && x21 && ~x66 && x19 && ~x20 && x16 && x12 )
						begin
							y8 = 1'b1;	y18 = 1'b1;	
							nx_state = s323;
						end
					else if( ~x65 && x21 && ~x66 && x19 && ~x20 && x16 && ~x12 && x17 )
						begin
							y8 = 1'b1;	y18 = 1'b1;	
							nx_state = s82;
						end
					else if( ~x65 && x21 && ~x66 && x19 && ~x20 && x16 && ~x12 && ~x17 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x65 && x21 && ~x66 && x19 && ~x20 && ~x16 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x65 && x21 && ~x66 && ~x19 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x65 && ~x21 && x66 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x21 && ~x66 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else nx_state = s72;
				s73 : if( x60 && x15 && x12 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x60 && x15 && x12 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s250;
						end
					else if( x60 && x15 && ~x12 && x7 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x60 && x15 && ~x12 && ~x7 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s262;
						end
					else if( x60 && ~x15 && x16 && x7 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s251;
						end
					else if( x60 && ~x15 && x16 && x7 && ~x12 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x60 && ~x15 && x16 && ~x7 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x60 && ~x15 && ~x16 && x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s318;
						end
					else if( x60 && ~x15 && ~x16 && ~x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s74;
						end
					else if( ~x60 && x61 && x15 && x12 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x60 && x61 && x15 && x12 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s250;
						end
					else if( ~x60 && x61 && x15 && ~x12 && x7 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x60 && x61 && x15 && ~x12 && ~x7 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s262;
						end
					else if( ~x60 && x61 && ~x15 && x16 && x7 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s251;
						end
					else if( ~x60 && x61 && ~x15 && x16 && x7 && ~x12 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x60 && x61 && ~x15 && x16 && ~x7 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x60 && x61 && ~x15 && ~x16 && x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s318;
						end
					else if( ~x60 && x61 && ~x15 && ~x16 && ~x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s74;
						end
					else if( ~x60 && ~x61 && x62 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y24 = 1'b1;	
							nx_state = s64;
						end
					else if( ~x60 && ~x61 && ~x62 )
						begin
							y25 = 1'b1;	
							nx_state = s324;
						end
					else nx_state = s73;
				s74 : if( x61 && x60 && x7 && x15 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x61 && x60 && x7 && ~x15 && x16 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s251;
						end
					else if( x61 && x60 && x7 && ~x15 && x16 && ~x12 && x3 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s258;
						end
					else if( x61 && x60 && x7 && ~x15 && x16 && ~x12 && ~x3 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( x61 && x60 && x7 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s253;
						end
					else if( x61 && x60 && ~x7 && x15 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s250;
						end
					else if( x61 && x60 && ~x7 && x15 && ~x12 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( x61 && x60 && ~x7 && ~x15 && x16 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x61 && x60 && ~x7 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x61 && ~x60 && x62 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x61 && ~x60 && ~x62 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x61 && x60 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x61 && ~x60 && x62 && x16 && x15 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x61 && ~x60 && x62 && x16 && ~x15 && x11 && x12 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x61 && ~x60 && x62 && x16 && ~x15 && x11 && ~x12 && x7 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x61 && ~x60 && x62 && x16 && ~x15 && x11 && ~x12 && ~x7 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x61 && ~x60 && x62 && x16 && ~x15 && ~x11 && x7 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x61 && ~x60 && x62 && x16 && ~x15 && ~x11 && ~x7 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x61 && ~x60 && x62 && ~x16 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x61 && ~x60 && ~x62 && x15 && x16 && x9 && x11 )
						nx_state = s40;
					else if( ~x61 && ~x60 && ~x62 && x15 && x16 && x9 && ~x11 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x61 && ~x60 && ~x62 && x15 && x16 && x9 && ~x11 && ~x7 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s261;
						end
					else if( ~x61 && ~x60 && ~x62 && x15 && x16 && ~x9 && x11 && x7 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s262;
						end
					else if( ~x61 && ~x60 && ~x62 && x15 && x16 && ~x9 && x11 && ~x7 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s260;
						end
					else if( ~x61 && ~x60 && ~x62 && x15 && x16 && ~x9 && ~x11 && x7 && x14 )
						nx_state = s316;
					else if( ~x61 && ~x60 && ~x62 && x15 && x16 && ~x9 && ~x11 && x7 && ~x14 )
						nx_state = s40;
					else if( ~x61 && ~x60 && ~x62 && x15 && x16 && ~x9 && ~x11 && ~x7 && x13 )
						nx_state = s316;
					else if( ~x61 && ~x60 && ~x62 && x15 && x16 && ~x9 && ~x11 && ~x7 && ~x13 )
						nx_state = s40;
					else if( ~x61 && ~x60 && ~x62 && x15 && ~x16 && x9 && x3 )
						nx_state = s40;
					else if( ~x61 && ~x60 && ~x62 && x15 && ~x16 && x9 && ~x3 && x7 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s325;
						end
					else if( ~x61 && ~x60 && ~x62 && x15 && ~x16 && x9 && ~x3 && ~x7 && x11 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s325;
						end
					else if( ~x61 && ~x60 && ~x62 && x15 && ~x16 && x9 && ~x3 && ~x7 && ~x11 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x61 && ~x60 && ~x62 && x15 && ~x16 && ~x9 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s69;
						end
					else if( ~x61 && ~x60 && ~x62 && x15 && ~x16 && ~x9 && ~x3 && x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x61 && ~x60 && ~x62 && x15 && ~x16 && ~x9 && ~x3 && ~x5 && x7 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s326;
						end
					else if( ~x61 && ~x60 && ~x62 && x15 && ~x16 && ~x9 && ~x3 && ~x5 && ~x7 && x11 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x61 && ~x60 && ~x62 && x15 && ~x16 && ~x9 && ~x3 && ~x5 && ~x7 && ~x11 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x61 && ~x60 && ~x62 && ~x15 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s69;
						end
					else if( ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && x11 && x9 )
						nx_state = s40;
					else if( ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && x11 && ~x9 && x7 && x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && x11 && ~x9 && x7 && ~x5 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s326;
						end
					else if( ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && x11 && ~x9 && ~x7 && x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s131;
						end
					else if( ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && x11 && ~x9 && ~x7 && ~x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s67;
						end
					else if( ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && x7 && x9 && x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s256;
						end
					else if( ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && x7 && x9 && ~x5 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && x7 && ~x9 && x8 && x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s256;
						end
					else if( ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && x7 && ~x9 && x8 && ~x5 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && x7 && ~x9 && ~x8 )
						nx_state = s40;
					else if( ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && ~x7 && x9 && x10 && x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s256;
						end
					else if( ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && ~x7 && x9 && x10 && ~x5 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && ~x7 && x9 && ~x10 )
						nx_state = s40;
					else if( ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && ~x7 && ~x9 && x12 && x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s256;
						end
					else if( ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && ~x7 && ~x9 && x12 && ~x5 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s252;
						end
					else if( ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && x16 && ~x11 && ~x7 && ~x9 && ~x12 )
						nx_state = s40;
					else if( ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && ~x16 && x5 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x61 && ~x60 && ~x62 && ~x15 && ~x3 && ~x16 && ~x5 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s68;
						end
					else nx_state = s74;
				s75 : if( x65 && x60 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( x65 && ~x60 && x61 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( x65 && ~x60 && ~x61 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x65 && x21 && x16 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s113;
						end
					else if( ~x65 && x21 && x16 && ~x10 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && x21 && ~x16 && x17 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x65 && x21 && ~x16 && ~x17 )
						begin
							y5 = 1'b1;	y17 = 1'b1;	
							nx_state = s115;
						end
					else if( ~x65 && ~x21 && x3 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s14;
						end
					else if( ~x65 && ~x21 && ~x3 && x19 && x16 && x10 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s67;
						end
					else if( ~x65 && ~x21 && ~x3 && x19 && x16 && ~x10 )
						begin
							y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s113;
						end
					else if( ~x65 && ~x21 && ~x3 && x19 && ~x16 && x17 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x65 && ~x21 && ~x3 && x19 && ~x16 && ~x17 )
						begin
							y5 = 1'b1;	y17 = 1'b1;	
							nx_state = s115;
						end
					else if( ~x65 && ~x21 && ~x3 && ~x19 )
						begin
							y13 = 1'b1;	y17 = 1'b1;	
							nx_state = s141;
						end
					else nx_state = s75;
				s76 : if( x65 && x61 && x60 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x61 && x60 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x61 && x60 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x61 && x60 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x61 && ~x60 && x62 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x15 && x16 && x7 && x12 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x15 && x16 && x7 && ~x12 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x15 && x16 && ~x7 && x12 && x14 && x11 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s260;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x15 && x16 && ~x7 && x12 && x14 && ~x11 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x15 && x16 && ~x7 && x12 && ~x14 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x15 && x16 && ~x7 && x12 && ~x14 && x18 && ~x13 )
						nx_state = s39;
					else if( x65 && x61 && ~x60 && ~x62 && x15 && x16 && ~x7 && x12 && ~x14 && ~x18 )
						nx_state = s39;
					else if( x65 && x61 && ~x60 && ~x62 && x15 && x16 && ~x7 && ~x12 && x13 && x11 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s261;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x15 && x16 && ~x7 && ~x12 && x13 && ~x11 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x15 && x16 && ~x7 && ~x12 && ~x13 && x18 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x15 && x16 && ~x7 && ~x12 && ~x13 && x18 && ~x14 )
						nx_state = s39;
					else if( x65 && x61 && ~x60 && ~x62 && x15 && x16 && ~x7 && ~x12 && ~x13 && ~x18 )
						nx_state = s39;
					else if( x65 && x61 && ~x60 && ~x62 && x15 && ~x16 && x11 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s327;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x15 && ~x16 && x11 && ~x7 && x12 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x15 && ~x16 && x11 && ~x7 && ~x12 )
						begin
							y4 = 1'b1;	
							nx_state = s318;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x15 && ~x16 && ~x11 && x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s328;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x15 && ~x16 && ~x11 && ~x4 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x15 && ~x16 && ~x11 && ~x4 && ~x2 && x12 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s329;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x15 && ~x16 && ~x11 && ~x4 && ~x2 && x12 && ~x7 )
						begin
							y4 = 1'b1;	
							nx_state = s318;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x15 && ~x16 && ~x11 && ~x4 && ~x2 && ~x12 && x7 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s263;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x15 && ~x16 && ~x11 && ~x4 && ~x2 && ~x12 && ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x61 && ~x60 && ~x62 && ~x15 && x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s328;
						end
					else if( x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && x7 && x12 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && x7 && x12 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s318;
						end
					else if( x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && x7 && ~x12 )
						begin
							y3 = 1'b1;	
							nx_state = s65;
						end
					else if( x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && x12 && x11 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && x12 && x11 && ~x2 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && x12 && ~x11 && x9 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && x12 && ~x11 && x9 && ~x2 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && x12 && ~x11 && ~x9 )
						nx_state = s1;
					else if( x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && x11 && x10 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && x11 && x10 && ~x2 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && x11 && ~x10 )
						nx_state = s1;
					else if( x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && ~x11 && x8 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && ~x11 && x8 && ~x2 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && ~x11 && ~x8 )
						nx_state = s1;
					else if( x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && ~x16 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && ~x16 && ~x2 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s318;
						end
					else if( x65 && x61 && ~x60 && ~x62 && ~x15 && ~x4 && ~x16 && ~x2 && ~x7 )
						begin
							y4 = 1'b1;	
							nx_state = s191;
						end
					else if( x65 && ~x61 && x60 && x15 && x16 && x7 && x12 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( x65 && ~x61 && x60 && x15 && x16 && x7 && ~x12 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( x65 && ~x61 && x60 && x15 && x16 && ~x7 && x12 && x14 && x11 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s260;
						end
					else if( x65 && ~x61 && x60 && x15 && x16 && ~x7 && x12 && x14 && ~x11 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x65 && ~x61 && x60 && x15 && x16 && ~x7 && x12 && ~x14 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x61 && x60 && x15 && x16 && ~x7 && x12 && ~x14 && x18 && ~x13 )
						nx_state = s39;
					else if( x65 && ~x61 && x60 && x15 && x16 && ~x7 && x12 && ~x14 && ~x18 )
						nx_state = s39;
					else if( x65 && ~x61 && x60 && x15 && x16 && ~x7 && ~x12 && x13 && x11 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s261;
						end
					else if( x65 && ~x61 && x60 && x15 && x16 && ~x7 && ~x12 && x13 && ~x11 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x65 && ~x61 && x60 && x15 && x16 && ~x7 && ~x12 && ~x13 && x18 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x61 && x60 && x15 && x16 && ~x7 && ~x12 && ~x13 && x18 && ~x14 )
						nx_state = s39;
					else if( x65 && ~x61 && x60 && x15 && x16 && ~x7 && ~x12 && ~x13 && ~x18 )
						nx_state = s39;
					else if( x65 && ~x61 && x60 && x15 && ~x16 && x11 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s327;
						end
					else if( x65 && ~x61 && x60 && x15 && ~x16 && x11 && ~x7 && x12 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( x65 && ~x61 && x60 && x15 && ~x16 && x11 && ~x7 && ~x12 )
						begin
							y4 = 1'b1;	
							nx_state = s318;
						end
					else if( x65 && ~x61 && x60 && x15 && ~x16 && ~x11 && x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s328;
						end
					else if( x65 && ~x61 && x60 && x15 && ~x16 && ~x11 && ~x4 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && ~x61 && x60 && x15 && ~x16 && ~x11 && ~x4 && ~x2 && x12 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s329;
						end
					else if( x65 && ~x61 && x60 && x15 && ~x16 && ~x11 && ~x4 && ~x2 && x12 && ~x7 )
						begin
							y4 = 1'b1;	
							nx_state = s318;
						end
					else if( x65 && ~x61 && x60 && x15 && ~x16 && ~x11 && ~x4 && ~x2 && ~x12 && x7 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s263;
						end
					else if( x65 && ~x61 && x60 && x15 && ~x16 && ~x11 && ~x4 && ~x2 && ~x12 && ~x7 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x61 && x60 && ~x15 && x4 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s328;
						end
					else if( x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && x7 && x12 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && x7 && x12 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s318;
						end
					else if( x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && x7 && ~x12 )
						begin
							y3 = 1'b1;	
							nx_state = s65;
						end
					else if( x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && x12 && x11 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && x12 && x11 && ~x2 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && x12 && ~x11 && x9 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && x12 && ~x11 && x9 && ~x2 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && x12 && ~x11 && ~x9 )
						nx_state = s1;
					else if( x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && x11 && x10 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && x11 && x10 && ~x2 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && x11 && ~x10 )
						nx_state = s1;
					else if( x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && ~x11 && x8 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && ~x11 && x8 && ~x2 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && ~x61 && x60 && ~x15 && ~x4 && x16 && ~x7 && ~x12 && ~x11 && ~x8 )
						nx_state = s1;
					else if( x65 && ~x61 && x60 && ~x15 && ~x4 && ~x16 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && ~x61 && x60 && ~x15 && ~x4 && ~x16 && ~x2 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s318;
						end
					else if( x65 && ~x61 && x60 && ~x15 && ~x4 && ~x16 && ~x2 && ~x7 )
						begin
							y4 = 1'b1;	
							nx_state = s191;
						end
					else if( x65 && ~x61 && ~x60 && x62 )
						nx_state = s40;
					else if( x65 && ~x61 && ~x60 && ~x62 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s74;
						end
					else if( ~x65 && x15 && x66 && x21 && x10 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s330;
						end
					else if( ~x65 && x15 && x66 && x21 && ~x10 && x12 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x65 && x15 && x66 && x21 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && x10 && x23 && x16 && x12 )
						begin
							y14 = 1'b1;	
							nx_state = s331;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && x10 && x23 && x16 && ~x12 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && x10 && x23 && ~x16 && x11 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && x10 && x23 && ~x16 && ~x11 && x12 )
						begin
							y14 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && x10 && x23 && ~x16 && ~x11 && ~x12 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && x10 && x23 && ~x16 && ~x11 && ~x12 && ~x2 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && x10 && x23 && ~x16 && ~x11 && ~x12 && ~x2 && ~x4 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s333;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && x10 && ~x23 && x11 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s334;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && x10 && ~x23 && ~x11 && x12 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s334;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && x10 && ~x23 && ~x11 && ~x12 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && x11 && x16 && x12 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s330;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && x11 && x16 && ~x12 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && x11 && ~x16 && x12 )
						begin
							y1 = 1'b1;	
							nx_state = s22;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && x11 && ~x16 && ~x12 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && x16 && x12 && x13 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s335;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && x16 && x12 && ~x13 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && x16 && x12 && ~x13 && x17 && ~x14 )
						nx_state = s1;
					else if( ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && x16 && x12 && ~x13 && ~x17 )
						nx_state = s1;
					else if( ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && x16 && ~x12 && x14 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s335;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && x16 && ~x12 && ~x14 && x17 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && x16 && ~x12 && ~x14 && x17 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && x16 && ~x12 && ~x14 && ~x17 )
						nx_state = s1;
					else if( ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && ~x16 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && ~x16 && ~x2 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && ~x16 && ~x2 && ~x4 && x12 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && x23 && ~x11 && ~x16 && ~x2 && ~x4 && ~x12 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s336;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && ~x23 && x12 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && ~x23 && x12 && ~x11 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x65 && x15 && x66 && ~x21 && x22 && ~x10 && ~x23 && ~x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && x9 && x7 && x23 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && x9 && x7 && ~x23 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && x9 && ~x7 && x8 && x23 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && x9 && ~x7 && x8 && ~x23 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s126;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && x9 && ~x7 && ~x8 && x13 && x23 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s337;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && x9 && ~x7 && ~x8 && x13 && ~x23 )
						begin
							y7 = 1'b1;	
							nx_state = s338;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && x9 && ~x7 && ~x8 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && ~x9 && x7 && x23 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && ~x9 && x7 && ~x23 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && ~x9 && ~x7 && x8 && x23 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s126;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && ~x9 && ~x7 && x8 && ~x23 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && ~x9 && ~x7 && ~x8 && x14 && x23 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s337;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && ~x9 && ~x7 && ~x8 && x14 && ~x23 )
						begin
							y7 = 1'b1;	
							nx_state = s338;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && x16 && ~x9 && ~x7 && ~x8 && ~x14 )
						nx_state = s1;
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && x8 && x9 && x7 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && x8 && x9 && ~x7 && x23 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s339;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && x8 && x9 && ~x7 && ~x23 )
						begin
							y14 = 1'b1;	
							nx_state = s331;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && x8 && ~x9 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && ~x8 && x7 && x9 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && ~x8 && x7 && ~x9 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && ~x8 && x7 && ~x9 && ~x2 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && ~x8 && x7 && ~x9 && ~x2 && ~x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s340;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && ~x8 && ~x7 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && ~x8 && ~x7 && ~x2 && x3 && x23 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && ~x8 && ~x7 && ~x2 && x3 && ~x23 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && ~x8 && ~x7 && ~x2 && ~x3 && x9 )
						begin
							y14 = 1'b1;	
							nx_state = s286;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && ~x8 && ~x7 && ~x2 && ~x3 && ~x9 && x23 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s341;
						end
					else if( ~x65 && x15 && x66 && ~x21 && ~x22 && ~x16 && ~x8 && ~x7 && ~x2 && ~x3 && ~x9 && ~x23 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x15 && ~x66 && x8 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && x15 && ~x66 && ~x8 && x6 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x65 && x15 && ~x66 && ~x8 && ~x6 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && ~x15 && x16 && x66 && x21 )
						begin
							y14 = 1'b1;	
							nx_state = s286;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && x12 && x8 && x2 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s341;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && x12 && x8 && ~x2 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && x12 && x8 && ~x2 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && x12 && x8 && ~x2 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && x12 && x8 && ~x2 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && x12 && ~x8 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && x12 && ~x8 && ~x2 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && x12 && ~x8 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && ~x12 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && ~x12 && ~x2 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && x23 && ~x12 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && ~x23 && x12 )
						begin
							y14 = 1'b1;	
							nx_state = s286;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && x10 && ~x23 && ~x12 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s341;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && x7 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && x7 && ~x2 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && x7 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && ~x7 && x11 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && ~x7 && x11 && ~x2 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && ~x7 && x11 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && ~x7 && ~x11 && x2 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s341;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && ~x7 && ~x11 && ~x2 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && ~x7 && ~x11 && ~x2 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && ~x7 && ~x11 && ~x2 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && x12 && ~x7 && ~x11 && ~x2 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && x11 && x9 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && x11 && x9 && ~x2 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && x11 && x9 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && x11 && ~x9 && x2 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s341;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && x11 && ~x9 && ~x2 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && x11 && ~x9 && ~x2 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && x11 && ~x9 && ~x2 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && x11 && ~x9 && ~x2 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && ~x11 && x8 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && ~x11 && x8 && ~x2 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && ~x11 && x8 && ~x2 && ~x4 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && ~x11 && ~x8 && x2 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s341;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && ~x11 && ~x8 && ~x2 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && ~x11 && ~x8 && ~x2 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && ~x11 && ~x8 && ~x2 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && x23 && ~x12 && ~x11 && ~x8 && ~x2 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && x22 && ~x10 && ~x23 )
						begin
							y14 = 1'b1;	
							nx_state = s286;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && x7 && x11 )
						nx_state = s1;
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && x7 && ~x11 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && x7 && ~x11 && ~x2 && x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && x7 && ~x11 && ~x2 && x23 && ~x3 )
						begin
							y14 = 1'b1;	
							nx_state = s331;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && x7 && ~x11 && ~x2 && ~x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && x7 && ~x11 && ~x2 && ~x23 && ~x3 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && x10 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && x10 && ~x2 && x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && x10 && ~x2 && x23 && ~x3 )
						begin
							y14 = 1'b1;	
							nx_state = s331;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && x10 && ~x2 && ~x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && x10 && ~x2 && ~x23 && ~x3 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && ~x10 && x8 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && ~x10 && x8 && ~x2 && x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && ~x10 && x8 && ~x2 && x23 && ~x3 )
						begin
							y14 = 1'b1;	
							nx_state = s331;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && ~x10 && x8 && ~x2 && ~x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && ~x10 && x8 && ~x2 && ~x23 && ~x3 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && x9 && ~x7 && ~x10 && ~x8 )
						nx_state = s1;
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && x7 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && x7 && ~x2 && x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && x7 && ~x2 && x23 && ~x3 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && x7 && ~x2 && ~x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s343;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && x7 && ~x2 && ~x23 && ~x3 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && x8 && x12 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && x8 && x12 && ~x2 && x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && x8 && x12 && ~x2 && x23 && ~x3 )
						begin
							y14 = 1'b1;	
							nx_state = s331;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && x8 && x12 && ~x2 && ~x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && x8 && x12 && ~x2 && ~x23 && ~x3 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && x8 && ~x12 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && x8 && ~x12 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && x8 && ~x12 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && x8 && ~x12 && x23 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && x8 && ~x12 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && ~x8 && x11 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && ~x8 && x11 && ~x2 && x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && ~x8 && x11 && ~x2 && x23 && ~x3 )
						begin
							y14 = 1'b1;	
							nx_state = s331;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && ~x8 && x11 && ~x2 && ~x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && ~x8 && x11 && ~x2 && ~x23 && ~x3 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x15 && x16 && x66 && ~x21 && ~x22 && ~x9 && ~x7 && ~x8 && ~x11 )
						nx_state = s1;
					else if( ~x65 && ~x15 && x16 && ~x66 && x8 && x7 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && ~x15 && x16 && ~x66 && x8 && ~x7 && x9 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && ~x15 && x16 && ~x66 && x8 && ~x7 && ~x9 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x15 && x16 && ~x66 && x8 && ~x7 && ~x9 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x15 && x16 && ~x66 && x8 && ~x7 && ~x9 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x15 && x16 && ~x66 && x8 && ~x7 && ~x9 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x15 && x16 && ~x66 && ~x8 && x7 && x11 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && ~x15 && x16 && ~x66 && ~x8 && x7 && ~x11 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x15 && x16 && ~x66 && ~x8 && x7 && ~x11 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x15 && x16 && ~x66 && ~x8 && x7 && ~x11 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x15 && x16 && ~x66 && ~x8 && x7 && ~x11 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x15 && x16 && ~x66 && ~x8 && ~x7 && x10 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && ~x15 && x16 && ~x66 && ~x8 && ~x7 && ~x10 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x15 && x16 && ~x66 && ~x8 && ~x7 && ~x10 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x15 && x16 && ~x66 && ~x8 && ~x7 && ~x10 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x15 && x16 && ~x66 && ~x8 && ~x7 && ~x10 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x15 && ~x16 && x66 && x21 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s340;
						end
					else if( ~x65 && ~x15 && ~x16 && x66 && ~x21 && x22 && x23 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x65 && ~x15 && ~x16 && x66 && ~x21 && x22 && x23 && ~x2 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && ~x15 && ~x16 && x66 && ~x21 && x22 && x23 && ~x2 && ~x4 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && ~x15 && ~x16 && x66 && ~x21 && x22 && ~x23 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s81;
						end
					else if( ~x65 && ~x15 && ~x16 && x66 && ~x21 && ~x22 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( ~x65 && ~x15 && ~x16 && x66 && ~x21 && ~x22 && ~x2 && x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && ~x15 && ~x16 && x66 && ~x21 && ~x22 && ~x2 && x23 && ~x3 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x65 && ~x15 && ~x16 && x66 && ~x21 && ~x22 && ~x2 && ~x23 && x3 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && ~x15 && ~x16 && x66 && ~x21 && ~x22 && ~x2 && ~x23 && ~x3 )
						begin
							y14 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x65 && ~x15 && ~x16 && ~x66 && x6 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x65 && ~x15 && ~x16 && ~x66 && ~x6 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else nx_state = s76;
				s77 : if( x65 && x66 && x67 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && x67 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && x67 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && x66 && x67 && x22 && ~x17 )
						nx_state = s1;
					else if( x65 && x66 && x67 && ~x22 && x18 && x13 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && x66 && x67 && ~x22 && x18 && x13 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x66 && x67 && ~x22 && x18 && ~x13 && x12 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && x66 && x67 && ~x22 && x18 && ~x13 && x12 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x66 && x67 && ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && x66 && x67 && ~x22 && ~x18 )
						nx_state = s1;
					else if( x65 && x66 && ~x67 && x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && ~x67 && x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && ~x67 && x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x66 && ~x67 && x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x65 && x66 && ~x67 && x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x66 && ~x67 && x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x66 && ~x67 && x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x66 && ~x67 && x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( x65 && x66 && ~x67 && ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x66 && ~x67 && ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x66 && ~x67 && ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x66 && ~x67 && ~x21 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x66 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x65 && ~x66 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && x23 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x23 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x23 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x23 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && x23 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x23 && x18 && x14 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x23 && x18 && ~x14 && x13 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x22 && x23 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && x23 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && x23 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x22 && x23 && ~x20 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x23 && x15 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x23 && ~x15 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x65 && x66 && x67 && x68 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && x66 && x67 && x68 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && x66 && x67 && x68 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && x68 && x21 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && x68 && ~x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s344;
						end
					else if( ~x65 && x66 && x67 && ~x68 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && x66 && x67 && ~x68 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && x66 && x67 && ~x68 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x68 && x62 && ~x61 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x68 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && x21 && x68 )
						begin
							y8 = 1'b1;	y18 = 1'b1;	
							nx_state = s82;
						end
					else if( ~x65 && x66 && ~x67 && x21 && ~x68 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s143;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && x68 && x22 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && x68 && x22 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && x68 && x22 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && ~x21 && x68 && x22 && ~x7 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && ~x21 && x68 && ~x22 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && x68 && ~x22 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && x68 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && ~x21 && x68 && ~x22 && ~x4 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && ~x21 && ~x68 && x23 && x22 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && ~x68 && x23 && ~x22 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && ~x68 && x23 && ~x22 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && ~x68 && x23 && ~x22 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && ~x21 && ~x68 && x23 && ~x22 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && ~x21 && ~x68 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && ~x66 && x68 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x66 && x68 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x66 && x68 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x68 && x20 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x68 && ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x66 && x68 && ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x66 && x68 && ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x68 && ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x68 && ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x65 && ~x66 && x68 && ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x65 && ~x66 && x68 && ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x68 && ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x68 && x24 && x26 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x65 && ~x66 && ~x68 && x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && ~x66 && ~x68 && x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && ~x66 && ~x68 && x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x68 && x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x68 && ~x24 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && ~x68 && ~x24 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && ~x68 && ~x24 && x25 && x19 && ~x14 && ~x13 && x26 )
						nx_state = s77;
					else if( ~x65 && ~x66 && ~x68 && ~x24 && x25 && x19 && ~x14 && ~x13 && ~x26 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x68 && ~x24 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && x4 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && x19 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && x20 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && ~x20 && x21 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && ~x20 && ~x21 && x22 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && ~x20 && ~x21 && ~x22 && x16 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && ~x20 && ~x21 && ~x22 && x16 && ~x11 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && ~x20 && ~x21 && ~x22 && x16 && ~x11 && ~x12 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && ~x20 && ~x21 && ~x22 && x16 && ~x11 && ~x12 && ~x10 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && ~x20 && ~x21 && ~x22 && ~x16 && x17 && x10 && x12 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && ~x20 && ~x21 && ~x22 && ~x16 && x17 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && ~x20 && ~x21 && ~x22 && ~x16 && x17 && ~x10 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && x26 && ~x4 && ~x19 && ~x20 && ~x21 && ~x22 && ~x16 && ~x17 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x68 && ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else nx_state = s77;
				s78 : if( x65 && x66 && x61 && x60 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x66 && x61 && x60 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x66 && x61 && x60 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x66 && x61 && x60 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x66 && x61 && ~x60 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x66 && x61 && ~x60 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x66 && x61 && ~x60 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x65 && x66 && x61 && ~x60 && x62 && ~x18 )
						nx_state = s1;
					else if( x65 && x66 && x61 && ~x60 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && x61 && ~x60 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && x61 && ~x60 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x65 && x66 && x61 && ~x60 && ~x62 && ~x18 )
						nx_state = s39;
					else if( x65 && x66 && ~x61 && x60 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && ~x61 && x60 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && ~x61 && x60 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x65 && x66 && ~x61 && x60 && ~x18 )
						nx_state = s39;
					else if( x65 && x66 && ~x61 && ~x60 && x62 )
						nx_state = s40;
					else if( x65 && x66 && ~x61 && ~x60 && ~x62 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s263;
						end
					else if( x65 && ~x66 && x67 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x67 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x67 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && ~x68 && x22 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && ~x68 && ~x22 )
						begin
							y28 = 1'b1;	
							nx_state = s94;
						end
					else if( ~x65 && x21 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && ~x21 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && ~x21 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x21 && ~x7 )
						nx_state = s1;
					else nx_state = s78;
				s79 : if( x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x21 && x22 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x10 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s226;
						end
					else if( ~x21 && ~x22 && ~x10 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x21 && ~x22 && ~x10 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x21 && ~x22 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x10 && ~x4 )
						nx_state = s1;
					else nx_state = s79;
				s80 : if( x22 )
						nx_state = s1;
					else if( ~x22 && x21 )
						nx_state = s1;
					else if( ~x22 && ~x21 && x23 && x15 && x7 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s81;
						end
					else if( ~x22 && ~x21 && x23 && x15 && ~x7 && x9 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x22 && ~x21 && x23 && x15 && ~x7 && ~x9 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x22 && ~x21 && x23 && ~x15 && x7 && x9 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s330;
						end
					else if( ~x22 && ~x21 && x23 && ~x15 && x7 && ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x22 && ~x21 && x23 && ~x15 && ~x7 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s330;
						end
					else if( ~x22 && ~x21 && ~x23 )
						begin
							y14 = 1'b1;	
							nx_state = s285;
						end
					else nx_state = s80;
				s81 : if( x21 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s336;
						end
					else if( ~x21 && x22 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x19 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else nx_state = s81;
				s82 : if( x21 && x66 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( x21 && ~x66 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( x21 && ~x66 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( x21 && ~x66 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x21 && ~x66 && ~x3 )
						nx_state = s1;
					else if( ~x21 && x66 && x22 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s232;
						end
					else if( ~x21 && x66 && ~x22 && x16 && x15 && x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s219;
						end
					else if( ~x21 && x66 && ~x22 && x16 && x15 && ~x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s309;
						end
					else if( ~x21 && x66 && ~x22 && x16 && ~x15 && x10 )
						begin
							y2 = 1'b1;	y16 = 1'b1;	y24 = 1'b1;	
							nx_state = s124;
						end
					else if( ~x21 && x66 && ~x22 && x16 && ~x15 && ~x10 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s310;
						end
					else if( ~x21 && x66 && ~x22 && ~x16 && x17 && x10 && x15 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s219;
						end
					else if( ~x21 && x66 && ~x22 && ~x16 && x17 && x10 && ~x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s308;
						end
					else if( ~x21 && x66 && ~x22 && ~x16 && x17 && ~x10 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s79;
						end
					else if( ~x21 && x66 && ~x22 && ~x16 && ~x17 && x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s219;
						end
					else if( ~x21 && x66 && ~x22 && ~x16 && ~x17 && ~x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s311;
						end
					else if( ~x21 && ~x66 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && ~x66 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && ~x66 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && ~x66 && ~x8 )
						nx_state = s1;
					else nx_state = s82;
				s83 : if( x65 && x66 && x68 && x21 && x20 )
						nx_state = s1;
					else if( x65 && x66 && x68 && x21 && ~x20 && x18 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y21 = 1'b1;	
							nx_state = s299;
						end
					else if( x65 && x66 && x68 && x21 && ~x20 && ~x18 && x15 && x10 && x11 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s192;
						end
					else if( x65 && x66 && x68 && x21 && ~x20 && ~x18 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s193;
						end
					else if( x65 && x66 && x68 && x21 && ~x20 && ~x18 && x15 && x10 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y13 = 1'b1;	
							nx_state = s192;
						end
					else if( x65 && x66 && x68 && x21 && ~x20 && ~x18 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s300;
						end
					else if( x65 && x66 && x68 && x21 && ~x20 && ~x18 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s192;
						end
					else if( x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && x10 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && x10 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && x10 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && x10 && ~x19 )
						nx_state = s1;
					else if( x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && ~x10 && x12 && x11 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s199;
						end
					else if( x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && ~x10 && x12 && ~x11 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && ~x10 && x12 && ~x11 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && ~x10 && x12 && ~x11 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && ~x10 && x12 && ~x11 && ~x19 )
						nx_state = s1;
					else if( x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && ~x10 && ~x12 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && ~x10 && ~x12 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && ~x10 && ~x12 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && x16 && ~x10 && ~x12 && ~x19 )
						nx_state = s1;
					else if( x65 && x66 && x68 && x21 && ~x20 && ~x18 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s201;
						end
					else if( x65 && x66 && x68 && ~x21 )
						nx_state = s1;
					else if( x65 && x66 && ~x68 && x60 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && x16 && x4 && x11 && x12 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s15;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && x16 && x4 && x11 && ~x12 && x13 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s345;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && x16 && x4 && x11 && ~x12 && ~x13 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && x16 && x4 && ~x11 && x13 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && x16 && x4 && ~x11 && ~x13 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && x16 && ~x4 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && x11 && x9 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && x11 && ~x9 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && x11 && ~x9 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && x11 && ~x9 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && x11 && ~x9 && ~x18 )
						nx_state = s1;
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && ~x11 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && ~x11 && ~x8 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && ~x11 && ~x8 && ~x12 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && ~x11 && ~x8 && ~x12 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && ~x11 && ~x8 && ~x12 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && x13 && ~x11 && ~x8 && ~x12 && ~x18 )
						nx_state = s1;
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && x11 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && ~x11 && x12 && x10 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && ~x11 && x12 && ~x10 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && ~x11 && x12 && ~x10 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && ~x11 && x12 && ~x10 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && ~x11 && x12 && ~x10 && ~x18 )
						nx_state = s1;
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && ~x11 && ~x12 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && ~x11 && ~x12 && ~x7 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && ~x11 && ~x12 && ~x7 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && ~x11 && ~x12 && ~x7 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && x17 && ~x13 && ~x11 && ~x12 && ~x7 && ~x18 )
						nx_state = s1;
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && ~x17 && x45 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x16 && ~x17 && ~x45 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && x66 && ~x68 && ~x60 && ~x61 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && x21 && x68 && x18 )
						begin
							y14 = 1'b1;	y19 = 1'b1;	
							nx_state = s116;
						end
					else if( x65 && ~x66 && x67 && x21 && x68 && ~x18 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s117;
						end
					else if( x65 && ~x66 && x67 && x21 && ~x68 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x67 && x21 && ~x68 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x67 && x21 && ~x68 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && x21 && ~x68 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && ~x21 && x22 && x68 && x8 && x23 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x66 && x67 && ~x21 && x22 && x68 && x8 && x23 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x66 && x67 && ~x21 && x22 && x68 && x8 && x23 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && ~x21 && x22 && x68 && x8 && ~x23 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x66 && x67 && ~x21 && x22 && x68 && x8 && ~x23 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x66 && x67 && ~x21 && x22 && x68 && x8 && ~x23 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && ~x21 && x22 && x68 && ~x8 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && ~x21 && x22 && ~x68 && x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x67 && ~x21 && x22 && ~x68 && x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x67 && ~x21 && x22 && ~x68 && x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && ~x21 && x22 && ~x68 && x19 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && ~x21 && x22 && ~x68 && ~x19 && x18 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x67 && ~x21 && x22 && ~x68 && ~x19 && x18 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x67 && ~x21 && x22 && ~x68 && ~x19 && x18 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && ~x21 && x22 && ~x68 && ~x19 && x18 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && ~x21 && x22 && ~x68 && ~x19 && ~x18 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && x67 && ~x21 && ~x22 && x68 && x23 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x66 && x67 && ~x21 && ~x22 && x68 && x23 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x66 && x67 && ~x21 && ~x22 && x68 && x23 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && ~x21 && ~x22 && x68 && x23 && ~x9 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && ~x21 && ~x22 && x68 && ~x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x66 && x67 && ~x21 && ~x22 && x68 && ~x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x66 && x67 && ~x21 && ~x22 && x68 && ~x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && ~x21 && ~x22 && x68 && ~x23 && ~x8 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && ~x21 && ~x22 && ~x68 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x67 && ~x21 && ~x22 && ~x68 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x67 && ~x21 && ~x22 && ~x68 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && ~x21 && ~x22 && ~x68 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && x17 && x20 && x16 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && x17 && x20 && ~x16 )
						begin
							y24 = 1'b1;	
							nx_state = s346;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && x17 && ~x20 && x16 )
						begin
							y13 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	y29 = 1'b1;	y30 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s347;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && x17 && ~x20 && ~x16 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && ~x17 && x16 && x4 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s348;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && ~x17 && x16 && ~x4 )
						begin
							y10 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s349;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && ~x17 && ~x16 && x20 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && ~x17 && ~x16 && x20 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && ~x17 && ~x16 && x20 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && ~x17 && ~x16 && x20 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && x14 && ~x17 && ~x16 && ~x20 )
						begin
							y15 = 1'b1;	y28 = 1'b1;	
							nx_state = s350;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && x15 && x17 && x20 && x16 )
						begin
							y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && x15 && x17 && x20 && ~x16 )
						begin
							y4 = 1'b1;	y12 = 1'b1;	y27 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && x15 && x17 && ~x20 && x16 )
						begin
							y24 = 1'b1;	
							nx_state = s346;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && x15 && x17 && ~x20 && ~x16 )
						begin
							y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && x15 && ~x17 && x16 )
						begin
							y15 = 1'b1;	y28 = 1'b1;	
							nx_state = s350;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && x15 && ~x17 && ~x16 && x13 )
						begin
							y15 = 1'b1;	y28 = 1'b1;	
							nx_state = s350;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && x15 && ~x17 && ~x16 && ~x13 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && x15 && ~x17 && ~x16 && ~x13 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && x15 && ~x17 && ~x16 && ~x13 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && x15 && ~x17 && ~x16 && ~x13 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && x17 && x6 && x16 && x7 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && x17 && x6 && x16 && ~x7 && x5 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && x17 && x6 && x16 && ~x7 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && x17 && x6 && ~x16 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && x17 && ~x6 && x7 && x16 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && x17 && ~x6 && x7 && ~x16 && x5 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && x17 && ~x6 && x7 && ~x16 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && x17 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && ~x17 && x16 && x12 )
						begin
							y15 = 1'b1;	y28 = 1'b1;	
							nx_state = s350;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && ~x17 && x16 && ~x12 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && ~x17 && x16 && ~x12 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && ~x17 && x16 && ~x12 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && ~x17 && x16 && ~x12 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && ~x17 && ~x16 && x11 )
						begin
							y15 = 1'b1;	y28 = 1'b1;	
							nx_state = s350;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && ~x17 && ~x16 && ~x11 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && ~x17 && ~x16 && ~x11 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && ~x17 && ~x16 && ~x11 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && x19 && ~x14 && ~x15 && ~x17 && ~x16 && ~x11 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && x20 && x14 && x13 )
						begin
							y10 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s349;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && x20 && x14 && ~x13 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && x20 && ~x14 && x13 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	y19 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s349;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && x20 && ~x14 && ~x13 && x6 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s102;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && x20 && ~x14 && ~x13 && ~x6 && x5 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && x20 && ~x14 && ~x13 && ~x6 && x5 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && x20 && ~x14 && ~x13 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && ~x20 && x15 && x14 )
						begin
							y10 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s349;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && ~x20 && x15 && ~x14 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s102;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && ~x20 && ~x15 && x14 )
						begin
							y15 = 1'b1;	y28 = 1'b1;	
							nx_state = s350;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && x17 && ~x20 && ~x15 && ~x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && x13 && x12 && x14 )
						begin
							y15 = 1'b1;	y28 = 1'b1;	
							nx_state = s350;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && x13 && x12 && ~x14 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && x13 && x12 && ~x14 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && x13 && x12 && ~x14 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && x13 && x12 && ~x14 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && x13 && ~x12 )
						begin
							y15 = 1'b1;	y28 = 1'b1;	
							nx_state = s350;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && ~x13 && x11 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && ~x13 && x11 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && ~x13 && x11 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && ~x13 && x11 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && x20 && ~x13 && ~x11 )
						begin
							y15 = 1'b1;	y28 = 1'b1;	
							nx_state = s350;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && x14 && x13 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s348;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && x14 && ~x13 && x15 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s348;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && x14 && ~x13 && ~x15 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && x14 && ~x13 && ~x15 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && x14 && ~x13 && ~x15 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && x14 && ~x13 && ~x15 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && ~x14 && x15 && x12 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s348;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && ~x14 && x15 && ~x12 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && ~x14 && x15 && ~x12 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && ~x14 && x15 && ~x12 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && ~x14 && x15 && ~x12 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && ~x14 && ~x15 && x11 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s348;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && ~x14 && ~x15 && ~x11 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && ~x14 && ~x15 && ~x11 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && ~x14 && ~x15 && ~x11 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && x18 && ~x19 && ~x17 && ~x20 && ~x14 && ~x15 && ~x11 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && x14 && x15 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && x14 && ~x15 && x16 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && x14 && ~x15 && ~x16 && x4 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s348;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && x14 && ~x15 && ~x16 && ~x4 )
						begin
							y4 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && ~x14 && x16 && x15 && x13 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && ~x14 && x16 && x15 && ~x13 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	y32 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && ~x14 && x16 && ~x15 && x4 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s348;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && ~x14 && x16 && ~x15 && ~x4 )
						begin
							y4 = 1'b1;	y17 = 1'b1;	y29 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && ~x14 && ~x16 && x15 )
						begin
							y4 = 1'b1;	y29 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && ~x14 && ~x16 && ~x15 && x4 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	y21 = 1'b1;	y28 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && x19 && ~x14 && ~x16 && ~x15 && ~x4 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && ~x19 && x16 && x14 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	y21 = 1'b1;	y28 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && ~x19 && x16 && ~x14 && x4 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && ~x19 && x16 && ~x14 && ~x4 )
						begin
							y16 = 1'b1;	y28 = 1'b1;	
							nx_state = s352;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && ~x19 && ~x16 && x13 && x14 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	y21 = 1'b1;	y28 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && ~x19 && ~x16 && x13 && x14 && ~x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && ~x19 && ~x16 && x13 && ~x14 && x4 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && ~x19 && ~x16 && x13 && ~x14 && ~x4 )
						begin
							y4 = 1'b1;	y12 = 1'b1;	y27 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && ~x19 && ~x16 && ~x13 && x4 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && x20 && ~x19 && ~x16 && ~x13 && ~x4 )
						begin
							y24 = 1'b1;	
							nx_state = s346;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && x14 && x19 && x15 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && x14 && x19 && ~x15 && x16 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && x14 && x19 && ~x15 && ~x16 && x4 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s348;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && x14 && x19 && ~x15 && ~x16 && ~x4 )
						begin
							y4 = 1'b1;	y29 = 1'b1;	y32 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && x14 && ~x19 && x16 )
						begin
							y24 = 1'b1;	
							nx_state = s346;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && x14 && ~x19 && ~x16 && x15 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && x14 && ~x19 && ~x16 && x15 && ~x13 )
						begin
							y4 = 1'b1;	y12 = 1'b1;	y27 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && x14 && ~x19 && ~x16 && ~x15 )
						begin
							y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && x15 && x16 && x19 && x13 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && x15 && x16 && x19 && ~x13 )
						begin
							y4 = 1'b1;	y29 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && x15 && x16 && ~x19 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && x15 && ~x16 && x4 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s348;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && x15 && ~x16 && ~x4 && x19 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && x15 && ~x16 && ~x4 && ~x19 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && ~x15 && x4 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s348;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && ~x15 && ~x4 && x19 && x16 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && ~x15 && ~x4 && x19 && ~x16 )
						begin
							y4 = 1'b1;	y12 = 1'b1;	y27 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && ~x15 && ~x4 && ~x19 && x16 )
						begin
							y16 = 1'b1;	y28 = 1'b1;	
							nx_state = s352;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && x17 && ~x20 && ~x14 && ~x15 && ~x4 && ~x19 && ~x16 )
						begin
							y13 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	y29 = 1'b1;	y30 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s347;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && ~x17 && x4 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s348;
						end
					else if( x65 && ~x66 && ~x67 && x68 && ~x3 && ~x18 && ~x17 && ~x4 )
						begin
							y4 = 1'b1;	y17 = 1'b1;	
							nx_state = s353;
						end
					else if( x65 && ~x66 && ~x67 && ~x68 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x65 && ~x66 && ~x67 && ~x68 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x67 && ~x68 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x67 && ~x68 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && ~x68 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && ~x68 && ~x21 && x23 && x22 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( x65 && ~x66 && ~x67 && ~x68 && ~x21 && x23 && x22 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x66 && ~x67 && ~x68 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x66 && ~x67 && ~x68 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && ~x68 && ~x21 && x23 && x22 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && ~x68 && ~x21 && x23 && ~x22 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x66 && ~x67 && ~x68 && ~x21 && x23 && ~x22 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x66 && ~x67 && ~x68 && ~x21 && x23 && ~x22 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && ~x68 && ~x21 && x23 && ~x22 && ~x20 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x23 && x18 && x14 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x23 && x18 && x14 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x23 && x18 && ~x14 && x13 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x23 && x18 && ~x14 && x13 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x67 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && x67 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && x67 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x67 && x62 && ~x61 )
						nx_state = s1;
					else if( ~x65 && x67 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && x67 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && x67 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && x67 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && x67 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x67 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( ~x65 && x67 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x67 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x67 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x67 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x67 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x67 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x67 )
						nx_state = s1;
					else nx_state = s83;
				s84 : if( x21 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x21 && x23 && x22 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s354;
						end
					else if( ~x21 && x23 && ~x22 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s80;
						end
					else if( ~x21 && ~x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s80;
						end
					else nx_state = s84;
				s85 : if( x65 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x65 && x22 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s340;
						end
					else if( ~x65 && ~x22 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s337;
						end
					else nx_state = s85;
				s86 : if( x65 && x66 && x67 && x23 )
						nx_state = s1;
					else if( x65 && x66 && x67 && ~x23 && x6 && x15 && x8 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x66 && x67 && ~x23 && x6 && x15 && ~x8 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x65 && x66 && x67 && ~x23 && x6 && ~x15 && x16 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x66 && x67 && ~x23 && x6 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s122;
						end
					else if( x65 && x66 && x67 && ~x23 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x66 && ~x67 && x60 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( x65 && x66 && ~x67 && ~x60 && x61 && x62 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && x66 && ~x67 && ~x60 && x61 && ~x62 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && x16 && x12 && x7 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s254;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && x16 && x12 && ~x7 && x14 && x11 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && x16 && x12 && ~x7 && x14 && ~x11 )
						begin
							y15 = 1'b1;	
							nx_state = s355;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && x16 && x12 && ~x7 && ~x14 )
						nx_state = s40;
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && x16 && ~x12 && x7 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && x16 && ~x12 && ~x7 && x13 && x11 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && x16 && ~x12 && ~x7 && x13 && ~x11 )
						begin
							y15 = 1'b1;	
							nx_state = s355;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && x16 && ~x12 && ~x7 && ~x13 )
						nx_state = s40;
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && ~x16 && x11 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s291;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && ~x16 && x11 && ~x7 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s231;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && ~x16 && x11 && ~x7 && ~x12 )
						begin
							y12 = 1'b1;	
							nx_state = s210;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && ~x16 && ~x11 && x6 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s74;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && ~x16 && ~x11 && ~x6 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && ~x16 && ~x11 && ~x6 && ~x2 && x12 && x7 )
						begin
							y11 = 1'b1;	
							nx_state = s356;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && ~x16 && ~x11 && ~x6 && ~x2 && x12 && ~x7 )
						begin
							y11 = 1'b1;	
							nx_state = s357;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && ~x16 && ~x11 && ~x6 && ~x2 && ~x12 && x7 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && x15 && ~x16 && ~x11 && ~x6 && ~x2 && ~x12 && ~x7 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && x6 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s74;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && x7 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && x7 && ~x2 && x12 )
						begin
							y11 = 1'b1;	
							nx_state = s357;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && x7 && ~x2 && ~x12 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && x12 && x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && x12 && x11 && ~x2 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s260;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && x12 && ~x11 && x9 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && x12 && ~x11 && x9 && ~x2 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s260;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && x12 && ~x11 && ~x9 )
						nx_state = s40;
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && ~x12 && x11 && x10 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && ~x12 && x11 && x10 && ~x2 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s260;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && ~x12 && x11 && ~x10 )
						nx_state = s40;
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && ~x12 && ~x11 && x8 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && ~x12 && ~x11 && x8 && ~x2 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s260;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && x16 && ~x7 && ~x12 && ~x11 && ~x8 )
						nx_state = s40;
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && ~x16 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && ~x16 && ~x2 && x7 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && x62 && ~x15 && ~x6 && ~x16 && ~x2 && ~x7 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s68;
						end
					else if( x65 && x66 && ~x67 && ~x60 && ~x61 && ~x62 )
						begin
							y3 = 1'b1;	
							nx_state = s65;
						end
					else if( x65 && ~x66 && x21 && x17 && x16 && x13 && x18 && x15 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && x21 && x17 && x16 && x13 && x18 && ~x15 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && ~x66 && x21 && x17 && x16 && x13 && ~x18 && x14 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && ~x66 && x21 && x17 && x16 && x13 && ~x18 && ~x14 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x65 && ~x66 && x21 && x17 && x16 && ~x13 && x14 && x18 && x15 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x65 && ~x66 && x21 && x17 && x16 && ~x13 && x14 && x18 && ~x15 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s288;
						end
					else if( x65 && ~x66 && x21 && x17 && x16 && ~x13 && x14 && ~x18 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s288;
						end
					else if( x65 && ~x66 && x21 && x17 && x16 && ~x13 && ~x14 && x18 && x15 && x6 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && x21 && x17 && x16 && ~x13 && ~x14 && x18 && x15 && ~x6 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x21 && x17 && x16 && ~x13 && ~x14 && x18 && x15 && ~x6 && x4 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && x21 && x17 && x16 && ~x13 && ~x14 && x18 && x15 && ~x6 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && x21 && x17 && x16 && ~x13 && ~x14 && x18 && ~x15 && x5 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && x21 && x17 && x16 && ~x13 && ~x14 && x18 && ~x15 && ~x5 && x4 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x21 && x17 && x16 && ~x13 && ~x14 && x18 && ~x15 && ~x5 && x4 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && x21 && x17 && x16 && ~x13 && ~x14 && x18 && ~x15 && ~x5 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && x21 && x17 && x16 && ~x13 && ~x14 && ~x18 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && x13 && x18 && x15 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && x13 && x18 && ~x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && x13 && x18 && ~x15 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && x13 && ~x18 && x14 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && x13 && ~x18 && x14 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && x13 && ~x18 && x14 && ~x2 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && x13 && ~x18 && ~x14 && x12 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && x13 && ~x18 && ~x14 && x12 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && x13 && ~x18 && ~x14 && x12 && ~x2 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && x13 && ~x18 && ~x14 && ~x12 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && x13 && ~x18 && ~x14 && ~x12 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && x13 && ~x18 && ~x14 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && x21 && x17 && ~x16 && x13 && ~x18 && ~x14 && ~x12 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && x18 && x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && x18 && x15 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && x18 && ~x15 && x12 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && x18 && ~x15 && x12 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && x18 && ~x15 && ~x12 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && x18 && ~x15 && ~x12 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && x18 && ~x15 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && x18 && ~x15 && ~x12 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && ~x18 && x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && ~x18 && x11 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && ~x18 && x11 && ~x2 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && ~x18 && ~x11 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && ~x18 && ~x11 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && ~x18 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && x14 && ~x18 && ~x11 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && x15 && x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && x15 && x11 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && x15 && ~x11 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && x15 && ~x11 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && x15 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && x15 && ~x11 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && ~x15 && x10 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && ~x15 && x10 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && ~x15 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && ~x15 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && ~x15 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && x18 && ~x15 && ~x10 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && ~x18 && x10 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && ~x18 && x10 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && ~x18 && x10 && ~x2 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && ~x18 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && ~x18 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && ~x18 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && x21 && x17 && ~x16 && ~x13 && ~x14 && ~x18 && ~x10 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && x21 && ~x17 && x16 && x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x66 && x21 && ~x17 && x16 && x14 && ~x13 && x15 && x18 && x12 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( x65 && ~x66 && x21 && ~x17 && x16 && x14 && ~x13 && x15 && x18 && ~x12 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s169;
						end
					else if( x65 && ~x66 && x21 && ~x17 && x16 && x14 && ~x13 && x15 && ~x18 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( x65 && ~x66 && x21 && ~x17 && x16 && x14 && ~x13 && ~x15 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s174;
						end
					else if( x65 && ~x66 && x21 && ~x17 && x16 && ~x14 && x15 && x18 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( x65 && ~x66 && x21 && ~x17 && x16 && ~x14 && x15 && x18 && ~x13 )
						begin
							y24 = 1'b1;	
							nx_state = s346;
						end
					else if( x65 && ~x66 && x21 && ~x17 && x16 && ~x14 && x15 && ~x18 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s346;
						end
					else if( x65 && ~x66 && x21 && ~x17 && x16 && ~x14 && x15 && ~x18 && ~x13 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s169;
						end
					else if( x65 && ~x66 && x21 && ~x17 && x16 && ~x14 && ~x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && x21 && ~x17 && x16 && ~x14 && ~x15 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && x21 && ~x17 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && x13 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && x21 && ~x17 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s300;
						end
					else if( x65 && ~x66 && x21 && ~x17 && ~x16 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && x21 && ~x17 && ~x16 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && x21 && ~x17 && ~x16 && ~x2 && ~x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s51;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && x10 && x15 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s288;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && x10 && ~x15 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s300;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && ~x10 && x15 && x6 && x14 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s360;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && ~x10 && x15 && x6 && ~x14 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && ~x10 && x15 && ~x6 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && ~x10 && x15 && ~x6 && x4 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && ~x10 && x15 && ~x6 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && ~x10 && ~x15 && x5 && x14 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && ~x10 && ~x15 && x5 && ~x14 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && ~x10 && ~x15 && ~x5 && x4 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && ~x10 && ~x15 && ~x5 && x4 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && x19 && ~x10 && ~x15 && ~x5 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && x13 && x15 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s300;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && x13 && ~x15 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s360;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && ~x13 && x15 && x6 && x14 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && ~x13 && x15 && x6 && ~x14 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && ~x13 && x15 && ~x6 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && ~x13 && x15 && ~x6 && x4 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && ~x13 && x15 && ~x6 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && ~x13 && ~x15 && x5 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && ~x13 && ~x15 && x5 && ~x14 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && ~x13 && ~x15 && ~x5 && x4 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && ~x13 && ~x15 && ~x5 && x4 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && x18 && ~x19 && ~x13 && ~x15 && ~x5 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && x13 && x15 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && x13 && ~x15 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s288;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && x14 && x19 && x15 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s300;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && x14 && x19 && ~x15 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s360;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && x14 && ~x19 && x15 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s360;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && x14 && ~x19 && ~x15 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && ~x14 && x15 && x6 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && ~x14 && x15 && ~x6 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && ~x14 && x15 && ~x6 && x4 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && ~x14 && x15 && ~x6 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && ~x14 && ~x15 && x5 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && ~x14 && ~x15 && ~x5 && x4 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && ~x14 && ~x15 && ~x5 && x4 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && x16 && ~x18 && ~x13 && ~x14 && ~x15 && ~x5 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && x19 && x10 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && x19 && ~x10 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && x19 && ~x10 && ~x2 && x14 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && x19 && ~x10 && ~x2 && x14 && ~x3 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && x19 && ~x10 && ~x2 && ~x14 && x12 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && x19 && ~x10 && ~x2 && ~x14 && x12 && ~x3 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && x19 && ~x10 && ~x2 && ~x14 && ~x12 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && x19 && ~x10 && ~x2 && ~x14 && ~x12 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && x19 && ~x10 && ~x2 && ~x14 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && x19 && ~x10 && ~x2 && ~x14 && ~x12 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && ~x19 && x13 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s288;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && ~x19 && ~x13 && x14 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && ~x19 && ~x13 && x14 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && ~x19 && ~x13 && x14 && ~x2 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && ~x19 && ~x13 && ~x14 && x11 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && ~x19 && ~x13 && ~x14 && ~x11 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && ~x19 && ~x13 && ~x14 && ~x11 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && ~x19 && ~x13 && ~x14 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && x15 && ~x19 && ~x13 && ~x14 && ~x11 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && x10 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && x14 && x13 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && x14 && x13 && ~x3 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && x14 && ~x13 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && x14 && ~x13 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && x14 && ~x13 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && x14 && ~x13 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && ~x14 && x11 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && ~x14 && x11 && ~x3 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && ~x14 && ~x11 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && ~x14 && ~x11 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && ~x14 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && x19 && ~x2 && ~x10 && ~x14 && ~x11 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && x13 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && x13 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && ~x13 && x14 && x12 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && ~x13 && x14 && ~x12 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && ~x13 && x14 && ~x12 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && ~x13 && x14 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && ~x13 && x14 && ~x12 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && ~x13 && ~x14 && x10 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && ~x13 && ~x14 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && ~x13 && ~x14 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && ~x13 && ~x14 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && x18 && ~x15 && ~x19 && ~x13 && ~x14 && ~x10 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && x13 && x15 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && x13 && ~x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && x13 && ~x15 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && x14 && x15 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && x14 && x15 && ~x3 && x19 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && x14 && x15 && ~x3 && ~x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && x14 && ~x15 && x12 && x19 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && x14 && ~x15 && x12 && x19 && ~x3 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && x14 && ~x15 && x12 && ~x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && x14 && ~x15 && ~x12 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && x14 && ~x15 && ~x12 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && x14 && ~x15 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && x14 && ~x15 && ~x12 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && x15 && x11 && x19 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && x15 && x11 && x19 && ~x3 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && x15 && x11 && ~x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && x15 && ~x11 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && x15 && ~x11 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && x15 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && x15 && ~x11 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && ~x15 && x10 && x19 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && ~x15 && x10 && x19 && ~x3 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && ~x15 && x10 && ~x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && ~x15 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && ~x15 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && ~x15 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && x22 && ~x16 && ~x18 && ~x13 && ~x2 && ~x14 && ~x15 && ~x10 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && x13 && x15 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && x13 && ~x15 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s288;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && ~x13 && x15 && x6 && x14 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s300;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && ~x13 && x15 && x6 && ~x14 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && ~x13 && x15 && ~x6 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && ~x13 && x15 && ~x6 && x4 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && ~x13 && x15 && ~x6 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && ~x13 && ~x15 && x5 && x14 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s360;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && ~x13 && ~x15 && x5 && ~x14 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && ~x13 && ~x15 && ~x5 && x4 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && ~x13 && ~x15 && ~x5 && x4 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && x18 && ~x13 && ~x15 && ~x5 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && ~x18 && x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && ~x18 && x14 && ~x13 && x15 && x16 )
						begin
							y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && ~x18 && x14 && ~x13 && x15 && ~x16 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && ~x18 && x14 && ~x13 && ~x15 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && ~x18 && ~x14 && x15 && x13 )
						begin
							y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && ~x18 && ~x14 && x15 && ~x13 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && ~x18 && ~x14 && ~x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && ~x18 && ~x14 && ~x15 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && ~x18 && ~x14 && ~x15 && ~x2 && ~x3 && x13 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	
							nx_state = s361;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && x19 && ~x18 && ~x14 && ~x15 && ~x2 && ~x3 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && x13 && x20 && x14 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && x13 && x20 && ~x14 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && x13 && ~x20 && x15 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && x13 && ~x20 && ~x15 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && x14 && x20 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s288;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && x14 && ~x20 && x15 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && x14 && ~x20 && ~x15 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s288;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && ~x14 && x20 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && ~x14 && ~x20 && x15 && x6 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && ~x14 && ~x20 && x15 && ~x6 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && ~x14 && ~x20 && x15 && ~x6 && x4 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && ~x14 && ~x20 && x15 && ~x6 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && ~x14 && ~x20 && ~x15 && x5 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && ~x14 && ~x20 && ~x15 && ~x5 && x4 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && ~x14 && ~x20 && ~x15 && ~x5 && x4 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && x16 && ~x13 && ~x14 && ~x20 && ~x15 && ~x5 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && x20 && x14 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && x20 && x14 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && x20 && x14 && ~x2 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && x20 && ~x14 && x12 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && x20 && ~x14 && x12 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && x20 && ~x14 && x12 && ~x2 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && x20 && ~x14 && ~x12 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && x20 && ~x14 && ~x12 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && x20 && ~x14 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && x20 && ~x14 && ~x12 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && ~x20 && x15 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && ~x20 && ~x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && x13 && ~x20 && ~x15 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && x20 && x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && x20 && x11 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && x20 && x11 && ~x2 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && x20 && ~x11 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && x20 && ~x11 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && x20 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && x20 && ~x11 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && ~x20 && x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && ~x20 && x15 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && ~x20 && ~x15 && x12 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && ~x20 && ~x15 && x12 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && ~x20 && ~x15 && ~x12 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && ~x20 && ~x15 && ~x12 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && ~x20 && ~x15 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && x14 && ~x20 && ~x15 && ~x12 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && x20 && x10 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && x20 && x10 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && x20 && x10 && ~x2 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && x20 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && x20 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && x20 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && x20 && ~x10 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && x15 && x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && x15 && x11 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && x15 && ~x11 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && x15 && ~x11 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && x15 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && x15 && ~x11 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && ~x15 && x10 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && ~x15 && x10 && ~x2 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && ~x15 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && ~x15 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && ~x15 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x17 && ~x22 && ~x19 && ~x16 && ~x13 && ~x14 && ~x20 && ~x15 && ~x10 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && x18 && x19 && x10 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && x18 && x19 && ~x10 && x15 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && x18 && x19 && ~x10 && ~x15 )
						begin
							y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && x18 && ~x19 && x13 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && x18 && ~x19 && ~x13 && x15 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	
							nx_state = s361;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && x18 && ~x19 && ~x13 && ~x15 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && ~x18 && x19 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && ~x18 && x19 && ~x13 && x15 )
						begin
							y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && ~x18 && x19 && ~x13 && ~x15 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && ~x18 && ~x19 && x13 )
						begin
							y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && ~x18 && ~x19 && ~x13 && x15 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && x14 && ~x18 && ~x19 && ~x13 && ~x15 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && x15 && x19 && x18 && x10 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	
							nx_state = s361;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && x15 && x19 && x18 && ~x10 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && x15 && x19 && ~x18 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && x15 && x19 && ~x18 && ~x13 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && x15 && ~x19 && x13 )
						nx_state = s40;
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && x15 && ~x19 && ~x13 && x18 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && x15 && ~x19 && ~x13 && x18 && ~x3 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && x15 && ~x19 && ~x13 && ~x18 && x3 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	
							nx_state = s361;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && x15 && ~x19 && ~x13 && ~x18 && ~x3 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && x2 && x18 && x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && x2 && x18 && ~x19 && x13 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && x2 && x18 && ~x19 && ~x13 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s362;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && x2 && ~x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && x19 && x18 && x10 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && x19 && x18 && ~x10 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && x19 && ~x18 && x13 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	
							nx_state = s361;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && x19 && ~x18 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && ~x19 && x13 )
						begin
							y20 = 1'b1;	
							nx_state = s363;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && ~x19 && ~x13 && x18 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && ~x19 && ~x13 && ~x18 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s362;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && ~x16 && x18 && x19 && x10 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && ~x16 && x18 && x19 && ~x10 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && ~x16 && x18 && x19 && ~x10 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && ~x16 && x18 && x19 && ~x10 && ~x2 && ~x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s51;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && ~x16 && x18 && ~x19 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && ~x16 && x18 && ~x19 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && ~x16 && x18 && ~x19 && ~x2 && ~x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s51;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && ~x16 && ~x18 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && ~x16 && ~x18 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && x22 && ~x16 && ~x18 && ~x2 && ~x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s51;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && x15 && x13 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && x15 && ~x13 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && x15 && ~x13 && ~x2 && x14 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && x15 && ~x13 && ~x2 && x14 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && x15 && ~x13 && ~x2 && ~x14 && x11 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && x15 && ~x13 && ~x2 && ~x14 && x11 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && x15 && ~x13 && ~x2 && ~x14 && ~x11 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && x15 && ~x13 && ~x2 && ~x14 && ~x11 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && x15 && ~x13 && ~x2 && ~x14 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && x15 && ~x13 && ~x2 && ~x14 && ~x11 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && x13 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && x14 && x12 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && x14 && x12 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && x14 && ~x12 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && x14 && ~x12 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && x14 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && x14 && ~x12 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && ~x14 && x10 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && ~x14 && x10 && ~x3 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && ~x14 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && ~x14 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && ~x14 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && x18 && ~x15 && ~x2 && ~x13 && ~x14 && ~x10 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && ~x18 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && ~x18 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && x19 && ~x18 && ~x2 && ~x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s51;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && x14 && ~x13 && x15 && x20 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && x14 && ~x13 && x15 && ~x20 && x12 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && x14 && ~x13 && x15 && ~x20 && ~x12 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && x14 && ~x13 && ~x15 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s362;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && ~x14 && x15 && x20 && x13 )
						begin
							y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && ~x14 && x15 && x20 && ~x13 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && ~x14 && x15 && ~x20 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && ~x14 && x15 && ~x20 && ~x13 )
						begin
							y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && ~x14 && ~x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && ~x14 && ~x15 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && x13 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && x16 && ~x14 && ~x15 && ~x2 && ~x3 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s300;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && ~x16 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && ~x16 && ~x2 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	
							nx_state = s359;
						end
					else if( x65 && ~x66 && ~x21 && ~x17 && ~x22 && ~x19 && ~x16 && ~x2 && ~x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x65 && x21 && x68 && x16 && x17 && x10 && x15 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && x21 && x68 && x16 && x17 && x10 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x65 && x21 && x68 && x16 && x17 && ~x10 && x15 && x7 && x14 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s288;
						end
					else if( ~x65 && x21 && x68 && x16 && x17 && ~x10 && x15 && x7 && ~x14 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && x21 && x68 && x16 && x17 && ~x10 && x15 && ~x7 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x21 && x68 && x16 && x17 && ~x10 && x15 && ~x7 && x9 && ~x8 && x14 )
						nx_state = s86;
					else if( ~x65 && x21 && x68 && x16 && x17 && ~x10 && x15 && ~x7 && x9 && ~x8 && ~x14 )
						nx_state = s1;
					else if( ~x65 && x21 && x68 && x16 && x17 && ~x10 && x15 && ~x7 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x21 && x68 && x16 && x17 && ~x10 && ~x15 && x8 && x14 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s310;
						end
					else if( ~x65 && x21 && x68 && x16 && x17 && ~x10 && ~x15 && x8 && ~x14 )
						begin
							y5 = 1'b1;	
							nx_state = s305;
						end
					else if( ~x65 && x21 && x68 && x16 && x17 && ~x10 && ~x15 && ~x8 && x9 && x14 )
						nx_state = s86;
					else if( ~x65 && x21 && x68 && x16 && x17 && ~x10 && ~x15 && ~x8 && x9 && ~x14 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x21 && x68 && x16 && x17 && ~x10 && ~x15 && ~x8 && x9 && ~x14 && ~x7 )
						nx_state = s1;
					else if( ~x65 && x21 && x68 && x16 && x17 && ~x10 && ~x15 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x21 && x68 && x16 && ~x17 && x14 && x10 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x21 && x68 && x16 && ~x17 && x14 && ~x10 && x15 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x65 && x21 && x68 && x16 && ~x17 && x14 && ~x10 && x15 && ~x13 )
						begin
							y11 = 1'b1;	
							nx_state = s122;
						end
					else if( ~x65 && x21 && x68 && x16 && ~x17 && x14 && ~x10 && ~x15 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	
							nx_state = s221;
						end
					else if( ~x65 && x21 && x68 && x16 && ~x17 && ~x14 && x2 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s322;
						end
					else if( ~x65 && x21 && x68 && x16 && ~x17 && ~x14 && ~x2 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x21 && x68 && x16 && ~x17 && ~x14 && ~x2 && ~x4 && x15 && x10 )
						begin
							y11 = 1'b1;	
							nx_state = s357;
						end
					else if( ~x65 && x21 && x68 && x16 && ~x17 && ~x14 && ~x2 && ~x4 && x15 && ~x10 )
						begin
							y11 = 1'b1;	
							nx_state = s357;
						end
					else if( ~x65 && x21 && x68 && x16 && ~x17 && ~x14 && ~x2 && ~x4 && ~x15 && x10 )
						begin
							y2 = 1'b1;	y16 = 1'b1;	y24 = 1'b1;	
							nx_state = s124;
						end
					else if( ~x65 && x21 && x68 && x16 && ~x17 && ~x14 && ~x2 && ~x4 && ~x15 && ~x10 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x65 && x21 && x68 && ~x16 && x2 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s322;
						end
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && x10 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && x10 && ~x4 )
						begin
							y11 = 1'b1;	
							nx_state = s297;
						end
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && x15 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && x15 && ~x4 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && x13 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && x13 && ~x4 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && ~x13 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && ~x13 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && ~x13 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && x14 && ~x15 && ~x13 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && x12 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && x12 && ~x4 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && ~x12 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && ~x12 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && ~x12 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && x15 && ~x12 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && x11 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && x11 && ~x4 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && ~x11 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && ~x11 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && ~x11 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && x17 && ~x10 && ~x14 && ~x15 && ~x11 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && ~x17 && x4 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && ~x17 && ~x4 && x10 )
						begin
							y11 = 1'b1;	
							nx_state = s296;
						end
					else if( ~x65 && x21 && x68 && ~x16 && ~x2 && ~x17 && ~x4 && ~x10 )
						begin
							y11 = 1'b1;	
							nx_state = s356;
						end
					else if( ~x65 && x21 && ~x68 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s143;
						end
					else if( ~x65 && ~x21 && x22 && x68 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && ~x21 && x22 && x68 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && ~x21 && x22 && x68 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x68 && ~x7 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x68 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x21 && x22 && ~x68 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x21 && x22 && ~x68 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x68 && x23 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x68 && ~x23 && x18 && x14 )
						nx_state = s40;
					else if( ~x65 && ~x21 && x22 && ~x68 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s40;
					else if( ~x65 && ~x21 && x22 && ~x68 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x68 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x21 && ~x22 && x68 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && ~x21 && ~x22 && ~x68 && x23 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s330;
						end
					else if( ~x65 && ~x21 && ~x22 && ~x68 && ~x23 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s333;
						end
					else nx_state = s86;
				s87 : if( x21 && x19 && x15 && x10 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s330;
						end
					else if( x21 && x19 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x21 && x19 && x15 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s48;
						end
					else if( x21 && x19 && ~x15 && x16 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x21 && x19 && ~x15 && ~x16 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s340;
						end
					else if( x21 && ~x19 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s84;
						end
					else if( ~x21 && x23 )
						nx_state = s1;
					else if( ~x21 && ~x23 && x22 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s84;
						end
					else if( ~x21 && ~x23 && ~x22 )
						nx_state = s1;
					else nx_state = s87;
				s88 : if( x21 && x66 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x21 && x66 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x21 && x66 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x21 && x66 && ~x9 )
						nx_state = s1;
					else if( x21 && ~x66 && x19 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s272;
						end
					else if( x21 && ~x66 && x19 && ~x12 && x17 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s272;
						end
					else if( x21 && ~x66 && x19 && ~x12 && ~x17 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x21 && ~x66 && ~x19 && x20 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s272;
						end
					else if( x21 && ~x66 && ~x19 && x20 && ~x12 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x21 && ~x66 && ~x19 && ~x20 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s270;
						end
					else if( x21 && ~x66 && ~x19 && ~x20 && ~x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x21 && x66 )
						nx_state = s1;
					else if( ~x21 && ~x66 && x22 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x21 && ~x66 && ~x22 )
						nx_state = s1;
					else nx_state = s88;
				s89 : if( x66 && x65 && x61 && x60 )
						nx_state = s40;
					else if( x66 && x65 && x61 && ~x60 && x62 )
						nx_state = s1;
					else if( x66 && x65 && x61 && ~x60 && ~x62 && x15 && x12 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x66 && x65 && x61 && ~x60 && ~x62 && x15 && x12 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s250;
						end
					else if( x66 && x65 && x61 && ~x60 && ~x62 && x15 && ~x12 && x7 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x66 && x65 && x61 && ~x60 && ~x62 && x15 && ~x12 && ~x7 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s262;
						end
					else if( x66 && x65 && x61 && ~x60 && ~x62 && ~x15 && x16 && x7 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s251;
						end
					else if( x66 && x65 && x61 && ~x60 && ~x62 && ~x15 && x16 && x7 && ~x12 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s252;
						end
					else if( x66 && x65 && x61 && ~x60 && ~x62 && ~x15 && x16 && ~x7 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s252;
						end
					else if( x66 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x16 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s253;
						end
					else if( x66 && x65 && x61 && ~x60 && ~x62 && ~x15 && ~x16 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x66 && x65 && ~x61 && x60 && x15 && x12 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x66 && x65 && ~x61 && x60 && x15 && x12 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s250;
						end
					else if( x66 && x65 && ~x61 && x60 && x15 && ~x12 && x7 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x66 && x65 && ~x61 && x60 && x15 && ~x12 && ~x7 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s262;
						end
					else if( x66 && x65 && ~x61 && x60 && ~x15 && x16 && x7 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s251;
						end
					else if( x66 && x65 && ~x61 && x60 && ~x15 && x16 && x7 && ~x12 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s252;
						end
					else if( x66 && x65 && ~x61 && x60 && ~x15 && x16 && ~x7 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s252;
						end
					else if( x66 && x65 && ~x61 && x60 && ~x15 && ~x16 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s253;
						end
					else if( x66 && x65 && ~x61 && x60 && ~x15 && ~x16 && ~x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x66 && x65 && ~x61 && ~x60 && x62 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( x66 && x65 && ~x61 && ~x60 && ~x62 )
						nx_state = s40;
					else if( x66 && ~x65 && x67 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x66 && ~x65 && x67 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x66 && ~x65 && x67 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x66 && ~x65 && x67 && x62 && ~x61 )
						nx_state = s1;
					else if( x66 && ~x65 && x67 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && ~x65 && x67 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( x66 && ~x65 && x67 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && ~x65 && x67 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( x66 && ~x65 && x67 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x66 && ~x65 && x67 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( x66 && ~x65 && x67 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x66 && ~x65 && x67 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x66 && ~x65 && x67 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x66 && ~x65 && x67 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x66 && ~x65 && x67 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x66 && ~x65 && x67 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && x21 && x68 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x66 && ~x65 && ~x67 && x21 && x68 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x66 && ~x65 && ~x67 && x21 && x68 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && x21 && x68 && ~x9 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && x21 && ~x68 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x66 && ~x65 && ~x67 && x21 && ~x68 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x66 && ~x65 && ~x67 && x21 && ~x68 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && x21 && ~x68 && ~x18 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && x22 && x68 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && x22 && x68 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && x22 && x68 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && x22 && x68 && ~x7 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && x22 && ~x68 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && x22 && ~x68 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && x22 && ~x68 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && x22 && ~x68 && x23 && ~x17 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && x18 && x14 )
						nx_state = s40;
					else if( x66 && ~x65 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s40;
					else if( x66 && ~x65 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && ~x18 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x22 && x68 && ~x4 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x22 && ~x68 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x22 && ~x68 && ~x23 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x66 && x65 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x4 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && x24 && x26 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x66 && ~x65 && x67 && x24 && x26 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x66 && ~x65 && x67 && x24 && x26 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && x24 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x66 && ~x65 && x67 && x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x66 && ~x65 && x67 && x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && ~x24 && x25 && x26 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x66 && ~x65 && x67 && ~x24 && x25 && x26 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x66 && ~x65 && x67 && ~x24 && x25 && x26 && x19 && ~x14 && ~x13 )
						nx_state = s89;
					else if( ~x66 && ~x65 && x67 && ~x24 && x25 && x26 && ~x19 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && ~x24 && x25 && ~x26 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x67 && x21 && x19 && x17 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s272;
						end
					else if( ~x66 && ~x65 && ~x67 && x21 && x19 && x17 && ~x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s272;
						end
					else if( ~x66 && ~x65 && ~x67 && x21 && x19 && ~x17 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && ~x65 && ~x67 && x21 && x19 && ~x17 && ~x12 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x66 && ~x65 && ~x67 && x21 && ~x19 && x20 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s272;
						end
					else if( ~x66 && ~x65 && ~x67 && x21 && ~x19 && x20 && ~x12 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s105;
						end
					else if( ~x66 && ~x65 && ~x67 && x21 && ~x19 && ~x20 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s270;
						end
					else if( ~x66 && ~x65 && ~x67 && x21 && ~x19 && ~x20 && ~x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s109;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && x12 && x4 && x18 && x17 )
						begin
							y18 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && x12 && x4 && x18 && ~x17 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s275;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && x12 && x4 && ~x18 && x19 && x17 )
						begin
							y18 = 1'b1;	
							nx_state = s272;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && x12 && x4 && ~x18 && x19 && ~x17 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s275;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && x12 && x4 && ~x18 && ~x19 )
						begin
							y18 = 1'b1;	
							nx_state = s272;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && x12 && ~x4 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s275;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && x18 && x4 && x17 )
						begin
							y18 = 1'b1;	
							nx_state = s234;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && x18 && x4 && ~x17 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && x18 && ~x4 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s275;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && x17 && x14 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s275;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && x17 && ~x14 && x16 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s275;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && x17 && ~x14 && ~x16 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && x17 && ~x14 && ~x16 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && x17 && ~x14 && ~x16 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && x17 && ~x14 && ~x16 && ~x6 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && ~x17 && x16 && x15 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s275;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && ~x17 && x16 && ~x15 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && ~x17 && x16 && ~x15 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && ~x17 && x16 && ~x15 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && ~x17 && x16 && ~x15 && ~x6 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && ~x17 && ~x16 && x13 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && ~x17 && ~x16 && x13 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && ~x17 && ~x16 && x13 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && ~x17 && ~x16 && x13 && ~x6 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && x19 && ~x17 && ~x16 && ~x13 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s275;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && ~x19 && x4 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && x22 && ~x12 && ~x18 && ~x19 && ~x4 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s275;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && x15 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && ~x15 && x19 && x18 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && ~x15 && x19 && ~x18 )
						begin
							y5 = 1'b1;	
							nx_state = s342;
						end
					else if( ~x66 && ~x65 && ~x67 && ~x21 && ~x22 && ~x15 && ~x19 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else nx_state = s89;
				s90 : if( 1'b1 )
						begin
							y2 = 1'b1;	y21 = 1'b1;	
							nx_state = s364;
						end
					else nx_state = s90;
				s91 : if( x65 && x21 && x18 && x20 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( x65 && x21 && x18 && ~x20 )
						nx_state = s91;
					else if( x65 && x21 && ~x18 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x21 && x22 && x15 && x9 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x65 && ~x21 && x22 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x65 && ~x21 && x22 && ~x15 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s205;
						end
					else if( x65 && ~x21 && ~x22 && x23 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x21 && ~x22 && x23 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x21 && ~x22 && x23 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x22 && x23 && ~x20 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && x14 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && x68 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && x67 && x66 && x68 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && x67 && x66 && x68 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && x68 && x21 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && x68 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x65 && x67 && x66 && x68 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x65 && x67 && x66 && x68 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && x68 && ~x21 && ~x20 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && x14 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && x14 && ~x8 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && ~x14 && x7 && x8 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && ~x14 && x7 && ~x8 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && ~x14 && ~x7 && x8 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s65;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && x17 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && x17 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && ~x17 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && ~x14 && ~x7 && ~x8 && x13 )
						begin
							y3 = 1'b1;	
							nx_state = s65;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && x17 && x12 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && x17 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && ~x17 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && x2 && x8 && x7 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && x2 && x8 && ~x7 && x9 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && x2 && x8 && ~x7 && ~x9 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && x2 && ~x8 && x7 && x11 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && x2 && ~x8 && x7 && ~x11 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && x2 && ~x8 && ~x7 && x10 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && x2 && ~x8 && ~x7 && ~x10 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && x7 && x8 && x1 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && x7 && x8 && ~x1 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && x7 && ~x8 && x11 && x1 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && x7 && ~x8 && x11 && ~x1 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && x7 && ~x8 && ~x11 && x17 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && x7 && ~x8 && ~x11 && x17 && ~x13 && x12 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && x7 && ~x8 && ~x11 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && x7 && ~x8 && ~x11 && ~x17 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && x8 && x9 && x1 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && x8 && x9 && ~x1 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && x8 && ~x9 && x17 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && x8 && ~x9 && x17 && ~x13 && x12 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && x8 && ~x9 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && x8 && ~x9 && ~x17 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && ~x8 && x10 && x1 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && ~x8 && x10 && ~x1 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && ~x8 && ~x10 && x17 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && ~x8 && ~x10 && x17 && ~x13 && x12 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && ~x8 && ~x10 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && x16 && ~x15 && ~x2 && ~x7 && ~x8 && ~x10 && ~x17 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && ~x16 && x15 && x7 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s159;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && ~x16 && x15 && ~x7 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && ~x16 && x15 && ~x7 && ~x2 && x1 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && ~x16 && x15 && ~x7 && ~x2 && ~x1 && x8 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && ~x16 && x15 && ~x7 && ~x2 && ~x1 && ~x8 )
						begin
							y18 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && ~x16 && ~x15 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && ~x16 && ~x15 && ~x2 && x1 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && x64 && ~x16 && ~x15 && ~x2 && ~x1 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y28 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x65 && x67 && x66 && ~x68 && x63 && ~x64 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && x16 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && x16 && ~x8 && x6 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && x16 && ~x8 && ~x6 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && x8 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && x8 && ~x7 && x9 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && x8 && ~x7 && ~x9 && x19 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && x8 && ~x7 && ~x9 && x19 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && x8 && ~x7 && ~x9 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && x8 && ~x7 && ~x9 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && ~x8 && x7 && x11 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && ~x8 && x7 && ~x11 && x19 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && ~x8 && x7 && ~x11 && x19 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && ~x8 && x7 && ~x11 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && ~x8 && x7 && ~x11 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && ~x8 && ~x7 && x10 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && ~x8 && ~x7 && ~x10 && x19 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && ~x8 && ~x7 && ~x10 && x19 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && ~x8 && ~x7 && ~x10 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && x4 && ~x8 && ~x7 && ~x10 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && ~x4 && x6 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y28 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && x64 && ~x16 && ~x4 && ~x6 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && ~x64 && x19 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && ~x64 && x19 && ~x13 && x12 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && ~x64 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x67 && x66 && ~x68 && ~x63 && ~x64 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x67 && ~x66 && x24 && x26 && x16 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x67 && ~x66 && x24 && x26 && ~x16 && x17 && x13 && x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x67 && ~x66 && x24 && x26 && ~x16 && x17 && x13 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s282;
						end
					else if( ~x65 && x67 && ~x66 && x24 && x26 && ~x16 && x17 && x13 && ~x11 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x67 && ~x66 && x24 && x26 && ~x16 && x17 && ~x13 && x11 )
						begin
							y17 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x65 && x67 && ~x66 && x24 && x26 && ~x16 && x17 && ~x13 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x67 && ~x66 && x24 && x26 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x65 && x67 && ~x66 && x24 && ~x26 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x65 && x67 && ~x66 && ~x24 && x25 && x26 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && x67 && ~x66 && ~x24 && x25 && x26 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && x67 && ~x66 && ~x24 && x25 && x26 && x19 && ~x14 && ~x13 )
						nx_state = s91;
					else if( ~x65 && x67 && ~x66 && ~x24 && x25 && x26 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x67 && ~x66 && ~x24 && x25 && ~x26 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && x67 && ~x66 && ~x24 && ~x25 && x26 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else if( ~x65 && x67 && ~x66 && ~x24 && ~x25 && ~x26 && x15 && x12 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && x67 && ~x66 && ~x24 && ~x25 && ~x26 && x15 && ~x12 && x11 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && x67 && ~x66 && ~x24 && ~x25 && ~x26 && x15 && ~x12 && ~x11 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && x67 && ~x66 && ~x24 && ~x25 && ~x26 && x15 && ~x12 && ~x11 && ~x10 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x65 && x67 && ~x66 && ~x24 && ~x25 && ~x26 && ~x15 && x16 && x10 && x12 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s46;
						end
					else if( ~x65 && x67 && ~x66 && ~x24 && ~x25 && ~x26 && ~x15 && x16 && x10 && ~x12 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && x67 && ~x66 && ~x24 && ~x25 && ~x26 && ~x15 && x16 && ~x10 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s46;
						end
					else if( ~x65 && x67 && ~x66 && ~x24 && ~x25 && ~x26 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x67 && x66 && x21 )
						nx_state = s1;
					else if( ~x65 && ~x67 && x66 && ~x21 && x22 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && ~x67 && x66 && ~x21 && x22 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && ~x67 && x66 && ~x21 && x22 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x67 && x66 && ~x21 && x22 && ~x7 )
						nx_state = s1;
					else if( ~x65 && ~x67 && x66 && ~x21 && ~x22 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && ~x67 && x66 && ~x21 && ~x22 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && ~x67 && x66 && ~x21 && ~x22 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x66 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x65 && ~x67 && ~x66 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x65 && ~x67 && ~x66 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x66 && ~x3 )
						nx_state = s1;
					else nx_state = s91;
				s92 : if( x65 && x67 && x21 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s365;
						end
					else if( x65 && x67 && ~x21 && x23 && x22 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x21 && x23 && x22 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x21 && x23 && x22 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && x67 && ~x21 && x23 && x22 && ~x8 )
						nx_state = s1;
					else if( x65 && x67 && ~x21 && x23 && ~x22 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x21 && x23 && ~x22 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x21 && x23 && ~x22 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && x67 && ~x21 && x23 && ~x22 && ~x9 )
						nx_state = s1;
					else if( x65 && x67 && ~x21 && ~x23 && x8 && x22 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x21 && ~x23 && x8 && x22 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x21 && ~x23 && x8 && x22 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x65 && x67 && ~x21 && ~x23 && x8 && ~x22 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x21 && ~x23 && x8 && ~x22 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && ~x21 && ~x23 && x8 && ~x22 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && x67 && ~x21 && ~x23 && ~x8 )
						nx_state = s1;
					else if( x65 && ~x67 && x68 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x67 && x68 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x67 && x68 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x67 && x68 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x68 && x21 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && x23 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && x23 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && x23 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && x23 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && x23 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && x7 && x9 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && x7 && ~x9 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && ~x7 && x8 && x9 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s157;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && ~x7 && x8 && ~x9 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s158;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && ~x7 && ~x8 && x9 && x13 )
						begin
							y4 = 1'b1;	
							nx_state = s191;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && ~x7 && ~x8 && x9 && ~x13 && x18 && x14 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && ~x7 && ~x8 && x9 && ~x13 && x18 && ~x14 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && ~x7 && ~x8 && x9 && ~x13 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && ~x7 && ~x8 && ~x9 && x14 )
						begin
							y4 = 1'b1;	
							nx_state = s191;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && ~x7 && ~x8 && ~x9 && ~x14 && x18 && x13 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && ~x7 && ~x8 && ~x9 && ~x14 && x18 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && x16 && ~x7 && ~x8 && ~x9 && ~x14 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && ~x16 && x7 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && ~x16 && ~x7 && x8 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && ~x16 && ~x7 && ~x8 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s22;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && ~x16 && ~x7 && ~x8 && ~x1 && x5 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && ~x16 && ~x7 && ~x8 && ~x1 && ~x5 && x9 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && x15 && ~x16 && ~x7 && ~x8 && ~x1 && ~x5 && ~x9 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && x1 )
						begin
							y1 = 1'b1;	
							nx_state = s22;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && x9 && x10 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && x9 && ~x10 && x8 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && x9 && ~x10 && ~x8 && x18 && x14 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && x9 && ~x10 && ~x8 && x18 && ~x14 && x13 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && x9 && ~x10 && ~x8 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && x9 && ~x10 && ~x8 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && ~x9 && x8 && x12 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && ~x9 && x8 && ~x12 && x18 && x14 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && ~x9 && x8 && ~x12 && x18 && ~x14 && x13 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && ~x9 && x8 && ~x12 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && ~x9 && x8 && ~x12 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && ~x9 && ~x8 && x11 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && ~x9 && ~x8 && ~x11 && x18 && x14 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && ~x9 && ~x8 && ~x11 && x18 && ~x14 && x13 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && ~x9 && ~x8 && ~x11 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && x16 && ~x9 && ~x8 && ~x11 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && ~x16 && x5 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && x22 && ~x23 && ~x15 && ~x1 && ~x16 && ~x5 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s205;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && ~x22 && x4 && x18 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && ~x22 && x4 && ~x18 && x19 )
						nx_state = s92;
					else if( x65 && ~x67 && ~x68 && ~x21 && ~x22 && x4 && ~x18 && ~x19 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							nx_state = s97;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && ~x22 && ~x4 && x3 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && ~x67 && ~x68 && ~x21 && ~x22 && ~x4 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x65 && x66 && x68 && x21 )
						nx_state = s1;
					else if( ~x65 && x66 && x68 && ~x21 && x16 && x10 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s67;
						end
					else if( ~x65 && x66 && x68 && ~x21 && x16 && ~x10 )
						begin
							y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s113;
						end
					else if( ~x65 && x66 && x68 && ~x21 && ~x16 )
						begin
							y5 = 1'b1;	y17 = 1'b1;	
							nx_state = s115;
						end
					else if( ~x65 && x66 && ~x68 && x63 && x64 && x6 && x15 && x8 )
						begin
							y21 = 1'b1;	
							nx_state = s298;
						end
					else if( ~x65 && x66 && ~x68 && x63 && x64 && x6 && x15 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && x66 && ~x68 && x63 && x64 && x6 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s298;
						end
					else if( ~x65 && x66 && ~x68 && x63 && x64 && x6 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x65 && x66 && ~x68 && x63 && x64 && ~x6 )
						begin
							y21 = 1'b1;	
							nx_state = s298;
						end
					else if( ~x65 && x66 && ~x68 && x63 && ~x64 && x5 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s20;
						end
					else if( ~x65 && x66 && ~x68 && x63 && ~x64 && ~x5 && x18 && x15 && x8 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && x66 && ~x68 && x63 && ~x64 && ~x5 && x18 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x65 && x66 && ~x68 && x63 && ~x64 && ~x5 && x18 && ~x15 && x16 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x65 && x66 && ~x68 && x63 && ~x64 && ~x5 && x18 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x65 && x66 && ~x68 && x63 && ~x64 && ~x5 && ~x18 )
						begin
							y31 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x65 && x66 && ~x68 && ~x63 && x64 && x19 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x66 && ~x68 && ~x63 && x64 && x19 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x66 && ~x68 && ~x63 && x64 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x68 && ~x63 && x64 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x68 && ~x63 && ~x64 && x4 )
						begin
							y31 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x65 && x66 && ~x68 && ~x63 && ~x64 && ~x4 && x17 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x65 && x66 && ~x68 && ~x63 && ~x64 && ~x4 && x17 && x15 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && x66 && ~x68 && ~x63 && ~x64 && ~x4 && x17 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s151;
						end
					else if( ~x65 && x66 && ~x68 && ~x63 && ~x64 && ~x4 && x17 && ~x15 && ~x16 && x14 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x65 && x66 && ~x68 && ~x63 && ~x64 && ~x4 && x17 && ~x15 && ~x16 && ~x14 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s152;
						end
					else if( ~x65 && x66 && ~x68 && ~x63 && ~x64 && ~x4 && ~x17 )
						begin
							y14 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x65 && ~x66 && x67 && x68 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x66 && x67 && x68 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x66 && x67 && x68 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x68 && x20 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x68 && ~x20 && x21 && x3 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s366;
						end
					else if( ~x65 && ~x66 && x67 && x68 && ~x20 && x21 && ~x3 && x17 && x15 && x8 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x65 && ~x66 && x67 && x68 && ~x20 && x21 && ~x3 && x17 && x15 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x65 && ~x66 && x67 && x68 && ~x20 && x21 && ~x3 && x17 && ~x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x65 && ~x66 && x67 && x68 && ~x20 && x21 && ~x3 && x17 && ~x15 && ~x16 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s209;
						end
					else if( ~x65 && ~x66 && x67 && x68 && ~x20 && x21 && ~x3 && ~x17 )
						nx_state = s40;
					else if( ~x65 && ~x66 && x67 && x68 && ~x20 && ~x21 && x15 && x8 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x66 && x67 && x68 && ~x20 && ~x21 && x15 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x65 && ~x66 && x67 && x68 && ~x20 && ~x21 && ~x15 && x16 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x65 && ~x66 && x67 && x68 && ~x20 && ~x21 && ~x15 && ~x16 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s209;
						end
					else if( ~x65 && ~x66 && x67 && ~x68 && x24 && x26 && x16 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x66 && x67 && ~x68 && x24 && x26 && x16 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x66 && x67 && ~x68 && x24 && x26 && x16 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && ~x68 && x24 && x26 && x16 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && ~x68 && x24 && x26 && ~x16 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s165;
						end
					else if( ~x65 && ~x66 && x67 && ~x68 && x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && ~x66 && x67 && ~x68 && x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x65 && ~x66 && x67 && ~x68 && x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && ~x68 && x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && ~x68 && ~x24 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && x67 && ~x68 && ~x24 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && x67 && ~x68 && ~x24 && x25 && x19 && ~x14 && ~x13 && x26 )
						nx_state = s92;
					else if( ~x65 && ~x66 && x67 && ~x68 && ~x24 && x25 && x19 && ~x14 && ~x13 && ~x26 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && ~x68 && ~x24 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && ~x68 && ~x24 && ~x25 && x26 )
						begin
							y17 = 1'b1;	
							nx_state = s17;
						end
					else if( ~x65 && ~x66 && x67 && ~x68 && ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x65 && ~x66 && x67 && ~x68 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x65 && ~x66 && x67 && ~x68 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && ~x68 && ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && x68 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x65 && ~x66 && ~x67 && x68 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x65 && ~x66 && ~x67 && x68 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && x68 && ~x3 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x68 && x21 && x9 && x3 )
						nx_state = s40;
					else if( ~x65 && ~x66 && ~x67 && ~x68 && x21 && x9 && ~x3 && x4 )
						nx_state = s40;
					else if( ~x65 && ~x66 && ~x67 && ~x68 && x21 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x68 && x21 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x5 && ~x4 && x22 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x5 && ~x4 && x22 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && x5 && ~x4 && ~x22 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x5 && x22 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x5 && ~x22 && x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x5 && ~x22 && x4 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x68 && ~x21 && ~x5 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s92;
				s93 : if( x22 && x20 && x19 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s93;
						end
					else if( x22 && x20 && ~x19 && x23 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x22 && x20 && ~x19 && ~x23 )
						nx_state = s93;
					else if( x22 && ~x20 && x23 && x19 )
						nx_state = s93;
					else if( x22 && ~x20 && x23 && ~x19 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x22 && ~x20 && ~x23 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x22 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else nx_state = s93;
				s94 : if( x22 && x4 && x19 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s93;
						end
					else if( x22 && x4 && ~x19 && x20 )
						nx_state = s94;
					else if( x22 && x4 && ~x19 && ~x20 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x22 && ~x4 && x3 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x22 && ~x4 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else if( ~x22 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	y29 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s94;
				s95 : if( x21 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && x18 && x15 && x9 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x21 && x22 && x23 && x18 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x21 && x22 && x23 && x18 && ~x15 && x16 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x21 && x22 && x23 && x18 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x21 && x22 && x23 && ~x18 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							nx_state = s97;
						end
					else if( ~x21 && x22 && ~x23 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							nx_state = s97;
						end
					else if( ~x21 && ~x22 && x23 && x15 && x9 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x21 && ~x22 && x23 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x21 && ~x22 && x23 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && x23 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x21 && ~x22 && ~x23 )
						nx_state = s1;
					else nx_state = s95;
				s96 : if( x65 && x21 && x17 && x15 && x9 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( x65 && x21 && x17 && x15 && ~x9 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( x65 && x21 && x17 && ~x15 && x16 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x65 && x21 && x17 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s212;
						end
					else if( x65 && x21 && ~x17 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s294;
						end
					else if( x65 && ~x21 && x23 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s294;
						end
					else if( x65 && ~x21 && ~x23 && x22 && x5 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s294;
						end
					else if( x65 && ~x21 && ~x23 && x22 && ~x5 && x17 && x15 && x9 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x21 && ~x23 && x22 && ~x5 && x17 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x65 && ~x21 && ~x23 && x22 && ~x5 && x17 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && ~x23 && x22 && ~x5 && x17 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s205;
						end
					else if( x65 && ~x21 && ~x23 && x22 && ~x5 && ~x17 )
						begin
							y35 = 1'b1;	
							nx_state = s26;
						end
					else if( x65 && ~x21 && ~x23 && ~x22 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x65 && x63 )
						begin
							y14 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x65 && ~x63 && x64 && x18 && x16 && x8 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && ~x63 && x64 && x18 && x16 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x63 && x64 && x18 && ~x16 && x4 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x65 && ~x63 && x64 && x18 && ~x16 && ~x4 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x65 && ~x63 && x64 && ~x18 )
						begin
							y14 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x65 && ~x63 && ~x64 && x17 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x65 && ~x63 && ~x64 && x17 && x15 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x63 && ~x64 && x17 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s151;
						end
					else if( ~x65 && ~x63 && ~x64 && x17 && ~x15 && ~x16 && x14 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x65 && ~x63 && ~x64 && x17 && ~x15 && ~x16 && ~x14 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s152;
						end
					else if( ~x65 && ~x63 && ~x64 && ~x17 )
						begin
							y14 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s18;
						end
					else nx_state = s96;
				s97 : if( x23 && x22 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s98;
						end
					else if( x23 && ~x22 )
						nx_state = s1;
					else if( ~x23 && x22 )
						begin
							y21 = 1'b1;	
							nx_state = s298;
						end
					else if( ~x23 && ~x22 && x4 && x20 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s98;
						end
					else if( ~x23 && ~x22 && x4 && ~x20 && x19 )
						nx_state = s97;
					else if( ~x23 && ~x22 && x4 && ~x20 && ~x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( ~x23 && ~x22 && ~x4 && x3 )
						begin
							y1 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s93;
						end
					else if( ~x23 && ~x22 && ~x4 && ~x3 )
						begin
							y1 = 1'b1;	
							nx_state = s24;
						end
					else nx_state = s97;
				s98 : if( x22 && x15 && x9 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x22 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x22 && ~x15 && x16 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x22 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x22 && x19 && x20 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s98;
						end
					else if( ~x22 && x19 && ~x20 )
						nx_state = s98;
					else if( ~x22 && ~x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else nx_state = s98;
				s99 : if( x23 && x22 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x23 && x22 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x23 && x22 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x23 && x22 && ~x17 )
						nx_state = s1;
					else if( x23 && ~x22 )
						nx_state = s1;
					else if( ~x23 )
						nx_state = s1;
					else nx_state = s99;
				s100 : if( x65 && x66 && x67 && x23 && x18 && x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && x66 && x67 && x23 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && x66 && x67 && x23 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && x66 && x67 && x23 && ~x18 )
						nx_state = s1;
					else if( x65 && x66 && x67 && ~x23 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x65 && x66 && ~x67 && x61 && x60 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x66 && ~x67 && x61 && x60 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x66 && ~x67 && x61 && x60 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x66 && ~x67 && x61 && x60 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x66 && ~x67 && x61 && ~x60 && x62 && x2 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x65 && x66 && ~x67 && x61 && ~x60 && x62 && ~x2 && x20 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	
							nx_state = s367;
						end
					else if( x65 && x66 && ~x67 && x61 && ~x60 && x62 && ~x2 && ~x20 && x16 && x11 && x12 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x65 && x66 && ~x67 && x61 && ~x60 && x62 && ~x2 && ~x20 && x16 && x11 && ~x12 && x13 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x65 && x66 && ~x67 && x61 && ~x60 && x62 && ~x2 && ~x20 && x16 && x11 && ~x12 && ~x13 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s154;
						end
					else if( x65 && x66 && ~x67 && x61 && ~x60 && x62 && ~x2 && ~x20 && x16 && ~x11 && x13 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s63;
						end
					else if( x65 && x66 && ~x67 && x61 && ~x60 && x62 && ~x2 && ~x20 && x16 && ~x11 && ~x13 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( x65 && x66 && ~x67 && x61 && ~x60 && x62 && ~x2 && ~x20 && ~x16 && x17 && x11 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x65 && x66 && ~x67 && x61 && ~x60 && x62 && ~x2 && ~x20 && ~x16 && x17 && x11 && ~x13 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( x65 && x66 && ~x67 && x61 && ~x60 && x62 && ~x2 && ~x20 && ~x16 && x17 && ~x11 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x65 && x66 && ~x67 && x61 && ~x60 && x62 && ~x2 && ~x20 && ~x16 && ~x17 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( x65 && x66 && ~x67 && x61 && ~x60 && ~x62 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x65 && x66 && ~x67 && x61 && ~x60 && ~x62 && ~x7 )
						nx_state = s39;
					else if( x65 && x66 && ~x67 && ~x61 && x60 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x65 && x66 && ~x67 && ~x61 && x60 && ~x7 )
						nx_state = s39;
					else if( x65 && x66 && ~x67 && ~x61 && ~x60 && x62 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( x65 && x66 && ~x67 && ~x61 && ~x60 && ~x62 )
						nx_state = s316;
					else if( x65 && ~x66 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x65 && ~x66 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && x15 && x9 )
						begin
							y31 = 1'b1;	
							nx_state = s96;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x15 && ~x9 && x6 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x15 && ~x9 && ~x6 )
						begin
							y31 = 1'b1;	
							nx_state = s96;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && x9 && x8 )
						begin
							y31 = 1'b1;	
							nx_state = s96;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && x9 && ~x8 && x10 )
						begin
							y31 = 1'b1;	
							nx_state = s96;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && x9 && ~x8 && ~x10 && x18 && x14 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && x9 && ~x8 && ~x10 && x18 && ~x14 && x13 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && x9 && ~x8 && ~x10 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && x9 && ~x8 && ~x10 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && ~x9 && x8 && x12 )
						begin
							y31 = 1'b1;	
							nx_state = s96;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && ~x9 && x8 && ~x12 && x18 && x14 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && ~x9 && x8 && ~x12 && x18 && ~x14 && x13 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && ~x9 && x8 && ~x12 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && ~x9 && x8 && ~x12 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && ~x9 && ~x8 && x11 )
						begin
							y31 = 1'b1;	
							nx_state = s96;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && ~x9 && ~x8 && ~x11 && x18 && x14 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && ~x9 && ~x8 && ~x11 && x18 && ~x14 && x13 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && ~x9 && ~x8 && ~x11 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x15 && x16 && ~x9 && ~x8 && ~x11 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x15 && ~x16 && x6 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s212;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x15 && ~x16 && ~x6 )
						begin
							y31 = 1'b1;	
							nx_state = s96;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 )
						begin
							y31 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x65 && x66 && x21 && x68 )
						nx_state = s1;
					else if( ~x65 && x66 && x21 && ~x68 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x65 && x66 && x21 && ~x68 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x65 && x66 && x21 && ~x68 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x66 && x21 && ~x68 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x21 && x22 && x68 && x17 && x10 && x15 && x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x65 && x66 && ~x21 && x22 && x68 && x17 && x10 && x15 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && x66 && ~x21 && x22 && x68 && x17 && x10 && ~x15 && x16 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x65 && x66 && ~x21 && x22 && x68 && x17 && x10 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && x66 && ~x21 && x22 && x68 && x17 && ~x10 && x6 )
						begin
							y13 = 1'b1;	y16 = 1'b1;	
							nx_state = s284;
						end
					else if( ~x65 && x66 && ~x21 && x22 && x68 && x17 && ~x10 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && x66 && ~x21 && x22 && x68 && ~x17 && x18 && x6 && x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s219;
						end
					else if( ~x65 && x66 && ~x21 && x22 && x68 && ~x17 && x18 && x6 && ~x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x65 && x66 && ~x21 && x22 && x68 && ~x17 && x18 && ~x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && x66 && ~x21 && x22 && x68 && ~x17 && ~x18 && x6 && x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s219;
						end
					else if( ~x65 && x66 && ~x21 && x22 && x68 && ~x17 && ~x18 && x6 && ~x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s28;
						end
					else if( ~x65 && x66 && ~x21 && x22 && x68 && ~x17 && ~x18 && ~x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x66 && ~x21 && x22 && ~x68 && x23 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x65 && x66 && ~x21 && x22 && ~x68 && ~x23 && x18 && x14 )
						nx_state = s40;
					else if( ~x65 && x66 && ~x21 && x22 && ~x68 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s40;
					else if( ~x65 && x66 && ~x21 && x22 && ~x68 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x21 && x22 && ~x68 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x21 && ~x22 && x68 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && x68 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && x68 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x21 && ~x22 && x68 && ~x4 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x21 && ~x22 && ~x68 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x66 && x67 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x66 && x67 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x20 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && ~x20 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x65 && ~x66 && ~x67 && x21 && x9 && x3 )
						nx_state = s40;
					else if( ~x65 && ~x66 && ~x67 && x21 && x9 && ~x3 && x4 )
						nx_state = s40;
					else if( ~x65 && ~x66 && ~x67 && x21 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && x21 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && ~x5 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x21 && ~x22 )
						nx_state = s1;
					else nx_state = s100;
				s101 : if( x65 && x66 && x22 && x20 && x15 && x8 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x66 && x22 && x20 && x15 && ~x8 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x65 && x66 && x22 && x20 && ~x15 && x16 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s302;
						end
					else if( x65 && x66 && x22 && x20 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s122;
						end
					else if( x65 && x66 && x22 && ~x20 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s368;
						end
					else if( x65 && x66 && ~x22 && x23 )
						nx_state = s1;
					else if( x65 && x66 && ~x22 && ~x23 && x3 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s368;
						end
					else if( x65 && x66 && ~x22 && ~x23 && ~x3 && x19 && x15 && x8 )
						begin
							y11 = 1'b1;	
							nx_state = s8;
						end
					else if( x65 && x66 && ~x22 && ~x23 && ~x3 && x19 && x15 && ~x8 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s111;
						end
					else if( x65 && x66 && ~x22 && ~x23 && ~x3 && x19 && ~x15 && x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x66 && ~x22 && ~x23 && ~x3 && x19 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( x65 && x66 && ~x22 && ~x23 && ~x3 && ~x19 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s314;
						end
					else if( x65 && ~x66 && x68 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x68 && x21 && x5 )
						begin
							y31 = 1'b1;	
							nx_state = s96;
						end
					else if( x65 && ~x66 && ~x68 && x21 && ~x5 && x17 && x15 && x9 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( x65 && ~x66 && ~x68 && x21 && ~x5 && x17 && x15 && ~x9 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( x65 && ~x66 && ~x68 && x21 && ~x5 && x17 && ~x15 && x16 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x65 && ~x66 && ~x68 && x21 && ~x5 && x17 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s212;
						end
					else if( x65 && ~x66 && ~x68 && x21 && ~x5 && ~x17 )
						begin
							y15 = 1'b1;	y32 = 1'b1;	y33 = 1'b1;	
							y34 = 1'b1;	
							nx_state = s294;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && x15 && x9 && x23 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && x15 && x9 && ~x23 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && x15 && ~x9 && x23 && x6 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && x15 && ~x9 && x23 && ~x6 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && x15 && ~x9 && ~x23 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && x9 && x8 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && x9 && ~x8 && x10 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && x9 && ~x8 && ~x10 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && x9 && ~x8 && ~x10 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && x9 && ~x8 && ~x10 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && x9 && ~x8 && ~x10 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && x9 && ~x8 && ~x10 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && x8 && x12 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && x8 && ~x12 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && x8 && ~x12 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && x8 && ~x12 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && x8 && ~x12 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && x8 && ~x12 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && ~x8 && x11 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && ~x8 && ~x11 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && ~x8 && ~x11 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && ~x8 && ~x11 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && ~x8 && ~x11 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && x16 && ~x9 && ~x8 && ~x11 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && ~x16 && x6 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s205;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && x23 && ~x16 && ~x6 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && x22 && ~x15 && ~x23 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s205;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && ~x22 && x23 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && ~x22 && x23 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && ~x22 && x23 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x68 && ~x21 && ~x22 && x23 && ~x20 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x68 && ~x21 && ~x22 && ~x23 && x18 && x14 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && ~x22 && ~x23 && x18 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x66 && ~x68 && ~x21 && ~x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x68 && ~x21 && ~x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && x62 && x6 && x15 && x8 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s369;
						end
					else if( ~x65 && x66 && x67 && x62 && x6 && x15 && ~x8 )
						begin
							y18 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x65 && x66 && x67 && x62 && x6 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s369;
						end
					else if( ~x65 && x66 && x67 && x62 && x6 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x65 && x66 && x67 && x62 && ~x6 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s369;
						end
					else if( ~x65 && x66 && x67 && ~x62 && x63 && x17 && x13 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && x66 && x67 && ~x62 && x63 && x17 && ~x13 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && x66 && x67 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && x14 && x8 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && x14 && ~x8 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && ~x14 && x7 && x8 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && ~x14 && x7 && ~x8 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s158;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && ~x14 && ~x7 && x8 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s65;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && ~x14 && ~x7 && x8 && ~x12 && x19 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && ~x14 && ~x7 && x8 && ~x12 && x19 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && ~x14 && ~x7 && x8 && ~x12 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && ~x14 && ~x7 && ~x8 && x13 )
						begin
							y3 = 1'b1;	
							nx_state = s65;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && ~x14 && ~x7 && ~x8 && ~x13 && x19 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && ~x14 && ~x7 && ~x8 && ~x13 && x19 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && x4 && ~x14 && ~x7 && ~x8 && ~x13 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && ~x4 && x7 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s159;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && ~x4 && ~x7 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s190;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && ~x4 && ~x7 && ~x3 && x8 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && x16 && ~x4 && ~x7 && ~x3 && ~x8 )
						begin
							y18 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && x3 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s190;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && x7 && x11 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && x7 && ~x11 && x8 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && x7 && ~x11 && ~x8 && x19 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && x7 && ~x11 && ~x8 && x19 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && x7 && ~x11 && ~x8 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && x7 && ~x11 && ~x8 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && ~x7 && x8 && x9 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && ~x7 && x8 && ~x9 && x19 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && ~x7 && x8 && ~x9 && x19 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && ~x7 && x8 && ~x9 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && ~x7 && x8 && ~x9 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && ~x7 && ~x8 && x10 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && ~x7 && ~x8 && ~x10 && x19 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && ~x7 && ~x8 && ~x10 && x19 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && ~x7 && ~x8 && ~x10 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && x4 && ~x7 && ~x8 && ~x10 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && ~x4 && x15 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && x64 && ~x16 && ~x3 && ~x4 && ~x15 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y30 = 1'b1;	
							nx_state = s204;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && ~x64 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && ~x64 && x15 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && ~x64 && ~x15 && x16 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && ~x64 && ~x15 && ~x16 && x14 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x65 && x66 && x67 && ~x62 && ~x63 && ~x64 && ~x15 && ~x16 && ~x14 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s152;
						end
					else if( ~x65 && x66 && ~x67 && x21 && x68 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x66 && ~x67 && x21 && x68 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x66 && ~x67 && x21 && x68 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && x21 && x68 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && x21 && ~x68 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x65 && x66 && ~x67 && x21 && ~x68 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x65 && x66 && ~x67 && x21 && ~x68 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && x21 && ~x68 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && x68 && x17 && x10 && x15 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && x68 && x17 && x10 && ~x15 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && x68 && x17 && ~x10 )
						begin
							y13 = 1'b1;	y16 = 1'b1;	
							nx_state = s284;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && x68 && ~x17 && x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s219;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && x68 && ~x17 && ~x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && x23 && ~x17 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && x10 && x12 && x18 && x14 )
						nx_state = s40;
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && x10 && x12 && x18 && ~x14 && x13 )
						nx_state = s40;
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && x10 && x12 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && x10 && x12 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && x10 && ~x12 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && ~x10 && x18 && x14 )
						nx_state = s40;
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && ~x10 && x18 && ~x14 && x13 )
						nx_state = s40;
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && ~x10 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && ~x21 && x22 && ~x68 && ~x23 && ~x10 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && ~x21 && ~x22 && x68 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x67 && ~x21 && ~x22 && ~x68 && x23 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s180;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x23 && x15 && x9 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s370;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x23 && x15 && ~x9 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x23 && ~x15 && x16 && x7 && x9 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s330;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x23 && ~x15 && x16 && x7 && ~x9 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s333;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x23 && ~x15 && x16 && ~x7 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s330;
						end
					else if( ~x65 && x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x23 && ~x15 && ~x16 )
						begin
							y14 = 1'b1;	
							nx_state = s285;
						end
					else if( ~x65 && ~x66 && x21 && x68 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	
							nx_state = s142;
						end
					else if( ~x65 && ~x66 && x21 && ~x68 && x19 && x13 && x20 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && ~x66 && x21 && ~x68 && x19 && x13 && x20 && ~x15 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && ~x66 && x21 && ~x68 && x19 && x13 && ~x20 )
						begin
							y2 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s371;
						end
					else if( ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && x20 && x14 && x15 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && x20 && x14 && ~x15 )
						begin
							y22 = 1'b1;	y25 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && x20 && ~x14 && x15 && x4 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s372;
						end
					else if( ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && x20 && ~x14 && x15 && ~x4 && x9 && x3 )
						nx_state = s40;
					else if( ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && x20 && ~x14 && x15 && ~x4 && x9 && ~x3 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && x20 && ~x14 && x15 && ~x4 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && x20 && ~x14 && ~x15 && x3 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s372;
						end
					else if( ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && x20 && ~x14 && ~x15 && ~x3 && x9 && x4 )
						nx_state = s40;
					else if( ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && x20 && ~x14 && ~x15 && ~x3 && x9 && ~x4 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && x20 && ~x14 && ~x15 && ~x3 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && ~x20 && x14 )
						begin
							y2 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s371;
						end
					else if( ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && ~x20 && ~x14 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s328;
						end
					else if( ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && ~x20 && ~x14 && ~x5 && x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y9 = 1'b1;	
							nx_state = s107;
						end
					else if( ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && ~x20 && ~x14 && ~x5 && ~x6 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x66 && x21 && ~x68 && x19 && ~x13 && ~x20 && ~x14 && ~x5 && ~x6 && ~x15 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x66 && x21 && ~x68 && ~x19 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s328;
						end
					else if( ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && x14 && x18 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && x14 && ~x18 && x15 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && x14 && ~x18 && ~x15 && x9 && x3 )
						nx_state = s40;
					else if( ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && x14 && ~x18 && ~x15 && x9 && ~x3 && x4 )
						nx_state = s40;
					else if( ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && x14 && ~x18 && ~x15 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && x14 && ~x18 && ~x15 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && ~x14 && x15 && x16 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && ~x14 && x15 && ~x16 && x9 && x3 )
						nx_state = s40;
					else if( ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && ~x14 && x15 && ~x16 && x9 && ~x3 && x4 )
						nx_state = s40;
					else if( ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && ~x14 && x15 && ~x16 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && ~x14 && x15 && ~x16 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && ~x14 && ~x15 && x17 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && ~x14 && ~x15 && ~x17 && x9 && x3 )
						nx_state = s40;
					else if( ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && ~x14 && ~x15 && ~x17 && x9 && ~x3 && x4 )
						nx_state = s40;
					else if( ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && ~x14 && ~x15 && ~x17 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && x20 && ~x14 && ~x15 && ~x17 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && ~x20 && x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y9 = 1'b1;	
							nx_state = s107;
						end
					else if( ~x65 && ~x66 && x21 && ~x68 && ~x19 && ~x5 && ~x20 && ~x6 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	y23 = 1'b1;	
							nx_state = s373;
						end
					else if( ~x65 && ~x66 && ~x21 && x68 && x22 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x65 && ~x66 && ~x21 && x68 && x22 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x65 && ~x66 && ~x21 && x68 && x22 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x21 && x68 && x22 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x21 && x68 && ~x22 && x15 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	
							nx_state = s142;
						end
					else if( ~x65 && ~x66 && ~x21 && x68 && ~x22 && ~x15 && x19 && x18 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	
							nx_state = s142;
						end
					else if( ~x65 && ~x66 && ~x21 && x68 && ~x22 && ~x15 && x19 && ~x18 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && ~x66 && ~x21 && x68 && ~x22 && ~x15 && x19 && ~x18 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && ~x66 && ~x21 && x68 && ~x22 && ~x15 && x19 && ~x18 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x21 && x68 && ~x22 && ~x15 && x19 && ~x18 && ~x8 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x21 && x68 && ~x22 && ~x15 && ~x19 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	
							nx_state = s142;
						end
					else if( ~x65 && ~x66 && ~x21 && ~x68 && x22 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x65 && ~x66 && ~x21 && ~x68 && ~x22 && x9 && x11 )
						nx_state = s40;
					else if( ~x65 && ~x66 && ~x21 && ~x68 && ~x22 && x9 && ~x11 && x2 )
						nx_state = s101;
					else if( ~x65 && ~x66 && ~x21 && ~x68 && ~x22 && x9 && ~x11 && ~x2 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x65 && ~x66 && ~x21 && ~x68 && ~x22 && ~x9 && x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s108;
						end
					else if( ~x65 && ~x66 && ~x21 && ~x68 && ~x22 && ~x9 && ~x8 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else nx_state = s101;
				s102 : if( x65 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x5 )
						nx_state = s1;
					else if( ~x65 && x21 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x16 && x12 && x19 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x16 && x12 && ~x19 && x18 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x65 && ~x21 && x22 && x16 && x12 && ~x19 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x16 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x16 )
						nx_state = s1;
					else if( ~x65 && ~x21 && ~x22 && x18 && x15 )
						begin
							y8 = 1'b1;	y18 = 1'b1;	
							nx_state = s82;
						end
					else if( ~x65 && ~x21 && ~x22 && x18 && ~x15 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s374;
						end
					else if( ~x65 && ~x21 && ~x22 && ~x18 && x19 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s320;
						end
					else if( ~x65 && ~x21 && ~x22 && ~x18 && x19 && ~x15 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && ~x21 && ~x22 && ~x18 && ~x19 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else nx_state = s102;
				s103 : if( x21 && x12 && x11 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( x21 && x12 && ~x11 && x10 )
						nx_state = s103;
					else if( x21 && x12 && ~x11 && ~x10 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s104;
						end
					else if( x21 && ~x12 && x2 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( x21 && ~x12 && ~x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x21 && x22 && x19 && x15 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y17 = 1'b1;	
							nx_state = s177;
						end
					else if( ~x21 && x22 && x19 && ~x15 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x21 && x22 && ~x19 && x20 && x14 && x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && x22 && ~x19 && x20 && x14 && ~x18 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && ~x19 && x20 && x14 && ~x18 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && ~x19 && x20 && x14 && ~x18 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x20 && x14 && ~x18 && ~x5 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x20 && ~x14 && x15 && x16 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x14 && x15 && ~x16 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x14 && x15 && ~x16 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x14 && x15 && ~x16 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x20 && ~x14 && x15 && ~x16 && ~x5 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x20 && ~x14 && ~x15 && x17 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x14 && ~x15 && ~x17 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x14 && ~x15 && ~x17 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x14 && ~x15 && ~x17 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x20 && ~x14 && ~x15 && ~x17 && ~x5 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && ~x20 )
						begin
							y21 = 1'b1;	
							nx_state = s151;
						end
					else if( ~x21 && ~x22 && x7 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x21 && ~x22 && ~x7 && x10 && x19 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x21 && ~x22 && ~x7 && x10 && x19 && ~x15 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x21 && ~x22 && ~x7 && x10 && ~x19 && x20 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x21 && ~x22 && ~x7 && x10 && ~x19 && ~x20 )
						begin
							y21 = 1'b1;	
							nx_state = s151;
						end
					else if( ~x21 && ~x22 && ~x7 && ~x10 )
						begin
							y10 = 1'b1;	y17 = 1'b1;	y20 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s104;
						end
					else nx_state = s103;
				s104 : if( x21 )
						nx_state = s1;
					else if( ~x21 && x22 && x19 && x15 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y17 = 1'b1;	
							nx_state = s177;
						end
					else if( ~x21 && x22 && x19 && ~x15 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x21 && x22 && ~x19 && x20 && x15 && x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && x22 && ~x19 && x20 && x15 && ~x14 && x16 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && x22 && ~x19 && x20 && x15 && ~x14 && ~x16 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && ~x19 && x20 && x15 && ~x14 && ~x16 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && ~x19 && x20 && x15 && ~x14 && ~x16 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x20 && x15 && ~x14 && ~x16 && ~x5 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x20 && ~x15 && x14 && x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x15 && x14 && ~x18 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x15 && x14 && ~x18 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x15 && x14 && ~x18 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x20 && ~x15 && x14 && ~x18 && ~x5 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x20 && ~x15 && ~x14 && x17 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && ~x5 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && ~x20 )
						begin
							y21 = 1'b1;	
							nx_state = s151;
						end
					else if( ~x21 && ~x22 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s176;
						end
					else nx_state = s104;
				s105 : if( x21 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( x21 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( x21 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x21 && ~x3 )
						nx_state = s1;
					else if( ~x21 && x22 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s375;
						end
					else if( ~x21 && ~x22 && x18 && x15 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s375;
						end
					else if( ~x21 && ~x22 && x18 && ~x15 && x4 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x21 && ~x22 && x18 && ~x15 && ~x4 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s375;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && x15 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s375;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && x17 && x13 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s375;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && x17 && ~x13 && x16 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s375;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && x17 && ~x13 && ~x16 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && x17 && ~x13 && ~x16 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && x17 && ~x13 && ~x16 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && x17 && ~x13 && ~x16 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && ~x17 && x16 && x14 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s375;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && ~x17 && x16 && ~x14 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && ~x17 && x16 && ~x14 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && ~x17 && x16 && ~x14 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && ~x17 && x16 && ~x14 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && x12 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s375;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && ~x12 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && ~x12 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && ~x12 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 && ~x17 && ~x16 && ~x12 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x18 && ~x19 && x4 )
						begin
							y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s376;
						end
					else if( ~x21 && ~x22 && ~x18 && ~x19 && ~x4 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s375;
						end
					else nx_state = s105;
				s106 : if( x21 && x8 && x19 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( x21 && x8 && ~x19 && x20 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s176;
						end
					else if( x21 && x8 && ~x19 && ~x20 )
						begin
							y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s377;
						end
					else if( x21 && ~x8 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	
							nx_state = s378;
						end
					else if( ~x21 && x22 && x11 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y9 = 1'b1;	
							nx_state = s107;
						end
					else if( ~x21 && x22 && x11 && ~x2 )
						nx_state = s40;
					else if( ~x21 && x22 && ~x11 && x9 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( ~x21 && x22 && ~x11 && ~x9 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x21 && ~x22 )
						nx_state = s1;
					else nx_state = s106;
				s107 : if( x21 && x19 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( x21 && ~x19 )
						begin
							y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s377;
						end
					else if( ~x21 && x22 && x3 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y9 = 1'b1;	
							nx_state = s107;
						end
					else if( ~x21 && x22 && x3 && ~x2 )
						nx_state = s40;
					else if( ~x21 && x22 && ~x3 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x21 && ~x22 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s379;
						end
					else nx_state = s107;
				s108 : if( x21 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s380;
						end
					else if( ~x21 && x22 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x21 && ~x22 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y9 = 1'b1;	
							nx_state = s107;
						end
					else nx_state = s108;
				s109 : if( x21 )
						begin
							y18 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x21 && x22 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x21 && x22 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x21 && x22 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 )
						nx_state = s1;
					else nx_state = s109;
				s110 : if( x66 && x21 && x5 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( x66 && x21 && ~x5 && x19 && x15 && x10 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s330;
						end
					else if( x66 && x21 && ~x5 && x19 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x66 && x21 && ~x5 && x19 && x15 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s48;
						end
					else if( x66 && x21 && ~x5 && x19 && ~x15 && x16 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x66 && x21 && ~x5 && x19 && ~x15 && ~x16 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s340;
						end
					else if( x66 && x21 && ~x5 && ~x19 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s84;
						end
					else if( x66 && ~x21 && x22 && x23 && x3 && x15 && x10 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s339;
						end
					else if( x66 && ~x21 && x22 && x23 && x3 && x15 && ~x10 && x12 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s126;
						end
					else if( x66 && ~x21 && x22 && x23 && x3 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( x66 && ~x21 && x22 && x23 && x3 && ~x15 && x16 && x10 && x12 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s370;
						end
					else if( x66 && ~x21 && x22 && x23 && x3 && ~x15 && x16 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s381;
						end
					else if( x66 && ~x21 && x22 && x23 && x3 && ~x15 && x16 && ~x10 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s370;
						end
					else if( x66 && ~x21 && x22 && x23 && x3 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s180;
						end
					else if( x66 && ~x21 && x22 && x23 && ~x3 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s339;
						end
					else if( x66 && ~x21 && x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x66 && ~x21 && ~x22 && x15 && x4 && x7 )
						nx_state = s40;
					else if( x66 && ~x21 && ~x22 && x15 && x4 && ~x7 && x23 && x9 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s370;
						end
					else if( x66 && ~x21 && ~x22 && x15 && x4 && ~x7 && x23 && ~x9 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( x66 && ~x21 && ~x22 && x15 && x4 && ~x7 && ~x23 && x9 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s341;
						end
					else if( x66 && ~x21 && ~x22 && x15 && x4 && ~x7 && ~x23 && ~x9 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s339;
						end
					else if( x66 && ~x21 && ~x22 && x15 && ~x4 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x66 && ~x21 && ~x22 && ~x15 && x16 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x66 && ~x21 && ~x22 && ~x15 && ~x16 && x23 && x4 )
						begin
							y14 = 1'b1;	
							nx_state = s285;
						end
					else if( x66 && ~x21 && ~x22 && ~x15 && ~x16 && x23 && ~x4 )
						begin
							y14 = 1'b1;	
							nx_state = s48;
						end
					else if( x66 && ~x21 && ~x22 && ~x15 && ~x16 && ~x23 && x4 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s336;
						end
					else if( x66 && ~x21 && ~x22 && ~x15 && ~x16 && ~x23 && ~x4 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x66 && x67 && x24 && x26 && x20 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x66 && x67 && x24 && x26 && ~x20 && x21 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x66 && x67 && x24 && x26 && ~x20 && ~x21 && x22 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x66 && x67 && x24 && x26 && ~x20 && ~x21 && ~x22 && x23 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x66 && x67 && x24 && x26 && ~x20 && ~x21 && ~x22 && ~x23 && x16 && x11 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x66 && x67 && x24 && x26 && ~x20 && ~x21 && ~x22 && ~x23 && x16 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x66 && x67 && x24 && x26 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && x13 && x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x66 && x67 && x24 && x26 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && x13 && ~x11 && x12 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x66 && x67 && x24 && x26 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && x13 && ~x11 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x66 && x67 && x24 && x26 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && ~x13 && x11 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x66 && x67 && x24 && x26 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && ~x13 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x66 && x67 && x24 && x26 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x66 && x67 && x24 && ~x26 && x16 && x11 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x66 && x67 && x24 && ~x26 && x16 && x11 && ~x12 )
						begin
							y6 = 1'b1;	
							nx_state = s172;
						end
					else if( ~x66 && x67 && x24 && ~x26 && x16 && ~x11 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x66 && x67 && x24 && ~x26 && ~x16 && x17 && x11 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x66 && x67 && x24 && ~x26 && ~x16 && x17 && x11 && ~x13 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s46;
						end
					else if( ~x66 && x67 && x24 && ~x26 && ~x16 && x17 && ~x11 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x66 && x67 && x24 && ~x26 && ~x16 && ~x17 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && x67 && ~x24 && x25 && x26 && x4 && x15 && x10 && x11 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x66 && x67 && ~x24 && x25 && x26 && x4 && x15 && x10 && ~x11 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s65;
						end
					else if( ~x66 && x67 && ~x24 && x25 && x26 && x4 && x15 && x10 && ~x11 && ~x12 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s161;
						end
					else if( ~x66 && x67 && ~x24 && x25 && x26 && x4 && x15 && ~x10 && x12 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s186;
						end
					else if( ~x66 && x67 && ~x24 && x25 && x26 && x4 && x15 && ~x10 && ~x12 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x66 && x67 && ~x24 && x25 && x26 && x4 && ~x15 && x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x66 && x67 && ~x24 && x25 && x26 && x4 && ~x15 && ~x16 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && x67 && ~x24 && x25 && x26 && ~x4 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x66 && x67 && ~x24 && x25 && ~x26 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x66 && x67 && ~x24 && x25 && ~x26 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x66 && x67 && ~x24 && x25 && ~x26 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && x25 && ~x26 && ~x19 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && x10 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && x10 && ~x12 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && ~x10 && x11 && x12 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s171;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && ~x10 && x11 && ~x12 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && ~x10 && ~x11 && x12 && x13 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s239;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && ~x10 && ~x11 && x12 && ~x13 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && ~x10 && ~x11 && x12 && ~x13 && x18 && ~x14 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && ~x10 && ~x11 && x12 && ~x13 && ~x18 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && ~x10 && ~x11 && ~x12 && x14 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s239;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && ~x10 && ~x11 && ~x12 && ~x14 && x18 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && ~x10 && ~x11 && ~x12 && ~x14 && x18 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && x17 && ~x10 && ~x11 && ~x12 && ~x14 && ~x18 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && x12 && x10 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && x12 && x10 && ~x2 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && x12 && x10 && ~x2 && ~x4 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s382;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && x12 && ~x10 && x11 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && x12 && ~x10 && ~x11 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && x12 && ~x10 && ~x11 && ~x2 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && x12 && ~x10 && ~x11 && ~x2 && ~x4 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s382;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && ~x12 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && ~x12 && ~x2 && x11 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && ~x12 && ~x2 && x11 && ~x4 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s382;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && ~x12 && ~x2 && ~x11 && x10 && x4 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && ~x12 && ~x2 && ~x11 && x10 && ~x4 )
						begin
							y14 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && ~x12 && ~x2 && ~x11 && ~x10 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && x26 && ~x17 && ~x12 && ~x2 && ~x11 && ~x10 && ~x4 )
						begin
							y8 = 1'b1;	y17 = 1'b1;	y23 = 1'b1;	
							nx_state = s164;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && x10 && x12 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && x10 && ~x12 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && ~x10 && x11 && x12 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && ~x10 && x11 && ~x12 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s171;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && ~x10 && ~x11 && x12 && x13 )
						begin
							y8 = 1'b1;	
							nx_state = s181;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && ~x10 && ~x11 && x12 && ~x13 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && ~x10 && ~x11 && x12 && ~x13 && x17 && ~x14 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && ~x10 && ~x11 && x12 && ~x13 && ~x17 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && ~x10 && ~x11 && ~x12 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s181;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && ~x10 && ~x11 && ~x12 && ~x14 && x17 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && ~x10 && ~x11 && ~x12 && ~x14 && x17 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && x15 && ~x10 && ~x11 && ~x12 && ~x14 && ~x17 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && x10 && x8 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && x10 && x8 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && x10 && x8 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && x10 && x8 && ~x17 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && x10 && ~x8 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && x10 && ~x8 && ~x3 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && x10 && ~x8 && ~x3 && ~x5 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && ~x10 && x7 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && ~x10 && x7 && ~x3 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && ~x10 && x7 && ~x3 && ~x5 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && ~x10 && ~x7 && x11 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && ~x10 && ~x7 && x11 && ~x3 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && ~x10 && ~x7 && x11 && ~x3 && ~x5 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && ~x10 && ~x7 && ~x11 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && ~x10 && ~x7 && ~x11 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && ~x10 && ~x7 && ~x11 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && x12 && ~x10 && ~x7 && ~x11 && ~x17 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && x10 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && x10 && ~x3 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s172;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && x10 && ~x3 && ~x5 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && x11 && x9 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && x11 && x9 && ~x3 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && x11 && x9 && ~x3 && ~x5 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && ~x17 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && ~x11 && x8 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && ~x11 && x8 && ~x3 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && ~x11 && x8 && ~x3 && ~x5 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && x16 && ~x26 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && ~x17 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && x10 && x8 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && x10 && x8 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && x10 && x8 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && x10 && x8 && ~x18 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && x10 && ~x8 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && x10 && ~x8 && ~x2 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && x10 && ~x8 && ~x2 && ~x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && ~x10 && x7 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && ~x10 && x7 && ~x2 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && ~x10 && x7 && ~x2 && ~x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && ~x10 && ~x7 && x11 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && ~x10 && ~x7 && x11 && ~x2 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && ~x10 && ~x7 && x11 && ~x2 && ~x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && ~x10 && ~x7 && ~x11 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && ~x10 && ~x7 && ~x11 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && ~x10 && ~x7 && ~x11 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && x12 && ~x10 && ~x7 && ~x11 && ~x18 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && x10 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && x10 && ~x2 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s297;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && x10 && ~x2 && ~x4 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && x11 && x9 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && x11 && x9 && ~x2 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && x11 && x9 && ~x2 && ~x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && x11 && ~x9 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && x11 && ~x9 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && x11 && ~x9 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && x11 && ~x9 && ~x18 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && ~x11 && x8 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && ~x11 && x8 && ~x2 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && ~x11 && x8 && ~x2 && ~x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && ~x11 && ~x8 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && ~x11 && ~x8 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && ~x11 && ~x8 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && x17 && ~x12 && ~x10 && ~x11 && ~x8 && ~x18 )
						nx_state = s1;
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && ~x17 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && ~x17 && ~x2 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && x26 && ~x17 && ~x2 && ~x4 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s382;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && x12 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && x12 && ~x3 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && x12 && ~x3 && ~x5 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && x15 && x11 && x10 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && x15 && x11 && x10 && ~x3 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && x15 && x11 && x10 && ~x3 && ~x5 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && x15 && x11 && ~x10 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && x15 && ~x11 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && x15 && ~x11 && ~x3 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && x15 && ~x11 && ~x3 && ~x5 && x10 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && x15 && ~x11 && ~x3 && ~x5 && ~x10 )
						begin
							y14 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && ~x15 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s242;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && ~x15 && ~x3 && x5 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && x67 && ~x24 && ~x25 && ~x16 && ~x26 && ~x12 && ~x15 && ~x3 && ~x5 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && ~x67 && x21 && x68 && x12 && x7 && x19 && x17 )
						begin
							y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s383;
						end
					else if( ~x66 && ~x67 && x21 && x68 && x12 && x7 && x19 && ~x17 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s385;
						end
					else if( ~x66 && ~x67 && x21 && x68 && x12 && x7 && ~x19 && x20 )
						begin
							y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s383;
						end
					else if( ~x66 && ~x67 && x21 && x68 && x12 && x7 && ~x19 && ~x20 )
						begin
							y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s384;
						end
					else if( ~x66 && ~x67 && x21 && x68 && x12 && ~x7 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s385;
						end
					else if( ~x66 && ~x67 && x21 && x68 && ~x12 && x19 && x7 && x17 )
						begin
							y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s383;
						end
					else if( ~x66 && ~x67 && x21 && x68 && ~x12 && x19 && x7 && ~x17 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x66 && ~x67 && x21 && x68 && ~x12 && x19 && ~x7 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s385;
						end
					else if( ~x66 && ~x67 && x21 && x68 && ~x12 && ~x19 && x20 && x17 && x14 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s385;
						end
					else if( ~x66 && ~x67 && x21 && x68 && ~x12 && ~x19 && x20 && x17 && ~x14 && x16 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s385;
						end
					else if( ~x66 && ~x67 && x21 && x68 && ~x12 && ~x19 && x20 && x17 && ~x14 && ~x16 )
						nx_state = s1;
					else if( ~x66 && ~x67 && x21 && x68 && ~x12 && ~x19 && x20 && ~x17 && x16 && x15 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s385;
						end
					else if( ~x66 && ~x67 && x21 && x68 && ~x12 && ~x19 && x20 && ~x17 && x16 && ~x15 )
						nx_state = s1;
					else if( ~x66 && ~x67 && x21 && x68 && ~x12 && ~x19 && x20 && ~x17 && ~x16 && x13 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s385;
						end
					else if( ~x66 && ~x67 && x21 && x68 && ~x12 && ~x19 && x20 && ~x17 && ~x16 && ~x13 )
						nx_state = s1;
					else if( ~x66 && ~x67 && x21 && x68 && ~x12 && ~x19 && ~x20 && x7 )
						begin
							y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s376;
						end
					else if( ~x66 && ~x67 && x21 && x68 && ~x12 && ~x19 && ~x20 && ~x7 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s385;
						end
					else if( ~x66 && ~x67 && x21 && ~x68 && x19 && x7 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y17 = 1'b1;	
							nx_state = s177;
						end
					else if( ~x66 && ~x67 && x21 && ~x68 && x19 && ~x7 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && x15 && x14 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && x15 && ~x14 && x16 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && x15 && ~x14 && ~x16 && x9 && x3 )
						nx_state = s40;
					else if( ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && x15 && ~x14 && ~x16 && x9 && ~x3 && x4 )
						nx_state = s40;
					else if( ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && x15 && ~x14 && ~x16 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && x15 && ~x14 && ~x16 && ~x9 )
						nx_state = s1;
					else if( ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && ~x15 && x14 && x18 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && ~x15 && x14 && ~x18 && x9 && x3 )
						nx_state = s40;
					else if( ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && ~x15 && x14 && ~x18 && x9 && ~x3 && x4 )
						nx_state = s40;
					else if( ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && ~x15 && x14 && ~x18 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && ~x15 && x14 && ~x18 && ~x9 )
						nx_state = s1;
					else if( ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && ~x15 && ~x14 && x17 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x9 && x3 )
						nx_state = s40;
					else if( ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x9 && ~x3 && x4 )
						nx_state = s40;
					else if( ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( ~x66 && ~x67 && x21 && ~x68 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && ~x9 )
						nx_state = s1;
					else if( ~x66 && ~x67 && x21 && ~x68 && ~x19 && ~x20 && x7 )
						begin
							y21 = 1'b1;	
							nx_state = s151;
						end
					else if( ~x66 && ~x67 && x21 && ~x68 && ~x19 && ~x20 && ~x7 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x66 && ~x67 && ~x21 && x22 && x68 && x12 && x18 && x17 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x66 && ~x67 && ~x21 && x22 && x68 && x12 && x18 && ~x17 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s386;
						end
					else if( ~x66 && ~x67 && ~x21 && x22 && x68 && x12 && ~x18 && x19 && x17 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x66 && ~x67 && ~x21 && x22 && x68 && x12 && ~x18 && x19 && ~x17 && x3 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s387;
						end
					else if( ~x66 && ~x67 && ~x21 && x22 && x68 && x12 && ~x18 && x19 && ~x17 && ~x3 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x66 && ~x67 && ~x21 && x22 && x68 && x12 && ~x18 && ~x19 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x66 && ~x67 && ~x21 && x22 && x68 && ~x12 && x18 && x17 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x66 && ~x67 && ~x21 && x22 && x68 && ~x12 && x18 && ~x17 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s374;
						end
					else if( ~x66 && ~x67 && ~x21 && x22 && x68 && ~x12 && ~x18 && x19 )
						begin
							y4 = 1'b1;	y21 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x66 && ~x67 && ~x21 && x22 && x68 && ~x12 && ~x18 && ~x19 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x66 && ~x67 && ~x21 && x22 && ~x68 )
						nx_state = s1;
					else if( ~x66 && ~x67 && ~x21 && ~x22 && x68 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && x13 && x20 && x15 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && x13 && x20 && ~x15 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && x13 && ~x20 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && x14 && x20 && x15 )
						begin
							y22 = 1'b1;	y25 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && x14 && x20 && ~x15 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	y23 = 1'b1;	
							nx_state = s373;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && x14 && ~x20 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && x20 && x15 && x6 )
						begin
							y8 = 1'b1;	
							nx_state = s181;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && x20 && x15 && ~x6 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && x20 && x15 && ~x6 && x4 && ~x5 )
						nx_state = s1;
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && x20 && x15 && ~x6 && ~x4 )
						nx_state = s1;
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && x20 && ~x15 && x5 )
						begin
							y8 = 1'b1;	
							nx_state = s181;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && x20 && ~x15 && ~x5 && x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && x20 && ~x15 && ~x5 && x4 && ~x6 )
						nx_state = s1;
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && x20 && ~x15 && ~x5 && ~x4 )
						nx_state = s1;
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && ~x20 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s328;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && ~x20 && ~x3 && x7 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y17 = 1'b1;	
							nx_state = s177;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && ~x20 && ~x3 && ~x7 && x15 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s126;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && x19 && ~x13 && ~x14 && ~x20 && ~x3 && ~x7 && ~x15 )
						begin
							y2 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s371;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s328;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && x14 && x18 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && x14 && ~x18 && x15 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && x14 && ~x18 && ~x15 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && x14 && ~x18 && ~x15 && x4 && ~x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && x14 && ~x18 && ~x15 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && x14 && ~x18 && ~x15 && ~x4 )
						nx_state = s1;
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && ~x14 && x15 && x16 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && ~x14 && x15 && ~x16 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && ~x14 && x15 && ~x16 && x4 && ~x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && ~x14 && x15 && ~x16 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && ~x14 && x15 && ~x16 && ~x4 )
						nx_state = s1;
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && ~x14 && ~x15 && x17 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && ~x14 && ~x15 && ~x17 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && ~x14 && ~x15 && ~x17 && x4 && ~x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && ~x14 && ~x15 && ~x17 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && x20 && ~x14 && ~x15 && ~x17 && ~x4 )
						nx_state = s1;
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && ~x20 && x7 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y17 = 1'b1;	
							nx_state = s177;
						end
					else if( ~x66 && ~x67 && ~x21 && ~x22 && ~x68 && ~x19 && ~x3 && ~x20 && ~x7 )
						begin
							y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s377;
						end
					else nx_state = s110;
				s111 : if( x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x22 && ~x17 )
						nx_state = s1;
					else if( ~x22 && x18 && x13 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x22 && x18 && x13 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x22 && x18 && ~x13 && x12 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x22 && x18 && ~x13 && x12 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x22 && ~x18 )
						nx_state = s1;
					else nx_state = s111;
				s112 : if( x65 && x66 && x22 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	
							nx_state = s111;
						end
					else if( x65 && x66 && ~x22 && x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && x66 && ~x22 && ~x23 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x65 && ~x66 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x5 )
						nx_state = s1;
					else if( ~x65 && x66 && x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x65 && x66 && x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x65 && x66 && x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x66 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x21 && x22 && x23 )
						begin
							y14 = 1'b1;	
							nx_state = s286;
						end
					else if( ~x65 && x66 && ~x21 && x22 && ~x23 && x18 && x14 )
						nx_state = s40;
					else if( ~x65 && x66 && ~x21 && x22 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s40;
					else if( ~x65 && x66 && ~x21 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x21 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x21 && ~x22 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x21 && ~x22 && x23 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x21 && ~x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && ~x66 && x20 && x15 && x16 && x8 && x14 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x65 && ~x66 && x20 && x15 && x16 && x8 && ~x14 && x7 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s126;
						end
					else if( ~x65 && ~x66 && x20 && x15 && x16 && x8 && ~x14 && ~x7 && x12 )
						begin
							y4 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x65 && ~x66 && x20 && x15 && x16 && x8 && ~x14 && ~x7 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x20 && x15 && x16 && ~x8 && x14 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x66 && x20 && x15 && x16 && ~x8 && ~x14 && x7 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	y20 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x65 && ~x66 && x20 && x15 && x16 && ~x8 && ~x14 && ~x7 && x13 )
						begin
							y4 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x65 && ~x66 && x20 && x15 && x16 && ~x8 && ~x14 && ~x7 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x20 && x15 && ~x16 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s191;
						end
					else if( ~x65 && ~x66 && x20 && x15 && ~x16 && ~x7 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x65 && ~x66 && x20 && x15 && ~x16 && ~x7 && ~x5 && x8 && x1 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x65 && ~x66 && x20 && x15 && ~x16 && ~x7 && ~x5 && x8 && ~x1 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( ~x65 && ~x66 && x20 && x15 && ~x16 && ~x7 && ~x5 && ~x8 && x1 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x65 && ~x66 && x20 && x15 && ~x16 && ~x7 && ~x5 && ~x8 && ~x1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && x7 && x8 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && x7 && x8 && ~x5 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && x7 && ~x8 && x11 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && x7 && ~x8 && x11 && ~x5 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && x7 && ~x8 && ~x11 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && x7 && ~x8 && ~x11 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && x7 && ~x8 && ~x11 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && x7 && ~x8 && ~x11 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && x8 && x9 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && x8 && x9 && ~x5 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && x8 && ~x9 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && x8 && ~x9 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && x8 && ~x9 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && x8 && ~x9 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && ~x8 && x10 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && ~x8 && x10 && ~x5 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && ~x8 && ~x10 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && ~x8 && ~x10 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && ~x8 && ~x10 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x20 && ~x15 && x16 && ~x7 && ~x8 && ~x10 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x20 && ~x15 && ~x16 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s44;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && ~x16 && ~x5 && x1 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x65 && ~x66 && x20 && ~x15 && ~x16 && ~x5 && ~x1 )
						begin
							y12 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x65 && ~x66 && ~x20 )
						nx_state = s1;
					else nx_state = s112;
				s113 : if( x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x21 && ~x19 )
						nx_state = s1;
					else if( ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x21 && ~x20 )
						nx_state = s1;
					else nx_state = s113;
				s114 : if( x67 && x65 && x21 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x67 && x65 && x21 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x67 && x65 && x21 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x67 && x65 && x21 && ~x8 )
						nx_state = s1;
					else if( x67 && x65 && ~x21 && x23 && x22 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x67 && x65 && ~x21 && x23 && x22 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x67 && x65 && ~x21 && x23 && x22 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x67 && x65 && ~x21 && x23 && x22 && ~x8 )
						nx_state = s1;
					else if( x67 && x65 && ~x21 && x23 && ~x22 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x67 && x65 && ~x21 && x23 && ~x22 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x67 && x65 && ~x21 && x23 && ~x22 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x67 && x65 && ~x21 && x23 && ~x22 && ~x9 )
						nx_state = s1;
					else if( x67 && x65 && ~x21 && ~x23 && x8 && x22 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x67 && x65 && ~x21 && ~x23 && x8 && x22 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x67 && x65 && ~x21 && ~x23 && x8 && x22 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x67 && x65 && ~x21 && ~x23 && x8 && ~x22 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x67 && x65 && ~x21 && ~x23 && x8 && ~x22 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x67 && x65 && ~x21 && ~x23 && x8 && ~x22 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x67 && x65 && ~x21 && ~x23 && ~x8 )
						nx_state = s1;
					else if( x67 && ~x65 && x66 && x68 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x67 && ~x65 && x66 && x68 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x67 && ~x65 && x66 && x68 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x67 && ~x65 && x66 && x68 && x21 && ~x19 )
						nx_state = s1;
					else if( x67 && ~x65 && x66 && x68 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x67 && ~x65 && x66 && x68 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x67 && ~x65 && x66 && x68 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x67 && ~x65 && x66 && x68 && ~x21 && ~x20 )
						nx_state = s1;
					else if( x67 && ~x65 && x66 && ~x68 )
						nx_state = s1;
					else if( x67 && ~x65 && ~x66 && x24 && x26 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y21 = 1'b1;	
							nx_state = s183;
						end
					else if( x67 && ~x65 && ~x66 && x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( x67 && ~x65 && ~x66 && x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( x67 && ~x65 && ~x66 && x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x67 && ~x65 && ~x66 && x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( x67 && ~x65 && ~x66 && ~x24 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( x67 && ~x65 && ~x66 && ~x24 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( x67 && ~x65 && ~x66 && ~x24 && x25 && x19 && ~x14 && ~x13 && x26 )
						nx_state = s114;
					else if( x67 && ~x65 && ~x66 && ~x24 && x25 && x19 && ~x14 && ~x13 && ~x26 )
						nx_state = s1;
					else if( x67 && ~x65 && ~x66 && ~x24 && x25 && ~x19 )
						nx_state = s1;
					else if( x67 && ~x65 && ~x66 && ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( x67 && ~x65 && ~x66 && ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( x67 && ~x65 && ~x66 && ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x67 && ~x65 && ~x66 && ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( x67 && ~x65 && ~x66 && ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( x67 && ~x65 && ~x66 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( x67 && ~x65 && ~x66 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x67 && ~x65 && ~x66 && ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else if( ~x67 && x65 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x67 && x65 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x67 && x65 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x67 && x65 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x67 && x65 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( ~x67 && x65 && ~x21 && x23 && x22 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( ~x67 && x65 && ~x21 && x23 && x22 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( ~x67 && x65 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( ~x67 && x65 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x67 && x65 && ~x21 && x23 && x22 && ~x19 && ~x17 )
						nx_state = s1;
					else if( ~x67 && x65 && ~x21 && x23 && ~x22 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( ~x67 && x65 && ~x21 && x23 && ~x22 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( ~x67 && x65 && ~x21 && x23 && ~x22 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x67 && x65 && ~x21 && x23 && ~x22 && ~x20 )
						nx_state = s1;
					else if( ~x67 && x65 && ~x21 && ~x23 && x18 && x14 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( ~x67 && x65 && ~x21 && ~x23 && x18 && x14 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x67 && x65 && ~x21 && ~x23 && x18 && ~x14 && x13 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( ~x67 && x65 && ~x21 && ~x23 && x18 && ~x14 && x13 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x67 && x65 && ~x21 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x67 && x65 && ~x21 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x67 && ~x65 && x21 && x66 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x67 && ~x65 && x21 && x66 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x67 && ~x65 && x21 && x66 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x67 && ~x65 && x21 && x66 && ~x9 )
						nx_state = s1;
					else if( ~x67 && ~x65 && x21 && ~x66 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x67 && ~x65 && x21 && ~x66 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x67 && ~x65 && x21 && ~x66 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x67 && ~x65 && x21 && ~x66 && ~x3 )
						nx_state = s1;
					else if( ~x67 && ~x65 && ~x21 && x22 && x66 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x67 && ~x65 && ~x21 && x22 && ~x66 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x67 && ~x65 && ~x21 && ~x22 && x66 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x67 && ~x65 && ~x21 && ~x22 && x66 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x67 && ~x65 && ~x21 && ~x22 && x66 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x67 && ~x65 && ~x21 && ~x22 && x66 && ~x4 )
						nx_state = s1;
					else if( ~x67 && ~x65 && ~x21 && ~x22 && ~x66 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x67 && ~x65 && ~x21 && ~x22 && ~x66 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x67 && ~x65 && ~x21 && ~x22 && ~x66 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x67 && ~x65 && ~x21 && ~x22 && ~x66 && ~x8 )
						nx_state = s1;
					else nx_state = s114;
				s115 : if( x21 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s344;
						end
					else nx_state = s115;
				s116 : if( x21 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( ~x21 && x22 && x8 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x8 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x12 && x23 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x21 && ~x22 && x12 && ~x23 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x21 && ~x22 && ~x12 && x23 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && ~x12 && x23 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && ~x12 && x23 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x12 && x23 && ~x9 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x12 && ~x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && ~x12 && ~x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && ~x12 && ~x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x12 && ~x23 && ~x8 )
						nx_state = s1;
					else nx_state = s116;
				s117 : if( x21 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( ~x21 && x22 && x23 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x21 && x22 && x23 && ~x12 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x23 && ~x12 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x23 && ~x12 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x12 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x8 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x8 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && ~x18 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s243;
						end
					else nx_state = s117;
				s118 : if( x60 && x61 && x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s38;
						end
					else if( x60 && x61 && ~x18 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( x60 && ~x61 )
						begin
							y11 = 1'b1;	
							nx_state = s356;
						end
					else if( ~x60 && x61 )
						begin
							y11 = 1'b1;	
							nx_state = s356;
						end
					else if( ~x60 && ~x61 && x62 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x60 && ~x61 && ~x62 )
						begin
							y7 = 1'b1;	
							nx_state = s338;
						end
					else nx_state = s118;
				s119 : if( x21 && x15 && x16 && x9 && x7 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && x15 && x16 && x9 && ~x7 && x8 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s157;
						end
					else if( x21 && x15 && x16 && x9 && ~x7 && ~x8 && x13 )
						begin
							y4 = 1'b1;	
							nx_state = s191;
						end
					else if( x21 && x15 && x16 && x9 && ~x7 && ~x8 && ~x13 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x21 && x15 && x16 && x9 && ~x7 && ~x8 && ~x13 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x21 && x15 && x16 && x9 && ~x7 && ~x8 && ~x13 && ~x18 && x19 && ~x14 )
						nx_state = s1;
					else if( x21 && x15 && x16 && x9 && ~x7 && ~x8 && ~x13 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x21 && x15 && x16 && ~x9 && x7 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x21 && x15 && x16 && ~x9 && ~x7 && x8 )
						begin
							y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s158;
						end
					else if( x21 && x15 && x16 && ~x9 && ~x7 && ~x8 && x14 )
						begin
							y4 = 1'b1;	
							nx_state = s191;
						end
					else if( x21 && x15 && x16 && ~x9 && ~x7 && ~x8 && ~x14 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( x21 && x15 && ~x16 && x7 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s147;
						end
					else if( x21 && x15 && ~x16 && ~x7 && x8 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s147;
						end
					else if( x21 && x15 && ~x16 && ~x7 && ~x8 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s22;
						end
					else if( x21 && x15 && ~x16 && ~x7 && ~x8 && ~x2 && x5 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x21 && x15 && ~x16 && ~x7 && ~x8 && ~x2 && ~x5 && x9 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x21 && x15 && ~x16 && ~x7 && ~x8 && ~x2 && ~x5 && ~x9 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( x21 && ~x15 && x2 )
						begin
							y1 = 1'b1;	
							nx_state = s22;
						end
					else if( x21 && ~x15 && ~x2 && x16 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && ~x15 && ~x2 && x16 && x9 && ~x10 && x8 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && ~x15 && ~x2 && x16 && x9 && ~x10 && ~x8 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x21 && ~x15 && ~x2 && x16 && x9 && ~x10 && ~x8 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x21 && ~x15 && ~x2 && x16 && x9 && ~x10 && ~x8 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x21 && ~x15 && ~x2 && x16 && x9 && ~x10 && ~x8 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x15 && ~x2 && x16 && x9 && ~x10 && ~x8 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x21 && ~x15 && ~x2 && x16 && ~x9 && x8 && x12 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && ~x15 && ~x2 && x16 && ~x9 && x8 && ~x12 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x21 && ~x15 && ~x2 && x16 && ~x9 && x8 && ~x12 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x21 && ~x15 && ~x2 && x16 && ~x9 && x8 && ~x12 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x21 && ~x15 && ~x2 && x16 && ~x9 && x8 && ~x12 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x15 && ~x2 && x16 && ~x9 && x8 && ~x12 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x21 && ~x15 && ~x2 && x16 && ~x9 && ~x8 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && ~x15 && ~x2 && x16 && ~x9 && ~x8 && ~x11 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x21 && ~x15 && ~x2 && x16 && ~x9 && ~x8 && ~x11 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x21 && ~x15 && ~x2 && x16 && ~x9 && ~x8 && ~x11 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x21 && ~x15 && ~x2 && x16 && ~x9 && ~x8 && ~x11 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x15 && ~x2 && x16 && ~x9 && ~x8 && ~x11 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x21 && ~x15 && ~x2 && ~x16 && x5 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x21 && ~x15 && ~x2 && ~x16 && ~x5 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x21 && x22 && x18 && x14 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( ~x21 && x22 && x18 && ~x14 && x13 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( ~x21 && x22 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x18 )
						nx_state = s1;
					else if( ~x21 && ~x22 )
						nx_state = s1;
					else nx_state = s119;
				s120 : if( x21 )
						begin
							y20 = 1'b1;	
							nx_state = s363;
						end
					else if( ~x21 && x23 && x22 && x5 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && x23 && x22 && ~x5 && x18 && x15 && x9 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x21 && x23 && x22 && ~x5 && x18 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x21 && x23 && x22 && ~x5 && x18 && ~x15 && x16 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x21 && x23 && x22 && ~x5 && x18 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x21 && x23 && x22 && ~x5 && ~x18 )
						begin
							y1 = 1'b1;	y5 = 1'b1;	y11 = 1'b1;	
							nx_state = s97;
						end
					else if( ~x21 && x23 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && ~x23 && x22 )
						nx_state = s1;
					else if( ~x21 && ~x23 && ~x22 && x15 && x9 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x21 && ~x23 && ~x22 && x15 && ~x9 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x15 && x16 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s205;
						end
					else nx_state = s120;
				s121 : if( x67 && x22 && x3 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x67 && x22 && x3 && x15 && ~x8 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s154;
						end
					else if( x67 && x22 && x3 && ~x15 && x16 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s255;
						end
					else if( x67 && x22 && x3 && ~x15 && ~x16 )
						begin
							y3 = 1'b1;	y11 = 1'b1;	
							nx_state = s6;
						end
					else if( x67 && x22 && ~x3 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s255;
						end
					else if( x67 && ~x22 && x23 && x18 && x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x67 && ~x22 && x23 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x67 && ~x22 && x23 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x67 && ~x22 && x23 && ~x18 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && x16 && x15 && x14 && x8 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( x67 && ~x22 && ~x23 && x16 && x15 && x14 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x67 && ~x22 && ~x23 && x16 && x15 && ~x14 && x7 && x8 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( x67 && ~x22 && ~x23 && x16 && x15 && ~x14 && x7 && ~x8 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s126;
						end
					else if( x67 && ~x22 && ~x23 && x16 && x15 && ~x14 && ~x7 && x8 && x12 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s125;
						end
					else if( x67 && ~x22 && ~x23 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && x18 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x67 && ~x22 && ~x23 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && x18 && ~x13 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && x16 && x15 && ~x14 && ~x7 && x8 && ~x12 && ~x18 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && x16 && x15 && ~x14 && ~x7 && ~x8 && x13 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s125;
						end
					else if( x67 && ~x22 && ~x23 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && x18 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x67 && ~x22 && ~x23 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && x18 && ~x12 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && x16 && x15 && ~x14 && ~x7 && ~x8 && ~x13 && ~x18 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && x8 && x9 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && x8 && x9 && ~x2 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && x8 && x9 && ~x2 && ~x3 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s111;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && x8 && ~x9 && x7 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && x8 && ~x9 && x7 && ~x2 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && x8 && ~x9 && x7 && ~x2 && ~x3 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s111;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && x8 && ~x9 && ~x7 && x18 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && x8 && ~x9 && ~x7 && x18 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && x8 && ~x9 && ~x7 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && x8 && ~x9 && ~x7 && ~x18 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && x7 && x11 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && x7 && x11 && ~x2 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && x7 && x11 && ~x2 && ~x3 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s111;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && x7 && ~x11 && x18 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && x7 && ~x11 && x18 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && x7 && ~x11 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && x7 && ~x11 && ~x18 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && ~x7 && x10 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && ~x7 && x10 && ~x2 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && ~x7 && x10 && ~x2 && ~x3 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s111;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && x18 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && x18 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && x16 && ~x15 && ~x8 && ~x7 && ~x10 && ~x18 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x23 && ~x16 && x15 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x67 && ~x22 && ~x23 && ~x16 && x15 && ~x7 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( x67 && ~x22 && ~x23 && ~x16 && x15 && ~x7 && ~x2 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x67 && ~x22 && ~x23 && ~x16 && x15 && ~x7 && ~x2 && ~x3 && x8 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y28 = 1'b1;	
							nx_state = s129;
						end
					else if( x67 && ~x22 && ~x23 && ~x16 && x15 && ~x7 && ~x2 && ~x3 && ~x8 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	
							nx_state = s111;
						end
					else if( x67 && ~x22 && ~x23 && ~x16 && ~x15 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else if( x67 && ~x22 && ~x23 && ~x16 && ~x15 && ~x2 && x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x67 && ~x22 && ~x23 && ~x16 && ~x15 && ~x2 && ~x3 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s127;
						end
					else if( ~x67 && x21 && x20 && x15 && x10 && x11 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x67 && x21 && x20 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s193;
						end
					else if( ~x67 && x21 && x20 && x15 && x10 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s194;
						end
					else if( ~x67 && x21 && x20 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s300;
						end
					else if( ~x67 && x21 && x20 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x67 && x21 && x20 && ~x15 && x16 && x10 && x12 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s259;
						end
					else if( ~x67 && x21 && x20 && ~x15 && x16 && x10 && ~x12 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x67 && x21 && x20 && ~x15 && x16 && ~x10 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s259;
						end
					else if( ~x67 && x21 && x20 && ~x15 && ~x16 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x67 && x21 && ~x20 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s57;
						end
					else if( ~x67 && ~x21 && x4 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s306;
						end
					else if( ~x67 && ~x21 && ~x4 && x18 && x15 && x10 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x67 && ~x21 && ~x4 && x18 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s301;
						end
					else if( ~x67 && ~x21 && ~x4 && x18 && x15 && x10 && ~x11 && ~x12 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s195;
						end
					else if( ~x67 && ~x21 && ~x4 && x18 && x15 && ~x10 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x67 && ~x21 && ~x4 && x18 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x67 && ~x21 && ~x4 && x18 && ~x15 && x16 && x10 && x12 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s259;
						end
					else if( ~x67 && ~x21 && ~x4 && x18 && ~x15 && x16 && x10 && ~x12 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x67 && ~x21 && ~x4 && x18 && ~x15 && x16 && ~x10 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s259;
						end
					else if( ~x67 && ~x21 && ~x4 && x18 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s303;
						end
					else if( ~x67 && ~x21 && ~x4 && ~x18 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s57;
						end
					else nx_state = s121;
				s122 : if( x65 && x22 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	
							nx_state = s111;
						end
					else if( x65 && ~x22 && x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x65 && ~x22 && ~x23 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x68 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x68 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x68 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && x68 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x68 && x23 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x68 && ~x23 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else nx_state = s122;
				s123 : if( x21 && x9 && x3 )
						nx_state = s40;
					else if( x21 && x9 && ~x3 && x4 )
						nx_state = s40;
					else if( x21 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( x21 && ~x9 )
						nx_state = s1;
					else if( ~x21 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x5 && ~x4 && x22 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x5 && ~x4 && x22 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x5 && ~x4 && ~x22 )
						nx_state = s1;
					else if( ~x21 && ~x5 && x22 )
						nx_state = s1;
					else if( ~x21 && ~x5 && ~x22 && x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && ~x5 && ~x22 && x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x5 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s123;
				s124 : if( x65 && x22 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s255;
						end
					else if( x65 && ~x22 && ~x23 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s389;
						end
					else if( ~x65 && x21 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x21 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x21 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && x21 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && ~x21 && x22 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && ~x21 && x22 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x7 )
						nx_state = s1;
					else if( ~x65 && ~x21 && ~x22 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s124;
				s125 : if( x67 && x22 )
						begin
							y2 = 1'b1;	y16 = 1'b1;	y24 = 1'b1;	
							nx_state = s124;
						end
					else if( x67 && ~x22 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x67 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s302;
						end
					else nx_state = s125;
				s126 : if( x65 && x67 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && x67 && x22 && ~x17 )
						nx_state = s1;
					else if( x65 && x67 && ~x22 && x18 && x13 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && x67 && ~x22 && x18 && x13 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x67 && ~x22 && x18 && ~x13 && x12 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && x67 && ~x22 && x18 && ~x13 && x12 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x67 && ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && x67 && ~x22 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x67 && x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x67 && x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x67 && x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x67 && x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && ~x67 && x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && ~x67 && x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x67 && ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x67 && ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x21 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && x21 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s143;
						end
					else if( ~x65 && x66 && ~x21 && x23 && x22 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x65 && x66 && ~x21 && x23 && ~x22 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x65 && x66 && ~x21 && x23 && ~x22 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x65 && x66 && ~x21 && x23 && ~x22 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x21 && x23 && ~x22 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x21 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && ~x66 && x67 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x66 && x67 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x66 && x67 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && x20 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x66 && x67 && ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x66 && x67 && ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x65 && ~x66 && x67 && ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x65 && ~x66 && x67 && ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x67 && ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && x21 && x19 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x67 && x21 && ~x19 && x20 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s176;
						end
					else if( ~x65 && ~x66 && ~x67 && x21 && ~x19 && ~x20 )
						begin
							y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s377;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && x13 && x20 && x15 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && x13 && x20 && ~x15 )
						begin
							y22 = 1'b1;	y25 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && x13 && ~x20 )
						begin
							y2 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s371;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && x20 && x14 && x15 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	y23 = 1'b1;	
							nx_state = s373;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && x20 && x14 && ~x15 )
						begin
							y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s377;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && x20 && ~x14 && x15 && x6 )
						begin
							y12 = 1'b1;	
							nx_state = s293;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && x20 && ~x14 && x15 && ~x6 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && x20 && ~x14 && x15 && ~x6 && x5 && ~x4 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && x20 && ~x14 && x15 && ~x6 && ~x5 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && x20 && ~x14 && ~x15 && x4 )
						begin
							y12 = 1'b1;	
							nx_state = s293;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && x20 && ~x14 && ~x15 && ~x4 && x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && x20 && ~x14 && ~x15 && ~x4 && x5 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && x20 && ~x14 && ~x15 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && ~x20 && x14 )
						begin
							y2 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s371;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && ~x20 && ~x14 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s329;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && ~x20 && ~x14 && ~x7 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && ~x20 && ~x14 && ~x7 && ~x8 && x15 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	
							nx_state = s378;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && x19 && ~x13 && ~x20 && ~x14 && ~x7 && ~x8 && ~x15 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && ~x19 && x7 )
						begin
							y4 = 1'b1;	
							nx_state = s329;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && ~x19 && ~x7 && x20 && x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && ~x19 && ~x7 && x20 && x15 && ~x14 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && ~x19 && ~x7 && x20 && ~x15 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && ~x19 && ~x7 && ~x20 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && x22 && ~x19 && ~x7 && ~x20 && ~x8 )
						begin
							y21 = 1'b1;	y24 = 1'b1;	
							nx_state = s225;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && ~x22 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x66 && ~x67 && ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x67 && ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s126;
				s127 : if( x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x22 && ~x17 )
						nx_state = s1;
					else if( ~x22 && x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x22 && ~x23 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else nx_state = s127;
				s128 : if( x65 && x67 && x22 && x15 && x8 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x67 && x22 && x15 && ~x8 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x65 && x67 && x22 && ~x15 && x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s50;
						end
					else if( x65 && x67 && x22 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s122;
						end
					else if( x65 && x67 && ~x22 && x15 && x8 && x23 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x67 && ~x22 && x15 && x8 && ~x23 )
						begin
							y11 = 1'b1;	
							nx_state = s8;
						end
					else if( x65 && x67 && ~x22 && x15 && ~x8 && x23 && x6 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s111;
						end
					else if( x65 && x67 && ~x22 && x15 && ~x8 && x23 && ~x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x67 && ~x22 && x15 && ~x8 && ~x23 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s111;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && x8 && x7 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && x8 && ~x7 && x9 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && x8 && ~x7 && ~x9 && x18 && x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && x8 && ~x7 && ~x9 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && x8 && ~x7 && ~x9 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && x8 && ~x7 && ~x9 && ~x18 )
						nx_state = s1;
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && ~x8 && x7 && x11 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && ~x8 && x7 && ~x11 && x18 && x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && ~x8 && x7 && ~x11 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && ~x8 && x7 && ~x11 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && ~x8 && x7 && ~x11 && ~x18 )
						nx_state = s1;
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && ~x8 && ~x7 && x10 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && ~x8 && ~x7 && ~x10 && x18 && x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && ~x8 && ~x7 && ~x10 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && ~x8 && ~x7 && ~x10 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && x67 && ~x22 && ~x15 && x16 && x23 && ~x8 && ~x7 && ~x10 && ~x18 )
						nx_state = s1;
					else if( x65 && x67 && ~x22 && ~x15 && x16 && ~x23 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s154;
						end
					else if( x65 && x67 && ~x22 && ~x15 && ~x16 && x23 && x6 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( x65 && x67 && ~x22 && ~x15 && ~x16 && x23 && ~x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x67 && ~x22 && ~x15 && ~x16 && ~x23 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( x65 && ~x67 && x61 && x60 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s67;
						end
					else if( x65 && ~x67 && x61 && ~x60 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( x65 && ~x67 && ~x61 && x60 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( x65 && ~x67 && ~x61 && ~x60 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && x22 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s79;
						end
					else if( ~x65 && ~x22 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else nx_state = s128;
				s129 : if( x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x22 && ~x17 )
						nx_state = s1;
					else if( ~x22 && x23 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( ~x22 && x23 && x15 && ~x8 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x22 && x23 && ~x15 && x16 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s111;
						end
					else if( ~x22 && x23 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s122;
						end
					else if( ~x22 && ~x23 && x18 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x22 && ~x23 && x18 && ~x13 && x12 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x22 && ~x23 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x22 && ~x23 && ~x18 )
						nx_state = s1;
					else nx_state = s129;
				s130 : if( x65 && x22 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s121;
						end
					else if( x65 && ~x22 && x23 && x15 && x16 && x14 && x8 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( x65 && ~x22 && x23 && x15 && x16 && x14 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x65 && ~x22 && x23 && x15 && x16 && ~x14 && x7 && x8 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( x65 && ~x22 && x23 && x15 && x16 && ~x14 && x7 && ~x8 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s126;
						end
					else if( x65 && ~x22 && x23 && x15 && x16 && ~x14 && ~x7 && x8 && x12 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s302;
						end
					else if( x65 && ~x22 && x23 && x15 && x16 && ~x14 && ~x7 && x8 && ~x12 && x18 && x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && ~x22 && x23 && x15 && x16 && ~x14 && ~x7 && x8 && ~x12 && x18 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 && x15 && x16 && ~x14 && ~x7 && x8 && ~x12 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 && x15 && x16 && ~x14 && ~x7 && ~x8 && x13 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s302;
						end
					else if( x65 && ~x22 && x23 && x15 && x16 && ~x14 && ~x7 && ~x8 && ~x13 && x18 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && ~x22 && x23 && x15 && x16 && ~x14 && ~x7 && ~x8 && ~x13 && x18 && ~x12 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 && x15 && x16 && ~x14 && ~x7 && ~x8 && ~x13 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 && x15 && ~x16 && x7 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x65 && ~x22 && x23 && x15 && ~x16 && ~x7 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s44;
						end
					else if( x65 && ~x22 && x23 && x15 && ~x16 && ~x7 && ~x2 && x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y28 = 1'b1;	
							nx_state = s129;
						end
					else if( x65 && ~x22 && x23 && x15 && ~x16 && ~x7 && ~x2 && ~x3 && x8 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s121;
						end
					else if( x65 && ~x22 && x23 && x15 && ~x16 && ~x7 && ~x2 && ~x3 && ~x8 )
						begin
							y9 = 1'b1;	y12 = 1'b1;	
							nx_state = s111;
						end
					else if( x65 && ~x22 && x23 && ~x15 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s44;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && x7 && x11 && x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y28 = 1'b1;	
							nx_state = s129;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && x7 && x11 && ~x3 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s154;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && x7 && ~x11 && x8 && x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y28 = 1'b1;	
							nx_state = s129;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && x7 && ~x11 && x8 && ~x3 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s154;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && x7 && ~x11 && ~x8 && x18 && x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && x7 && ~x11 && ~x8 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && x7 && ~x11 && ~x8 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && x7 && ~x11 && ~x8 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && x8 && x9 && x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y28 = 1'b1;	
							nx_state = s129;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && x8 && x9 && ~x3 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s154;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && x8 && ~x9 && x18 && x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && x8 && ~x9 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && x8 && ~x9 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && x8 && ~x9 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && x10 && x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y28 = 1'b1;	
							nx_state = s129;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && x10 && ~x3 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s154;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && ~x10 && x18 && x13 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && ~x10 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && ~x10 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && ~x10 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && ~x16 && x3 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y28 = 1'b1;	
							nx_state = s129;
						end
					else if( x65 && ~x22 && x23 && ~x15 && ~x2 && ~x16 && ~x3 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y12 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s127;
						end
					else if( x65 && ~x22 && ~x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x65 && x67 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x65 && x67 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x65 && x67 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s151;
						end
					else if( ~x65 && x67 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y28 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x65 && ~x67 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else nx_state = s130;
				s131 : if( x68 && x6 && x15 && x10 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s301;
						end
					else if( x68 && x6 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s192;
						end
					else if( x68 && x6 && x15 && x10 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s60;
						end
					else if( x68 && x6 && x15 && ~x10 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s196;
						end
					else if( x68 && x6 && x15 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	
							nx_state = s61;
						end
					else if( x68 && x6 && ~x15 && x16 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s60;
						end
					else if( x68 && x6 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s303;
						end
					else if( x68 && ~x6 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s60;
						end
					else if( ~x68 && x60 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s68;
						end
					else if( ~x68 && ~x60 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else nx_state = s131;
				s132 : if( x21 && x15 && x20 && x10 && x11 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s192;
						end
					else if( x21 && x15 && x20 && x10 && ~x11 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s193;
						end
					else if( x21 && x15 && x20 && ~x10 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s300;
						end
					else if( x21 && x15 && x20 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s192;
						end
					else if( x21 && x15 && ~x20 && x5 && x10 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s301;
						end
					else if( x21 && x15 && ~x20 && x5 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s192;
						end
					else if( x21 && x15 && ~x20 && x5 && x10 && ~x11 && ~x12 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( x21 && x15 && ~x20 && x5 && ~x10 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s196;
						end
					else if( x21 && x15 && ~x20 && x5 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	
							nx_state = s61;
						end
					else if( x21 && x15 && ~x20 && ~x5 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( x21 && ~x15 && x16 && x10 && x12 && x20 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y11 = 1'b1;	
							nx_state = s192;
						end
					else if( x21 && ~x15 && x16 && x10 && x12 && ~x20 && x8 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( x21 && ~x15 && x16 && x10 && x12 && ~x20 && ~x8 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x15 && x16 && x10 && x12 && ~x20 && ~x8 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x15 && x16 && x10 && x12 && ~x20 && ~x8 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x15 && x16 && x10 && x12 && ~x20 && ~x8 && ~x19 )
						nx_state = s1;
					else if( x21 && ~x15 && x16 && x10 && ~x12 && x20 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( x21 && ~x15 && x16 && x10 && ~x12 && ~x20 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( x21 && ~x15 && x16 && ~x10 && x20 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y11 = 1'b1;	
							nx_state = s192;
						end
					else if( x21 && ~x15 && x16 && ~x10 && ~x20 && x12 && x7 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( x21 && ~x15 && x16 && ~x10 && ~x20 && x12 && ~x7 && x11 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( x21 && ~x15 && x16 && ~x10 && ~x20 && x12 && ~x7 && ~x11 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x15 && x16 && ~x10 && ~x20 && x12 && ~x7 && ~x11 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x15 && x16 && ~x10 && ~x20 && x12 && ~x7 && ~x11 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x15 && x16 && ~x10 && ~x20 && x12 && ~x7 && ~x11 && ~x19 )
						nx_state = s1;
					else if( x21 && ~x15 && x16 && ~x10 && ~x20 && ~x12 && x11 && x9 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( x21 && ~x15 && x16 && ~x10 && ~x20 && ~x12 && x11 && ~x9 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x15 && x16 && ~x10 && ~x20 && ~x12 && x11 && ~x9 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x15 && x16 && ~x10 && ~x20 && ~x12 && x11 && ~x9 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x15 && x16 && ~x10 && ~x20 && ~x12 && x11 && ~x9 && ~x19 )
						nx_state = s1;
					else if( x21 && ~x15 && x16 && ~x10 && ~x20 && ~x12 && ~x11 && x8 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x15 && x16 && ~x10 && ~x20 && ~x12 && ~x11 && x8 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x15 && x16 && ~x10 && ~x20 && ~x12 && ~x11 && x8 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x15 && x16 && ~x10 && ~x20 && ~x12 && ~x11 && x8 && ~x19 )
						nx_state = s1;
					else if( x21 && ~x15 && x16 && ~x10 && ~x20 && ~x12 && ~x11 && ~x8 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( x21 && ~x15 && ~x16 && x20 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x21 && ~x15 && ~x16 && ~x20 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x21 && ~x15 && ~x16 && ~x20 && ~x5 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x21 && x3 && x15 && x10 && x11 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x21 && x3 && x15 && x10 && ~x11 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s193;
						end
					else if( ~x21 && x3 && x15 && x10 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y13 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x21 && x3 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s300;
						end
					else if( ~x21 && x3 && x15 && ~x10 && ~x12 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x21 && x3 && ~x15 && x16 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s121;
						end
					else if( ~x21 && x3 && ~x15 && ~x16 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s390;
						end
					else if( ~x21 && ~x3 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s121;
						end
					else nx_state = s132;
				s133 : if( x65 && x66 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x66 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x66 && x20 && ~x17 )
						nx_state = s1;
					else if( x65 && x66 && ~x20 && x15 && x10 && x11 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s192;
						end
					else if( x65 && x66 && ~x20 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s193;
						end
					else if( x65 && x66 && ~x20 && x15 && x10 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y13 = 1'b1;	
							nx_state = s192;
						end
					else if( x65 && x66 && ~x20 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s300;
						end
					else if( x65 && x66 && ~x20 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s192;
						end
					else if( x65 && x66 && ~x20 && ~x15 && x16 && x10 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s306;
						end
					else if( x65 && x66 && ~x20 && ~x15 && x16 && ~x10 && x12 && x11 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s259;
						end
					else if( x65 && x66 && ~x20 && ~x15 && x16 && ~x10 && x12 && ~x11 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s306;
						end
					else if( x65 && x66 && ~x20 && ~x15 && x16 && ~x10 && ~x12 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s306;
						end
					else if( x65 && x66 && ~x20 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s201;
						end
					else if( x65 && ~x66 && x21 && x68 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x65 && ~x66 && x21 && ~x68 && x7 && x16 && x13 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && x21 && ~x68 && x7 && x16 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && x21 && ~x68 && x7 && ~x16 && x17 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && x21 && ~x68 && x7 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && x21 && ~x68 && ~x7 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x68 && x8 && x23 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x68 && x8 && x23 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x68 && x8 && x23 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && x68 && x8 && ~x23 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x68 && x8 && ~x23 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x68 && x8 && ~x23 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && x68 && ~x8 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && x16 && x18 && x19 && x10 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && x16 && x18 && x19 && ~x10 && x7 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && x16 && x18 && x19 && ~x10 && ~x7 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && x16 && x18 && ~x19 && x7 && x13 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && x16 && x18 && ~x19 && x7 && ~x13 )
						begin
							y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && x16 && x18 && ~x19 && ~x7 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && x16 && ~x18 && x13 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && x16 && ~x18 && ~x13 && x7 && x19 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s362;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && x16 && ~x18 && ~x13 && x7 && ~x19 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && x16 && ~x18 && ~x13 && ~x7 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && x10 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && x15 && x12 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && x15 && ~x12 && x14 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && x15 && ~x12 && ~x14 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && x15 && ~x12 && ~x14 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && x15 && ~x12 && ~x14 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && x15 && ~x12 && ~x14 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && ~x15 && x14 && x13 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && ~x15 && x14 && ~x13 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && ~x15 && x14 && ~x13 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && ~x15 && x14 && ~x13 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && ~x15 && x14 && ~x13 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && ~x15 && ~x14 && x11 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && ~x15 && ~x14 && ~x11 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && ~x15 && ~x14 && ~x11 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && ~x15 && ~x14 && ~x11 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && x19 && ~x10 && ~x15 && ~x14 && ~x11 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && ~x19 && x7 && x13 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && ~x19 && x7 && ~x13 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && x18 && ~x19 && ~x7 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && x13 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && x15 && x11 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && x15 && ~x11 && x14 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && x15 && ~x11 && ~x14 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && x15 && ~x11 && ~x14 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && x15 && ~x11 && ~x14 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && x15 && ~x11 && ~x14 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && x14 && x12 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && x14 && ~x12 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && x14 && ~x12 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && x14 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && x14 && ~x12 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && ~x14 && x10 && x19 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && ~x14 && x10 && ~x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && ~x14 && x10 && ~x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && ~x14 && x10 && ~x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && ~x14 && x10 && ~x19 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && ~x14 && ~x10 && x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && ~x14 && ~x10 && x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && ~x14 && ~x10 && x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && ~x14 && ~x10 && x19 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && x17 && ~x18 && ~x13 && ~x15 && ~x14 && ~x10 && ~x19 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && ~x17 && x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x68 && ~x16 && ~x17 && ~x7 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && x68 && x23 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && x68 && x23 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && x68 && x23 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x22 && x68 && x23 && ~x9 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x22 && x68 && ~x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && x68 && ~x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && x68 && ~x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x22 && x68 && ~x23 && ~x8 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && x17 && x13 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && x17 && ~x13 && x7 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s362;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && x17 && ~x13 && ~x7 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && x13 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && x15 && x11 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && x15 && ~x11 && x14 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && x15 && ~x11 && ~x14 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && x15 && ~x11 && ~x14 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && x15 && ~x11 && ~x14 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && x15 && ~x11 && ~x14 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && ~x15 && x14 && x12 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && ~x15 && x14 && ~x12 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && ~x15 && x14 && ~x12 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && ~x15 && x14 && ~x12 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && ~x15 && x14 && ~x12 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && ~x15 && ~x14 && x10 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && ~x15 && ~x14 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && ~x15 && ~x14 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && ~x15 && ~x14 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && x18 && ~x13 && ~x15 && ~x14 && ~x10 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && ~x18 && x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && x19 && ~x17 && ~x18 && ~x7 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && ~x19 && x16 && x13 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && ~x19 && x16 && ~x13 && x7 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && ~x19 && x16 && ~x13 && ~x7 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && ~x19 && ~x16 && x17 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && ~x19 && ~x16 && ~x17 && x7 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s146;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x68 && ~x19 && ~x16 && ~x17 && ~x7 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y14 = 1'b1;	
							nx_state = s391;
						end
					else if( ~x65 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x20 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x20 && x21 && x15 && x16 && x14 && x8 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s126;
						end
					else if( ~x65 && ~x20 && x21 && x15 && x16 && x14 && ~x8 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	y20 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x65 && ~x20 && x21 && x15 && x16 && ~x14 && x7 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s210;
						end
					else if( ~x65 && ~x20 && x21 && x15 && x16 && ~x14 && x7 && ~x8 )
						begin
							y7 = 1'b1;	y12 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x65 && ~x20 && x21 && x15 && x16 && ~x14 && ~x7 && x8 && x12 )
						begin
							y17 = 1'b1;	
							nx_state = s279;
						end
					else if( ~x65 && ~x20 && x21 && x15 && x16 && ~x14 && ~x7 && x8 && ~x12 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x20 && x21 && x15 && x16 && ~x14 && ~x7 && x8 && ~x12 && x18 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x20 && x21 && x15 && x16 && ~x14 && ~x7 && x8 && ~x12 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x20 && x21 && x15 && x16 && ~x14 && ~x7 && ~x8 && x13 )
						begin
							y17 = 1'b1;	
							nx_state = s279;
						end
					else if( ~x65 && ~x20 && x21 && x15 && x16 && ~x14 && ~x7 && ~x8 && ~x13 && x18 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x20 && x21 && x15 && x16 && ~x14 && ~x7 && ~x8 && ~x13 && x18 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x20 && x21 && x15 && x16 && ~x14 && ~x7 && ~x8 && ~x13 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x20 && x21 && x15 && ~x16 && x7 && x8 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x65 && ~x20 && x21 && x15 && ~x16 && x7 && ~x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && ~x20 && x21 && x15 && ~x16 && ~x7 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s392;
						end
					else if( ~x65 && ~x20 && x21 && x15 && ~x16 && ~x7 && ~x2 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x65 && ~x20 && x21 && x15 && ~x16 && ~x7 && ~x2 && ~x3 && x8 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x20 && x21 && x15 && ~x16 && ~x7 && ~x2 && ~x3 && ~x8 )
						begin
							y2 = 1'b1;	y13 = 1'b1;	
							nx_state = s206;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && x2 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s392;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && x7 && x11 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && x7 && x11 && ~x3 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && x7 && ~x11 && x8 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && x7 && ~x11 && x8 && ~x3 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && x7 && ~x11 && ~x8 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && x7 && ~x11 && ~x8 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && x7 && ~x11 && ~x8 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && x7 && ~x11 && ~x8 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && x8 && x9 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && x8 && x9 && ~x3 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && x8 && ~x9 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && x8 && ~x9 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && x8 && ~x9 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && x8 && ~x9 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && x10 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && x10 && ~x3 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && ~x10 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && ~x10 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && ~x10 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && x16 && ~x7 && ~x8 && ~x10 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && ~x16 && x3 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y7 = 1'b1;	
							nx_state = s41;
						end
					else if( ~x65 && ~x20 && x21 && ~x15 && ~x2 && ~x16 && ~x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s393;
						end
					else if( ~x65 && ~x20 && ~x21 && x6 && x15 && x8 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s366;
						end
					else if( ~x65 && ~x20 && ~x21 && x6 && x15 && ~x8 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s207;
						end
					else if( ~x65 && ~x20 && ~x21 && x6 && ~x15 && x16 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s366;
						end
					else if( ~x65 && ~x20 && ~x21 && x6 && ~x15 && ~x16 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s393;
						end
					else if( ~x65 && ~x20 && ~x21 && ~x6 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s366;
						end
					else nx_state = s133;
				s134 : if( x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( ~x21 && x15 && x10 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x21 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s301;
						end
					else if( ~x21 && x15 && x10 && ~x11 && ~x12 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s195;
						end
					else if( ~x21 && x15 && ~x10 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x21 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x21 && ~x15 && x16 && x10 && x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y11 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x21 && ~x15 && x16 && x10 && ~x12 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x21 && ~x15 && x16 && ~x10 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y11 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x21 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s303;
						end
					else nx_state = s134;
				s135 : if( x62 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s159;
						end
					else if( ~x62 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else nx_state = s135;
				s136 : if( x21 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && x18 && x19 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x21 && x22 && ~x23 && x18 && x19 && x15 && ~x17 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x21 && x22 && ~x23 && x18 && x19 && ~x15 && x16 && x17 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x21 && x22 && ~x23 && x18 && x19 && ~x15 && x16 && ~x17 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y20 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x21 && x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && x8 && x9 && x17 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && x8 && x9 && ~x17 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s117;
						end
					else if( ~x21 && x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && x8 && ~x9 && x10 && x17 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s117;
						end
					else if( ~x21 && x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && x8 && ~x9 && x10 && ~x17 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && x18 && x19 && ~x15 && ~x16 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && x18 && ~x19 && x16 && x15 )
						begin
							y18 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x21 && x22 && ~x23 && x18 && ~x19 && x16 && ~x15 && x17 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x21 && x22 && ~x23 && x18 && ~x19 && x16 && ~x15 && ~x17 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s233;
						end
					else if( ~x21 && x22 && ~x23 && x18 && ~x19 && ~x16 && x17 && x15 )
						begin
							y18 = 1'b1;	
							nx_state = s234;
						end
					else if( ~x21 && x22 && ~x23 && x18 && ~x19 && ~x16 && x17 && ~x15 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s235;
						end
					else if( ~x21 && x22 && ~x23 && x18 && ~x19 && ~x16 && ~x17 && x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s31;
						end
					else if( ~x21 && x22 && ~x23 && x18 && ~x19 && ~x16 && ~x17 && ~x5 && x3 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x21 && x22 && ~x23 && x18 && ~x19 && ~x16 && ~x17 && ~x5 && ~x3 && x15 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x21 && x22 && ~x23 && x18 && ~x19 && ~x16 && ~x17 && ~x5 && ~x3 && ~x15 )
						begin
							y16 = 1'b1;	y20 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && x15 && x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s31;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && x15 && ~x5 && x3 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && x15 && ~x5 && ~x3 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s228;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && x16 && x14 && x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s31;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && x16 && x14 && ~x5 && x3 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && x16 && x14 && ~x5 && ~x3 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && x16 && ~x14 && x17 && x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s31;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && x16 && ~x14 && x17 && ~x5 && x3 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && x16 && ~x14 && x17 && ~x5 && ~x3 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && x16 && ~x14 && ~x17 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && ~x16 && x17 && x13 && x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s31;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && ~x16 && x17 && x13 && ~x5 && x3 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && ~x16 && x17 && x13 && ~x5 && ~x3 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && ~x16 && x17 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && ~x16 && ~x17 && x12 && x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s31;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && ~x16 && ~x17 && x12 && ~x5 && x3 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && ~x16 && ~x17 && x12 && ~x5 && ~x3 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && x19 && ~x15 && ~x16 && ~x17 && ~x12 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && ~x18 && ~x19 && x5 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s31;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && ~x19 && ~x5 && x3 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s36;
						end
					else if( ~x21 && x22 && ~x23 && ~x18 && ~x19 && ~x5 && ~x3 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x21 && ~x22 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s161;
						end
					else nx_state = s136;
				s137 : if( x21 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x21 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x21 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x21 && ~x9 )
						nx_state = s1;
					else if( ~x21 && x22 )
						nx_state = s1;
					else if( ~x21 && ~x22 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else nx_state = s137;
				s138 : if( x21 && x19 && x20 && x17 && x5 )
						begin
							y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s269;
						end
					else if( x21 && x19 && x20 && x17 && ~x5 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( x21 && x19 && x20 && x17 && ~x5 && x3 && ~x4 )
						nx_state = s1;
					else if( x21 && x19 && x20 && x17 && ~x5 && ~x3 )
						nx_state = s1;
					else if( x21 && x19 && x20 && ~x17 && x4 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s273;
						end
					else if( x21 && x19 && x20 && ~x17 && ~x4 && x3 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( x21 && x19 && x20 && ~x17 && ~x4 && x3 && ~x5 )
						nx_state = s1;
					else if( x21 && x19 && x20 && ~x17 && ~x4 && ~x3 )
						nx_state = s1;
					else if( x21 && x19 && ~x20 && x12 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( x21 && x19 && ~x20 && x12 && ~x2 && x17 && x8 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && x19 && ~x20 && x12 && ~x2 && x17 && ~x8 )
						begin
							y18 = 1'b1;	
							nx_state = s272;
						end
					else if( x21 && x19 && ~x20 && x12 && ~x2 && ~x17 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( x21 && x19 && ~x20 && x12 && ~x2 && ~x17 && ~x8 )
						begin
							y6 = 1'b1;	
							nx_state = s172;
						end
					else if( x21 && x19 && ~x20 && ~x12 && x16 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x21 && x19 && ~x20 && ~x12 && ~x16 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s62;
						end
					else if( x21 && x19 && ~x20 && ~x12 && ~x16 && ~x2 && x8 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && x19 && ~x20 && ~x12 && ~x16 && ~x2 && ~x8 && x17 )
						begin
							y18 = 1'b1;	
							nx_state = s234;
						end
					else if( x21 && x19 && ~x20 && ~x12 && ~x16 && ~x2 && ~x8 && ~x17 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s374;
						end
					else if( x21 && ~x19 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s328;
						end
					else if( x21 && ~x19 && ~x2 && x20 && x12 && x8 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && ~x19 && ~x2 && x20 && x12 && ~x8 )
						begin
							y18 = 1'b1;	
							nx_state = s272;
						end
					else if( x21 && ~x19 && ~x2 && x20 && ~x12 && x17 && x16 && x8 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && ~x19 && ~x2 && x20 && ~x12 && x17 && x16 && ~x8 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s273;
						end
					else if( x21 && ~x19 && ~x2 && x20 && ~x12 && x17 && ~x16 && x14 && x8 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && ~x19 && ~x2 && x20 && ~x12 && x17 && ~x16 && x14 && ~x8 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s273;
						end
					else if( x21 && ~x19 && ~x2 && x20 && ~x12 && x17 && ~x16 && ~x14 )
						nx_state = s1;
					else if( x21 && ~x19 && ~x2 && x20 && ~x12 && ~x17 && x16 && x15 && x8 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && ~x19 && ~x2 && x20 && ~x12 && ~x17 && x16 && x15 && ~x8 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s273;
						end
					else if( x21 && ~x19 && ~x2 && x20 && ~x12 && ~x17 && x16 && ~x15 )
						nx_state = s1;
					else if( x21 && ~x19 && ~x2 && x20 && ~x12 && ~x17 && ~x16 && x13 && x8 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && ~x19 && ~x2 && x20 && ~x12 && ~x17 && ~x16 && x13 && ~x8 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	
							nx_state = s273;
						end
					else if( x21 && ~x19 && ~x2 && x20 && ~x12 && ~x17 && ~x16 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x19 && ~x2 && ~x20 && x8 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( x21 && ~x19 && ~x2 && ~x20 && ~x8 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s394;
						end
					else if( x21 && ~x19 && ~x2 && ~x20 && ~x8 && ~x12 )
						begin
							y18 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x21 && x22 )
						nx_state = s1;
					else if( ~x21 && ~x22 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else nx_state = s138;
				s139 : if( 1'b1 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else nx_state = s139;
				s140 : if( x65 && x66 && x68 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x65 && x66 && ~x68 && x60 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && x62 && x20 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	
							nx_state = s367;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && x62 && ~x20 && x16 && x11 && x12 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && x62 && ~x20 && x16 && x11 && ~x12 && x13 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s153;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && x62 && ~x20 && x16 && x11 && ~x12 && ~x13 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s154;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && x62 && ~x20 && x16 && ~x11 && x13 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s63;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && x62 && ~x20 && x16 && ~x11 && ~x13 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && x62 && ~x20 && ~x16 && x17 && x11 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && x62 && ~x20 && ~x16 && x17 && x11 && ~x13 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && x62 && ~x20 && ~x16 && x17 && ~x11 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && x62 && ~x20 && ~x16 && ~x17 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( x65 && x66 && ~x68 && ~x60 && x61 && ~x62 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x65 && x66 && ~x68 && ~x60 && ~x61 )
						begin
							y2 = 1'b1;	y19 = 1'b1;	y24 = 1'b1;	
							nx_state = s321;
						end
					else if( x65 && ~x66 && x67 && x21 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x65 && ~x66 && x67 && x21 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x65 && ~x66 && x67 && x21 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && x21 && ~x8 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && ~x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s32;
						end
					else if( x65 && ~x66 && ~x67 && x20 && x19 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x20 && x19 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x20 && x19 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x20 && x19 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x20 && ~x19 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	y25 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && ~x66 && ~x67 && ~x20 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	y25 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x65 && x67 && x68 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && x67 && x68 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && x67 && x68 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && x67 && x68 && x21 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x67 && x68 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x65 && x67 && x68 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x65 && x67 && x68 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && x67 && x68 && ~x21 && ~x20 )
						nx_state = s1;
					else if( ~x65 && x67 && ~x68 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && x67 && ~x68 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && x67 && ~x68 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x67 && ~x68 && x62 && ~x61 )
						nx_state = s1;
					else if( ~x65 && x67 && ~x68 && ~x62 && x63 && x17 && x13 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && x67 && ~x68 && ~x62 && x63 && x17 && ~x13 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && x67 && ~x68 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x67 && ~x68 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( ~x65 && x67 && ~x68 && ~x62 && ~x63 && x64 && x4 )
						begin
							y31 = 1'b1;	
							nx_state = s96;
						end
					else if( ~x65 && x67 && ~x68 && ~x62 && ~x63 && x64 && ~x4 && x18 && x16 && x8 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && x67 && ~x68 && ~x62 && ~x63 && x64 && ~x4 && x18 && x16 && ~x8 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && x67 && ~x68 && ~x62 && ~x63 && x64 && ~x4 && x18 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x65 && x67 && ~x68 && ~x62 && ~x63 && x64 && ~x4 && ~x18 )
						begin
							y14 = 1'b1;	y28 = 1'b1;	y32 = 1'b1;	
							y33 = 1'b1;	
							nx_state = s18;
						end
					else if( ~x65 && x67 && ~x68 && ~x62 && ~x63 && ~x64 && x19 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x67 && ~x68 && ~x62 && ~x63 && ~x64 && x19 && ~x13 && x12 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x67 && ~x68 && ~x62 && ~x63 && ~x64 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x67 && ~x68 && ~x62 && ~x63 && ~x64 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x67 && x21 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s143;
						end
					else if( ~x65 && ~x67 && ~x21 && x23 && x22 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x65 && ~x67 && ~x21 && x23 && ~x22 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x65 && ~x67 && ~x21 && x23 && ~x22 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x65 && ~x67 && ~x21 && x23 && ~x22 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && x23 && ~x22 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else nx_state = s140;
				s141 : if( x21 && x20 && x16 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s113;
						end
					else if( x21 && x20 && x16 && ~x10 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x21 && x20 && ~x16 && x17 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x21 && x20 && ~x16 && ~x17 )
						begin
							y5 = 1'b1;	y17 = 1'b1;	
							nx_state = s115;
						end
					else if( x21 && ~x20 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s317;
						end
					else if( ~x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s317;
						end
					else nx_state = s141;
				s142 : if( x66 && x16 && x17 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && x16 && x17 && x8 && ~x10 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x66 && x16 && x17 && ~x8 && x9 && x10 )
						begin
							y23 = 1'b1;	y24 = 1'b1;	
							nx_state = s269;
						end
					else if( x66 && x16 && x17 && ~x8 && x9 && ~x10 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y15 = 1'b1;	
							y18 = 1'b1;	y25 = 1'b1;	
							nx_state = s113;
						end
					else if( x66 && x16 && x17 && ~x8 && ~x9 && x21 && x10 && x14 )
						begin
							y6 = 1'b1;	
							nx_state = s188;
						end
					else if( x66 && x16 && x17 && ~x8 && ~x9 && x21 && x10 && ~x14 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && x16 && x17 && ~x8 && ~x9 && x21 && x10 && ~x14 && x19 && ~x15 )
						nx_state = s1;
					else if( x66 && x16 && x17 && ~x8 && ~x9 && x21 && x10 && ~x14 && ~x19 )
						nx_state = s1;
					else if( x66 && x16 && x17 && ~x8 && ~x9 && x21 && ~x10 && x15 )
						begin
							y6 = 1'b1;	
							nx_state = s188;
						end
					else if( x66 && x16 && x17 && ~x8 && ~x9 && x21 && ~x10 && ~x15 && x19 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && x16 && x17 && ~x8 && ~x9 && x21 && ~x10 && ~x15 && x19 && ~x14 )
						nx_state = s1;
					else if( x66 && x16 && x17 && ~x8 && ~x9 && x21 && ~x10 && ~x15 && ~x19 )
						nx_state = s1;
					else if( x66 && x16 && x17 && ~x8 && ~x9 && ~x21 && x10 && x14 )
						begin
							y6 = 1'b1;	
							nx_state = s188;
						end
					else if( x66 && x16 && x17 && ~x8 && ~x9 && ~x21 && x10 && ~x14 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x66 && x16 && x17 && ~x8 && ~x9 && ~x21 && x10 && ~x14 && x20 && ~x15 )
						nx_state = s1;
					else if( x66 && x16 && x17 && ~x8 && ~x9 && ~x21 && x10 && ~x14 && ~x20 )
						nx_state = s1;
					else if( x66 && x16 && x17 && ~x8 && ~x9 && ~x21 && ~x10 && x15 )
						begin
							y6 = 1'b1;	
							nx_state = s188;
						end
					else if( x66 && x16 && x17 && ~x8 && ~x9 && ~x21 && ~x10 && ~x15 && x20 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x66 && x16 && x17 && ~x8 && ~x9 && ~x21 && ~x10 && ~x15 && x20 && ~x14 )
						nx_state = s1;
					else if( x66 && x16 && x17 && ~x8 && ~x9 && ~x21 && ~x10 && ~x15 && ~x20 )
						nx_state = s1;
					else if( x66 && x16 && ~x17 && x9 && x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s344;
						end
					else if( x66 && x16 && ~x17 && x9 && ~x21 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( x66 && x16 && ~x17 && ~x9 && x8 && x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s344;
						end
					else if( x66 && x16 && ~x17 && ~x9 && x8 && ~x21 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( x66 && x16 && ~x17 && ~x9 && ~x8 && x2 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( x66 && x16 && ~x17 && ~x9 && ~x8 && ~x2 && x21 && x3 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x66 && x16 && ~x17 && ~x9 && ~x8 && ~x2 && x21 && ~x3 && x10 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x66 && x16 && ~x17 && ~x9 && ~x8 && ~x2 && x21 && ~x3 && ~x10 )
						begin
							y4 = 1'b1;	y18 = 1'b1;	
							nx_state = s395;
						end
					else if( x66 && x16 && ~x17 && ~x9 && ~x8 && ~x2 && ~x21 && x3 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && x16 && ~x17 && ~x9 && ~x8 && ~x2 && ~x21 && ~x3 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s113;
						end
					else if( x66 && x16 && ~x17 && ~x9 && ~x8 && ~x2 && ~x21 && ~x3 && ~x10 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x66 && ~x16 && x2 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( x66 && ~x16 && ~x2 && x17 && x10 && x11 )
						begin
							y7 = 1'b1;	y12 = 1'b1;	
							nx_state = s211;
						end
					else if( x66 && ~x16 && ~x2 && x17 && x10 && ~x11 && x9 )
						begin
							y7 = 1'b1;	y12 = 1'b1;	
							nx_state = s211;
						end
					else if( x66 && ~x16 && ~x2 && x17 && x10 && ~x11 && ~x9 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && ~x16 && ~x2 && x17 && x10 && ~x11 && ~x9 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && ~x16 && ~x2 && x17 && x10 && ~x11 && ~x9 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x66 && ~x16 && ~x2 && x17 && x10 && ~x11 && ~x9 && x21 && ~x19 )
						nx_state = s1;
					else if( x66 && ~x16 && ~x2 && x17 && x10 && ~x11 && ~x9 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x66 && ~x16 && ~x2 && x17 && x10 && ~x11 && ~x9 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x66 && ~x16 && ~x2 && x17 && x10 && ~x11 && ~x9 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x66 && ~x16 && ~x2 && x17 && x10 && ~x11 && ~x9 && ~x21 && ~x20 )
						nx_state = s1;
					else if( x66 && ~x16 && ~x2 && x17 && ~x10 && x9 && x13 )
						begin
							y7 = 1'b1;	y12 = 1'b1;	
							nx_state = s211;
						end
					else if( x66 && ~x16 && ~x2 && x17 && ~x10 && x9 && ~x13 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && ~x16 && ~x2 && x17 && ~x10 && x9 && ~x13 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && ~x16 && ~x2 && x17 && ~x10 && x9 && ~x13 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x66 && ~x16 && ~x2 && x17 && ~x10 && x9 && ~x13 && x21 && ~x19 )
						nx_state = s1;
					else if( x66 && ~x16 && ~x2 && x17 && ~x10 && x9 && ~x13 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x66 && ~x16 && ~x2 && x17 && ~x10 && x9 && ~x13 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x66 && ~x16 && ~x2 && x17 && ~x10 && x9 && ~x13 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x66 && ~x16 && ~x2 && x17 && ~x10 && x9 && ~x13 && ~x21 && ~x20 )
						nx_state = s1;
					else if( x66 && ~x16 && ~x2 && x17 && ~x10 && ~x9 && x12 )
						begin
							y7 = 1'b1;	y12 = 1'b1;	
							nx_state = s211;
						end
					else if( x66 && ~x16 && ~x2 && x17 && ~x10 && ~x9 && ~x12 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && ~x16 && ~x2 && x17 && ~x10 && ~x9 && ~x12 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && ~x16 && ~x2 && x17 && ~x10 && ~x9 && ~x12 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x66 && ~x16 && ~x2 && x17 && ~x10 && ~x9 && ~x12 && x21 && ~x19 )
						nx_state = s1;
					else if( x66 && ~x16 && ~x2 && x17 && ~x10 && ~x9 && ~x12 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x66 && ~x16 && ~x2 && x17 && ~x10 && ~x9 && ~x12 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x66 && ~x16 && ~x2 && x17 && ~x10 && ~x9 && ~x12 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x66 && ~x16 && ~x2 && x17 && ~x10 && ~x9 && ~x12 && ~x21 && ~x20 )
						nx_state = s1;
					else if( x66 && ~x16 && ~x2 && ~x17 && x3 && x21 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x66 && ~x16 && ~x2 && ~x17 && x3 && ~x21 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && ~x16 && ~x2 && ~x17 && ~x3 )
						begin
							y17 = 1'b1;	
							nx_state = s279;
						end
					else if( ~x66 && x21 && x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s328;
						end
					else if( ~x66 && x21 && ~x19 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s396;
						end
					else if( ~x66 && ~x21 && x22 && x18 && x17 && x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x66 && ~x21 && x22 && x18 && x17 && ~x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x66 && ~x21 && x22 && x18 && ~x17 && x12 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s386;
						end
					else if( ~x66 && ~x21 && x22 && x18 && ~x17 && ~x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s374;
						end
					else if( ~x66 && ~x21 && x22 && ~x18 && x19 && x12 && x17 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x66 && ~x21 && x22 && ~x18 && x19 && x12 && ~x17 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x66 && ~x21 && x22 && ~x18 && x19 && ~x12 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x66 && ~x21 && x22 && ~x18 && ~x19 && x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x66 && ~x21 && x22 && ~x18 && ~x19 && ~x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x66 && ~x21 && ~x22 )
						nx_state = s1;
					else nx_state = s142;
				s143 : if( x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x18 )
						nx_state = s1;
					else if( ~x21 && x23 && x15 && x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x21 && x23 && x15 && ~x10 && x12 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && x23 && x15 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s285;
						end
					else if( ~x21 && x23 && ~x15 && x16 && x10 && x12 )
						begin
							y14 = 1'b1;	
							nx_state = s286;
						end
					else if( ~x21 && x23 && ~x15 && x16 && x10 && ~x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x21 && x23 && ~x15 && x16 && ~x10 )
						begin
							y14 = 1'b1;	
							nx_state = s286;
						end
					else if( ~x21 && x23 && ~x15 && ~x16 )
						nx_state = s40;
					else if( ~x21 && ~x23 && x15 && x10 && x11 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s334;
						end
					else if( ~x21 && ~x23 && x15 && x10 && ~x11 && x12 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s334;
						end
					else if( ~x21 && ~x23 && x15 && x10 && ~x11 && ~x12 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x21 && ~x23 && x15 && ~x10 && x12 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x21 && ~x23 && x15 && ~x10 && x12 && ~x11 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && ~x23 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x21 && ~x23 && ~x15 && x16 && x10 && x12 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x21 && ~x23 && ~x15 && x16 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s341;
						end
					else if( ~x21 && ~x23 && ~x15 && x16 && ~x10 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x21 && ~x23 && ~x15 && ~x16 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s81;
						end
					else nx_state = s143;
				s144 : if( x65 && x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x65 && x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x66 && x21 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x21 && x22 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && x66 && ~x21 && x22 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && x66 && ~x21 && x22 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x21 && x22 && x23 && ~x17 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x21 && x22 && ~x23 && x19 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s304;
						end
					else if( ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && x20 && x15 && x10 && x11 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s334;
						end
					else if( ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && x20 && x15 && x10 && ~x11 && x12 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s334;
						end
					else if( ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && x20 && x15 && x10 && ~x11 && ~x12 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && x20 && x15 && ~x10 && x12 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && x20 && x15 && ~x10 && x12 && ~x11 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && x20 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && x20 && ~x15 && x16 && x10 && x12 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && x20 && ~x15 && x16 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s341;
						end
					else if( ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && x20 && ~x15 && x16 && ~x10 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && x20 && ~x15 && ~x16 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s81;
						end
					else if( ~x65 && x66 && ~x21 && x22 && ~x23 && ~x19 && ~x20 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && x23 && x3 )
						begin
							y3 = 1'b1;	
							nx_state = s320;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && x23 && ~x3 && x18 && x15 && x7 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s81;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && x23 && ~x3 && x18 && x15 && ~x7 && x9 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && x23 && ~x3 && x18 && x15 && ~x7 && ~x9 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && x23 && ~x3 && x18 && ~x15 && x7 && x9 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s330;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && x23 && ~x3 && x18 && ~x15 && x7 && ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && x23 && ~x3 && x18 && ~x15 && ~x7 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s330;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && x23 && ~x3 && ~x18 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s84;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && ~x23 && x15 && x7 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s81;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && ~x23 && x15 && ~x7 && x9 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s370;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && ~x23 && x15 && ~x7 && ~x9 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && ~x23 && ~x15 && x7 && x9 )
						begin
							y3 = 1'b1;	
							nx_state = s320;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && ~x23 && ~x15 && x7 && ~x9 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s333;
						end
					else if( ~x65 && x66 && ~x21 && ~x22 && ~x23 && ~x15 && ~x7 )
						begin
							y3 = 1'b1;	
							nx_state = s320;
						end
					else if( ~x65 && ~x66 && x24 && x26 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x66 && x24 && x26 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && ~x66 && x24 && x26 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x24 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x24 && ~x26 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x26 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x26 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x66 && ~x24 && x25 && x26 && x19 && ~x14 && ~x13 )
						nx_state = s144;
					else if( ~x65 && ~x66 && ~x24 && x25 && x26 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x24 && x25 && ~x26 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x65 && ~x66 && ~x24 && ~x25 && x26 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && ~x66 && ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x65 && ~x66 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x65 && ~x66 && ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else nx_state = s144;
				s145 : if( x21 && x15 && x10 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s330;
						end
					else if( x21 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x21 && x15 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s48;
						end
					else if( x21 && ~x15 && x16 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x21 && ~x15 && ~x16 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s340;
						end
					else if( ~x21 && x22 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s143;
						end
					else if( ~x21 && ~x22 )
						nx_state = s1;
					else nx_state = s145;
				s146 : if( x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x4 )
						nx_state = s1;
					else nx_state = s146;
				s147 : if( x21 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && x23 && x22 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && x23 && ~x22 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( ~x21 && x23 && ~x22 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( ~x21 && x23 && ~x22 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x23 && ~x22 && ~x20 )
						nx_state = s1;
					else if( ~x21 && ~x23 && x18 && x14 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( ~x21 && ~x23 && x18 && x14 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && ~x23 && x18 && ~x14 && x13 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( ~x21 && ~x23 && x18 && ~x14 && x13 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x23 && ~x18 )
						nx_state = s1;
					else nx_state = s147;
				s148 : if( x20 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x20 && x21 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x20 && ~x21 )
						nx_state = s1;
					else nx_state = s148;
				s149 : if( x66 && x65 && x61 && x60 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && x65 && x61 && x60 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x66 && x65 && x61 && x60 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x66 && x65 && x61 && x60 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x66 && x65 && x61 && ~x60 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x66 && x65 && x61 && ~x60 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x66 && x65 && x61 && ~x60 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x66 && x65 && x61 && ~x60 && x62 && ~x18 )
						nx_state = s1;
					else if( x66 && x65 && x61 && ~x60 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && x65 && x61 && ~x60 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && x65 && x61 && ~x60 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x66 && x65 && x61 && ~x60 && ~x62 && ~x18 )
						nx_state = s39;
					else if( x66 && x65 && ~x61 && x60 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && x65 && ~x61 && x60 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && x65 && ~x61 && x60 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x66 && x65 && ~x61 && x60 && ~x18 )
						nx_state = s39;
					else if( x66 && x65 && ~x61 && ~x60 && x62 && x11 && x10 && x15 )
						nx_state = s40;
					else if( x66 && x65 && ~x61 && ~x60 && x62 && x11 && x10 && ~x15 && x7 )
						nx_state = s40;
					else if( x66 && x65 && ~x61 && ~x60 && x62 && x11 && x10 && ~x15 && ~x7 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( x66 && x65 && ~x61 && ~x60 && x62 && x11 && ~x10 )
						nx_state = s40;
					else if( x66 && x65 && ~x61 && ~x60 && x62 && ~x11 && x12 && x9 && x15 )
						nx_state = s40;
					else if( x66 && x65 && ~x61 && ~x60 && x62 && ~x11 && x12 && x9 && ~x15 && x7 )
						nx_state = s40;
					else if( x66 && x65 && ~x61 && ~x60 && x62 && ~x11 && x12 && x9 && ~x15 && ~x7 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( x66 && x65 && ~x61 && ~x60 && x62 && ~x11 && x12 && ~x9 )
						nx_state = s40;
					else if( x66 && x65 && ~x61 && ~x60 && x62 && ~x11 && ~x12 && x8 && x15 )
						nx_state = s40;
					else if( x66 && x65 && ~x61 && ~x60 && x62 && ~x11 && ~x12 && x8 && ~x15 && x7 )
						nx_state = s40;
					else if( x66 && x65 && ~x61 && ~x60 && x62 && ~x11 && ~x12 && x8 && ~x15 && ~x7 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( x66 && x65 && ~x61 && ~x60 && x62 && ~x11 && ~x12 && ~x8 )
						nx_state = s40;
					else if( x66 && x65 && ~x61 && ~x60 && ~x62 )
						nx_state = s40;
					else if( x66 && ~x65 && x67 && x62 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s159;
						end
					else if( x66 && ~x65 && x67 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && ~x65 && x67 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( x66 && ~x65 && x67 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && ~x65 && x67 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( x66 && ~x65 && x67 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x66 && ~x65 && x67 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( x66 && ~x65 && x67 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x66 && ~x65 && x67 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x66 && ~x65 && x67 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x66 && ~x65 && x67 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x66 && ~x65 && x67 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x66 && ~x65 && x67 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x66 && ~x65 && ~x67 && x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x66 && ~x65 && ~x67 && x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && x21 && ~x18 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && x23 && x22 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && x23 && x22 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && x23 && x22 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && x23 && x22 && ~x17 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && x23 && ~x22 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && x23 && ~x22 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( x66 && ~x65 && ~x67 && ~x21 && x23 && ~x22 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && x23 && ~x22 && ~x19 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x23 && x22 && x18 && x14 )
						nx_state = s40;
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x23 && x22 && x18 && ~x14 && x13 )
						nx_state = s40;
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x23 && x22 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x23 && x22 && ~x18 )
						nx_state = s1;
					else if( x66 && ~x65 && ~x67 && ~x21 && ~x23 && ~x22 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x66 && x65 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x66 && x65 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x66 && x65 && ~x4 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && x24 && x26 && x11 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x66 && ~x65 && x67 && x24 && x26 && ~x11 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x66 && ~x65 && x67 && x24 && x26 && ~x11 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x66 && ~x65 && x67 && x24 && x26 && ~x11 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && x24 && x26 && ~x11 && ~x18 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && x24 && ~x26 && x19 && x16 && x11 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x66 && ~x65 && x67 && x24 && ~x26 && x19 && x16 && x11 && ~x12 && x13 )
						begin
							y6 = 1'b1;	
							nx_state = s172;
						end
					else if( ~x66 && ~x65 && x67 && x24 && ~x26 && x19 && x16 && x11 && ~x12 && ~x13 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x66 && ~x65 && x67 && x24 && ~x26 && x19 && x16 && ~x11 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x66 && ~x65 && x67 && x24 && ~x26 && x19 && ~x16 && x17 && x11 && x13 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else if( ~x66 && ~x65 && x67 && x24 && ~x26 && x19 && ~x16 && x17 && x11 && ~x13 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s46;
						end
					else if( ~x66 && ~x65 && x67 && x24 && ~x26 && x19 && ~x16 && x17 && ~x11 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else if( ~x66 && ~x65 && x67 && x24 && ~x26 && x19 && ~x16 && ~x17 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && ~x65 && x67 && x24 && ~x26 && ~x19 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x66 && ~x65 && x67 && ~x24 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x66 && ~x65 && x67 && ~x24 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x66 && ~x65 && x67 && ~x24 && x25 && x19 && ~x14 && ~x13 && x26 )
						nx_state = s149;
					else if( ~x66 && ~x65 && x67 && ~x24 && x25 && x19 && ~x14 && ~x13 && ~x26 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && ~x24 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && x10 && x12 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && x10 && x12 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && x10 && x12 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && x10 && x12 && ~x18 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && x10 && ~x12 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s165;
						end
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && ~x10 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && ~x10 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && ~x10 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && x26 && ~x10 && ~x18 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && x10 && x12 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && x10 && x12 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && x10 && x12 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && x10 && x12 && ~x17 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && x10 && ~x12 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && ~x10 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && ~x10 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && ~x10 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x66 && ~x65 && x67 && ~x24 && ~x25 && ~x26 && ~x10 && ~x17 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x67 && x21 && x9 && x3 )
						nx_state = s40;
					else if( ~x66 && ~x65 && ~x67 && x21 && x9 && ~x3 && x4 )
						nx_state = s40;
					else if( ~x66 && ~x65 && ~x67 && x21 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x67 && x21 && ~x9 )
						nx_state = s1;
					else if( ~x66 && ~x65 && ~x67 && ~x21 )
						nx_state = s1;
					else nx_state = s149;
				s150 : if( 1'b1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else nx_state = s150;
				s151 : if( x66 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x66 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x66 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x66 && x62 && ~x61 )
						nx_state = s1;
					else if( x66 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( x66 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x66 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( x66 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x66 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( x66 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x66 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x66 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x66 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x66 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x66 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else if( ~x66 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s123;
						end
					else nx_state = s151;
				s152 : if( x64 && x63 )
						begin
							y3 = 1'b1;	y22 = 1'b1;	y37 = 1'b1;	
							nx_state = s397;
						end
					else if( x64 && ~x63 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s20;
						end
					else if( ~x64 && x63 )
						nx_state = s1;
					else if( ~x64 && ~x63 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else nx_state = s152;
				s153 : if( 1'b1 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else nx_state = s153;
				s154 : if( x67 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x67 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x67 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x67 && x22 && ~x17 )
						nx_state = s1;
					else if( x67 && ~x22 && x18 && x13 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x67 && ~x22 && x18 && x13 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x67 && ~x22 && x18 && ~x13 && x12 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x67 && ~x22 && x18 && ~x13 && x12 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x67 && ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x67 && ~x22 && ~x18 )
						nx_state = s1;
					else if( ~x67 && x61 && x60 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x67 && x61 && ~x60 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x67 && x61 && ~x60 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x67 && x61 && ~x60 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( ~x67 && x61 && ~x60 && x62 && ~x18 )
						nx_state = s1;
					else if( ~x67 && x61 && ~x60 && ~x62 && x15 )
						nx_state = s73;
					else if( ~x67 && x61 && ~x60 && ~x62 && ~x15 && x16 )
						begin
							y12 = 1'b1;	
							nx_state = s291;
						end
					else if( ~x67 && x61 && ~x60 && ~x62 && ~x15 && ~x16 )
						nx_state = s73;
					else if( ~x67 && ~x61 && x60 && x15 )
						nx_state = s73;
					else if( ~x67 && ~x61 && x60 && ~x15 && x16 )
						begin
							y12 = 1'b1;	
							nx_state = s291;
						end
					else if( ~x67 && ~x61 && x60 && ~x15 && ~x16 )
						nx_state = s73;
					else if( ~x67 && ~x61 && ~x60 && x62 )
						nx_state = s1;
					else if( ~x67 && ~x61 && ~x60 && ~x62 && x15 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x67 && ~x61 && ~x60 && ~x62 && x15 && ~x7 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x67 && ~x61 && ~x60 && ~x62 && x15 && ~x7 && ~x11 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && x4 )
						nx_state = s40;
					else if( ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && ~x4 && x11 && x9 )
						nx_state = s40;
					else if( ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && ~x4 && x11 && ~x9 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && ~x4 && x11 && ~x9 && ~x7 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s118;
						end
					else if( ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && ~x4 && ~x11 && x9 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && ~x4 && ~x11 && x9 && ~x7 && x10 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && ~x4 && ~x11 && x9 && ~x7 && ~x10 )
						nx_state = s40;
					else if( ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && x7 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && x7 && ~x8 )
						nx_state = s40;
					else if( ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && ~x7 && x12 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && ~x7 && ~x12 )
						nx_state = s40;
					else if( ~x67 && ~x61 && ~x60 && ~x62 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else nx_state = s154;
				s155 : if( x65 && x60 && x61 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s252;
						end
					else if( x65 && x60 && ~x61 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x60 && ~x61 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x60 && ~x61 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x65 && x60 && ~x61 && ~x18 )
						nx_state = s39;
					else if( x65 && ~x60 && x62 && x61 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x65 && ~x60 && x62 && ~x61 )
						nx_state = s316;
					else if( x65 && ~x60 && ~x62 && x61 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x60 && ~x62 && x61 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x60 && ~x62 && x61 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x65 && ~x60 && ~x62 && x61 && ~x18 )
						nx_state = s39;
					else if( x65 && ~x60 && ~x62 && ~x61 )
						nx_state = s40;
					else if( ~x65 && x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x65 && x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x65 && x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x21 && x22 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x21 && x22 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x23 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x23 && x18 && x14 )
						nx_state = s40;
					else if( ~x65 && ~x21 && x22 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s40;
					else if( ~x65 && ~x21 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x21 && ~x22 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s180;
						end
					else nx_state = s155;
				s156 : if( x63 && x64 && x18 && x15 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( x63 && x64 && x18 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x63 && x64 && x18 && ~x15 && x16 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( x63 && x64 && x18 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s135;
						end
					else if( x63 && x64 && ~x18 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s152;
						end
					else if( x63 && ~x64 )
						begin
							y19 = 1'b1;	
							nx_state = s213;
						end
					else if( ~x63 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else nx_state = s156;
				s157 : if( x65 && x21 && x67 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x65 && x21 && x67 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x65 && x21 && x67 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x65 && x21 && x67 && ~x8 )
						nx_state = s1;
					else if( x65 && x21 && ~x67 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x65 && x21 && ~x67 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x21 && ~x67 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x21 && ~x67 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x21 && ~x67 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x21 && x23 && x22 && x67 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && x23 && x22 && x67 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && x23 && x22 && x67 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && ~x21 && x23 && x22 && x67 && ~x8 )
						nx_state = s1;
					else if( x65 && ~x21 && x23 && x22 && ~x67 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( x65 && ~x21 && x23 && x22 && ~x67 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x21 && x23 && x22 && ~x67 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x21 && x23 && x22 && ~x67 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x21 && x23 && x22 && ~x67 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x21 && x23 && ~x22 && x67 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && x23 && ~x22 && x67 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && x23 && ~x22 && x67 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && ~x21 && x23 && ~x22 && x67 && ~x9 )
						nx_state = s1;
					else if( x65 && ~x21 && x23 && ~x22 && ~x67 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x21 && x23 && ~x22 && ~x67 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x21 && x23 && ~x22 && ~x67 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x21 && x23 && ~x22 && ~x67 && ~x20 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x23 && x67 && x8 && x22 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && ~x23 && x67 && x8 && x22 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && ~x23 && x67 && x8 && x22 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x23 && x67 && x8 && ~x22 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && ~x23 && x67 && x8 && ~x22 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && ~x23 && x67 && x8 && ~x22 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x23 && x67 && ~x8 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x23 && ~x67 && x18 && x14 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x21 && ~x23 && ~x67 && x18 && x14 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x21 && ~x23 && ~x67 && x18 && ~x14 && x13 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x21 && ~x23 && ~x67 && x18 && ~x14 && x13 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x21 && ~x23 && ~x67 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x23 && ~x67 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x62 && ~x61 )
						nx_state = s1;
					else if( ~x65 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else nx_state = s157;
				s158 : if( x65 && x21 && x18 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x65 && x21 && ~x18 && x19 && x14 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x21 && ~x18 && x19 && ~x14 && x13 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x21 && ~x18 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x21 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x21 && x23 && x22 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( x65 && ~x21 && x23 && x22 && ~x19 && x17 && x14 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && x13 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( x65 && ~x21 && x23 && x22 && ~x19 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x21 && x23 && x22 && ~x19 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x21 && x23 && ~x22 && x20 && x14 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x21 && x23 && ~x22 && x20 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( x65 && ~x21 && x23 && ~x22 && x20 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x21 && x23 && ~x22 && ~x20 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x23 && x18 && x14 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x21 && ~x23 && x18 && x14 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x21 && ~x23 && x18 && ~x14 && x13 && x22 )
						begin
							y37 = 1'b1;	
							nx_state = s120;
						end
					else if( x65 && ~x21 && ~x23 && x18 && ~x14 && x13 && ~x22 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x21 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x65 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x62 && ~x61 )
						nx_state = s1;
					else if( ~x65 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else nx_state = s158;
				s159 : if( x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x62 && ~x61 )
						nx_state = s1;
					else if( ~x62 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else nx_state = s159;
				s160 : if( x24 && x26 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( x24 && x26 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( x24 && x26 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x24 && x26 && ~x18 )
						nx_state = s1;
					else if( x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x24 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x25 && x19 && ~x14 && ~x13 && x26 )
						nx_state = s160;
					else if( ~x24 && x25 && x19 && ~x14 && ~x13 && ~x26 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else nx_state = s160;
				s161 : if( x65 && x21 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x65 && ~x21 && x22 && x8 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && x22 && x8 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && x22 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x65 && ~x21 && x22 && ~x8 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x22 && x23 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && ~x22 && x23 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && ~x22 && x23 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x22 && x23 && ~x9 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x22 && ~x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && ~x22 && ~x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x22 && ~x23 && ~x8 )
						nx_state = s1;
					else if( ~x65 && x24 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x65 && ~x24 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x24 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x65 && ~x24 && x19 && ~x14 && ~x13 )
						nx_state = s161;
					else if( ~x65 && ~x24 && ~x19 )
						nx_state = s1;
					else nx_state = s161;
				s162 : if( x24 && x26 )
						nx_state = s1;
					else if( x24 && ~x26 )
						begin
							y11 = 1'b1;	y16 = 1'b1;	y25 = 1'b1;	
							nx_state = s281;
						end
					else if( ~x24 && x25 && x15 && x10 && x11 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x24 && x25 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s398;
						end
					else if( ~x24 && x25 && x15 && x10 && ~x11 && ~x12 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x24 && x25 && x15 && ~x10 && x12 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s399;
						end
					else if( ~x24 && x25 && x15 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x24 && x25 && ~x15 && x16 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x24 && x25 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else if( ~x24 && ~x25 && x26 )
						begin
							y11 = 1'b1;	y16 = 1'b1;	y25 = 1'b1;	
							nx_state = s281;
						end
					else if( ~x24 && ~x25 && ~x26 && x18 && x15 && x12 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && ~x25 && ~x26 && x18 && x15 && ~x12 && x11 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && ~x25 && ~x26 && x18 && x15 && ~x12 && ~x11 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x24 && ~x25 && ~x26 && x18 && x15 && ~x12 && ~x11 && ~x10 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x24 && ~x25 && ~x26 && x18 && ~x15 && x16 && x10 && x12 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s282;
						end
					else if( ~x24 && ~x25 && ~x26 && x18 && ~x15 && x16 && x10 && ~x12 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s392;
						end
					else if( ~x24 && ~x25 && ~x26 && x18 && ~x15 && x16 && ~x10 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s282;
						end
					else if( ~x24 && ~x25 && ~x26 && x18 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x18 )
						begin
							y11 = 1'b1;	y16 = 1'b1;	y25 = 1'b1;	
							nx_state = s281;
						end
					else nx_state = s162;
				s163 : if( x65 )
						begin
							y15 = 1'b1;	y21 = 1'b1;	y28 = 1'b1;	
							nx_state = s313;
						end
					else if( ~x65 && x66 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x65 && ~x66 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else nx_state = s163;
				s164 : if( x24 && x26 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( x24 && x26 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( x24 && x26 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x24 && x26 && ~x18 )
						nx_state = s1;
					else if( x24 && ~x26 )
						nx_state = s1;
					else if( ~x24 && x25 && x26 && x18 )
						nx_state = s1;
					else if( ~x24 && x25 && x26 && ~x18 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x24 && x25 && ~x26 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x25 && ~x26 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x25 && ~x26 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x26 && ~x19 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 )
						nx_state = s1;
					else nx_state = s164;
				s165 : if( x24 && x26 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( x24 && x26 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( x24 && x26 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x24 && x26 && ~x18 )
						nx_state = s1;
					else if( x24 && ~x26 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x24 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x25 && x19 && ~x14 && ~x13 && x26 )
						nx_state = s165;
					else if( ~x24 && x25 && x19 && ~x14 && ~x13 && ~x26 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && x5 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x5 && x18 && x15 && x12 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x5 && x18 && x15 && ~x12 && x11 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x5 && x18 && x15 && ~x12 && ~x11 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x5 && x18 && x15 && ~x12 && ~x11 && ~x10 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x5 && x18 && ~x15 && x16 && x10 && x12 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s282;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x5 && x18 && ~x15 && x16 && x10 && ~x12 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s392;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x5 && x18 && ~x15 && x16 && ~x10 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s282;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x5 && x18 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x5 && ~x18 )
						begin
							y11 = 1'b1;	y16 = 1'b1;	y25 = 1'b1;	
							nx_state = s281;
						end
					else nx_state = s165;
				s166 : if( x24 && x26 && x11 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s160;
						end
					else if( x24 && x26 && ~x11 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( x24 && x26 && ~x11 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( x24 && x26 && ~x11 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x24 && x26 && ~x11 && ~x18 )
						nx_state = s1;
					else if( x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x24 && x26 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x26 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x26 && x25 && x19 && ~x14 && ~x13 )
						nx_state = s166;
					else if( ~x24 && x26 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x24 && x26 && ~x25 && x10 && x12 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x24 && x26 && ~x25 && x10 && x12 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x24 && x26 && ~x25 && x10 && x12 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && x26 && ~x25 && x10 && x12 && ~x18 )
						nx_state = s1;
					else if( ~x24 && x26 && ~x25 && x10 && ~x12 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s165;
						end
					else if( ~x24 && x26 && ~x25 && ~x10 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x24 && x26 && ~x25 && ~x10 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x24 && x26 && ~x25 && ~x10 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && x26 && ~x25 && ~x10 && ~x18 )
						nx_state = s1;
					else if( ~x24 && ~x26 && x10 && x12 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && ~x26 && x10 && x12 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && ~x26 && x10 && x12 && x25 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x26 && x10 && x12 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x24 && ~x26 && x10 && x12 && ~x25 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x24 && ~x26 && x10 && x12 && ~x25 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x24 && ~x26 && x10 && x12 && ~x25 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x26 && x10 && x12 && ~x25 && ~x17 )
						nx_state = s1;
					else if( ~x24 && ~x26 && x10 && ~x12 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x24 && ~x26 && ~x10 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && ~x26 && ~x10 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && ~x26 && ~x10 && x25 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x26 && ~x10 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x24 && ~x26 && ~x10 && ~x25 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x24 && ~x26 && ~x10 && ~x25 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x24 && ~x26 && ~x10 && ~x25 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x26 && ~x10 && ~x25 && ~x17 )
						nx_state = s1;
					else nx_state = s166;
				s167 : if( x24 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s282;
						end
					else if( ~x24 )
						begin
							y8 = 1'b1;	y17 = 1'b1;	y23 = 1'b1;	
							nx_state = s164;
						end
					else nx_state = s167;
				s168 : if( x66 && x42 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x66 && x42 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x66 && x42 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s151;
						end
					else if( x66 && x42 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y28 = 1'b1;	
							nx_state = s135;
						end
					else if( x66 && ~x42 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s400;
						end
					else if( ~x66 && x24 )
						nx_state = s1;
					else if( ~x66 && ~x24 && x25 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x66 && ~x24 && ~x25 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else nx_state = s168;
				s169 : if( x65 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x4 )
						nx_state = s1;
					else if( ~x65 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else nx_state = s169;
				s170 : if( 1'b1 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else nx_state = s170;
				s171 : if( x24 && x26 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( x24 && x26 && ~x4 && x20 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( x24 && x26 && ~x4 && ~x20 && x21 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( x24 && x26 && ~x4 && ~x20 && ~x21 && x22 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( x24 && x26 && ~x4 && ~x20 && ~x21 && ~x22 && x23 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( x24 && x26 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && x16 && x11 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s49;
						end
					else if( x24 && x26 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && x16 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x24 && x26 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && x13 && x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x24 && x26 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && x13 && ~x11 && x12 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( x24 && x26 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && x13 && ~x11 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x24 && x26 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && ~x13 && x11 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( x24 && x26 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && ~x13 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x24 && x26 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s51;
						end
					else if( x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x24 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x25 && x19 && ~x14 && ~x13 && x26 )
						nx_state = s171;
					else if( ~x24 && x25 && x19 && ~x14 && ~x13 && ~x26 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x24 && ~x25 && ~x26 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x24 && ~x25 && ~x26 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && ~x17 )
						nx_state = s1;
					else nx_state = s171;
				s172 : if( x67 && x24 && x26 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x67 && x24 && ~x26 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( x67 && ~x24 && x25 && x26 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x67 && ~x24 && x25 && ~x26 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( x67 && ~x24 && ~x25 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x67 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x67 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x67 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x67 && ~x3 )
						nx_state = s1;
					else nx_state = s172;
				s173 : if( x67 )
						begin
							y15 = 1'b1;	
							nx_state = s355;
						end
					else if( ~x67 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s105;
						end
					else nx_state = s173;
				s174 : if( x65 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x4 )
						nx_state = s1;
					else if( ~x65 && x24 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x65 && ~x24 && x15 && x10 && x11 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s187;
						end
					else if( ~x65 && ~x24 && x15 && x10 && ~x11 && x12 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x65 && ~x24 && x15 && x10 && ~x11 && ~x12 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x65 && ~x24 && x15 && ~x10 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && ~x24 && ~x15 && x16 && x10 && x12 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s282;
						end
					else if( ~x65 && ~x24 && ~x15 && x16 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && ~x24 && ~x15 && x16 && ~x10 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s282;
						end
					else if( ~x65 && ~x24 && ~x15 && ~x16 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else nx_state = s174;
				s175 : if( x24 && x26 )
						begin
							y11 = 1'b1;	y16 = 1'b1;	y25 = 1'b1;	
							nx_state = s281;
						end
					else if( x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x24 && x25 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else nx_state = s175;
				s176 : if( x21 && x9 && x3 )
						nx_state = s40;
					else if( x21 && x9 && ~x3 && x4 )
						nx_state = s40;
					else if( x21 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( x21 && ~x9 )
						nx_state = s1;
					else if( ~x21 && x22 && x10 && x19 && x15 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y17 = 1'b1;	
							nx_state = s177;
						end
					else if( ~x21 && x22 && x10 && x19 && ~x15 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && x15 && x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && x15 && ~x14 && x16 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && x15 && ~x14 && ~x16 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && x15 && ~x14 && ~x16 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && x15 && ~x14 && ~x16 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && x10 && ~x19 && x20 && x15 && ~x14 && ~x16 && ~x5 )
						nx_state = s1;
					else if( ~x21 && x22 && x10 && ~x19 && x20 && ~x15 && x14 && x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && ~x15 && x14 && ~x18 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && ~x15 && x14 && ~x18 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && ~x15 && x14 && ~x18 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && x10 && ~x19 && x20 && ~x15 && x14 && ~x18 && ~x5 )
						nx_state = s1;
					else if( ~x21 && x22 && x10 && ~x19 && x20 && ~x15 && ~x14 && x17 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							y6 = 1'b1;	
							nx_state = s178;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && x10 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && x10 && ~x19 && x20 && ~x15 && ~x14 && ~x17 && ~x5 )
						nx_state = s1;
					else if( ~x21 && x22 && x10 && ~x19 && ~x20 )
						begin
							y21 = 1'b1;	
							nx_state = s151;
						end
					else if( ~x21 && x22 && ~x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && x19 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x21 && ~x22 && x19 && ~x15 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x21 && ~x22 && ~x19 && x20 )
						begin
							y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s179;
						end
					else if( ~x21 && ~x22 && ~x19 && ~x20 )
						begin
							y21 = 1'b1;	
							nx_state = s151;
						end
					else nx_state = s176;
				s177 : if( x21 && x9 && x3 )
						nx_state = s40;
					else if( x21 && x9 && ~x3 && x4 )
						nx_state = s40;
					else if( x21 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( x21 && ~x9 )
						nx_state = s1;
					else if( ~x21 && x22 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x5 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x19 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x21 && ~x22 && x19 && ~x15 )
						begin
							y2 = 1'b1;	y18 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x21 && ~x22 && ~x19 )
						begin
							y21 = 1'b1;	
							nx_state = s151;
						end
					else nx_state = s177;
				s178 : if( x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x5 )
						nx_state = s1;
					else nx_state = s178;
				s179 : if( x21 && x6 )
						begin
							y8 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s106;
						end
					else if( x21 && ~x6 && x8 && x19 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( x21 && ~x6 && x8 && ~x19 && x20 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							y17 = 1'b1;	
							nx_state = s176;
						end
					else if( x21 && ~x6 && x8 && ~x19 && ~x20 )
						begin
							y17 = 1'b1;	y21 = 1'b1;	
							nx_state = s377;
						end
					else if( x21 && ~x6 && ~x8 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	
							nx_state = s378;
						end
					else if( ~x21 && x22 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s179;
				s180 : if( x21 && x16 && x15 && x10 && x12 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( x21 && x16 && x15 && x10 && ~x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( x21 && x16 && x15 && ~x10 && x11 && x12 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s339;
						end
					else if( x21 && x16 && x15 && ~x10 && x11 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s331;
						end
					else if( x21 && x16 && x15 && ~x10 && ~x11 && x12 && x13 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s335;
						end
					else if( x21 && x16 && x15 && ~x10 && ~x11 && x12 && ~x13 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x16 && x15 && ~x10 && ~x11 && x12 && ~x13 && x18 && ~x14 )
						nx_state = s1;
					else if( x21 && x16 && x15 && ~x10 && ~x11 && x12 && ~x13 && ~x18 )
						nx_state = s1;
					else if( x21 && x16 && x15 && ~x10 && ~x11 && ~x12 && x14 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s335;
						end
					else if( x21 && x16 && x15 && ~x10 && ~x11 && ~x12 && ~x14 && x18 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x16 && x15 && ~x10 && ~x11 && ~x12 && ~x14 && x18 && ~x13 )
						nx_state = s1;
					else if( x21 && x16 && x15 && ~x10 && ~x11 && ~x12 && ~x14 && ~x18 )
						nx_state = s1;
					else if( x21 && x16 && ~x15 && x12 && x10 && x8 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x16 && ~x15 && x12 && x10 && x8 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x16 && ~x15 && x12 && x10 && x8 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x16 && ~x15 && x12 && x10 && x8 && ~x18 )
						nx_state = s1;
					else if( x21 && x16 && ~x15 && x12 && x10 && ~x8 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( x21 && x16 && ~x15 && x12 && x10 && ~x8 && ~x3 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( x21 && x16 && ~x15 && x12 && x10 && ~x8 && ~x3 && ~x5 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( x21 && x16 && ~x15 && x12 && ~x10 && x7 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( x21 && x16 && ~x15 && x12 && ~x10 && x7 && ~x3 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( x21 && x16 && ~x15 && x12 && ~x10 && x7 && ~x3 && ~x5 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( x21 && x16 && ~x15 && x12 && ~x10 && ~x7 && x11 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( x21 && x16 && ~x15 && x12 && ~x10 && ~x7 && x11 && ~x3 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( x21 && x16 && ~x15 && x12 && ~x10 && ~x7 && x11 && ~x3 && ~x5 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( x21 && x16 && ~x15 && x12 && ~x10 && ~x7 && ~x11 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x16 && ~x15 && x12 && ~x10 && ~x7 && ~x11 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x16 && ~x15 && x12 && ~x10 && ~x7 && ~x11 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x16 && ~x15 && x12 && ~x10 && ~x7 && ~x11 && ~x18 )
						nx_state = s1;
					else if( x21 && x16 && ~x15 && ~x12 && x10 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( x21 && x16 && ~x15 && ~x12 && x10 && ~x3 && x5 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s315;
						end
					else if( x21 && x16 && ~x15 && ~x12 && x10 && ~x3 && ~x5 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s370;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && x11 && x9 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && x11 && x9 && ~x3 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && x11 && x9 && ~x3 && ~x5 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && ~x18 )
						nx_state = s1;
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && ~x11 && x8 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && ~x11 && x8 && ~x3 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && ~x11 && x8 && ~x3 && ~x5 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x16 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && ~x18 )
						nx_state = s1;
					else if( x21 && ~x16 && x15 && x10 && x11 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( x21 && ~x16 && x15 && x10 && ~x11 && x12 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s126;
						end
					else if( x21 && ~x16 && x15 && x10 && ~x11 && ~x12 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( x21 && ~x16 && x15 && x10 && ~x11 && ~x12 && ~x3 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( x21 && ~x16 && x15 && x10 && ~x11 && ~x12 && ~x3 && ~x5 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( x21 && ~x16 && x15 && ~x10 && x11 && x12 )
						begin
							y14 = 1'b1;	
							nx_state = s285;
						end
					else if( x21 && ~x16 && x15 && ~x10 && x11 && ~x12 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x21 && ~x16 && x15 && ~x10 && ~x11 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( x21 && ~x16 && x15 && ~x10 && ~x11 && ~x3 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( x21 && ~x16 && x15 && ~x10 && ~x11 && ~x3 && ~x5 && x12 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s333;
						end
					else if( x21 && ~x16 && x15 && ~x10 && ~x11 && ~x3 && ~x5 && ~x12 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s332;
						end
					else if( x21 && ~x16 && ~x15 && x3 )
						begin
							y1 = 1'b1;	
							nx_state = s163;
						end
					else if( x21 && ~x16 && ~x15 && ~x3 && x5 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( x21 && ~x16 && ~x15 && ~x3 && ~x5 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s5;
						end
					else if( ~x21 && x22 && x23 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x21 && x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x19 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 && x18 && x14 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x21 && ~x22 && ~x23 && x18 && ~x14 && x13 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x21 && ~x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 && ~x18 )
						nx_state = s1;
					else nx_state = s180;
				s181 : if( 1'b1 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else nx_state = s181;
				s182 : if( x68 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x68 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x68 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x68 && x20 && ~x18 )
						nx_state = s1;
					else if( x68 && ~x20 && x21 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( x68 && ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( x68 && ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( x68 && ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x68 && ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else if( ~x68 && x24 && x26 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x68 && x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x68 && x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x68 && x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x68 && x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x68 && ~x24 && x25 && x26 && x15 && x10 && x11 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x68 && ~x24 && x25 && x26 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s398;
						end
					else if( ~x68 && ~x24 && x25 && x26 && x15 && x10 && ~x11 && ~x12 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x68 && ~x24 && x25 && x26 && x15 && ~x10 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s399;
						end
					else if( ~x68 && ~x24 && x25 && x26 && ~x15 && x16 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s282;
						end
					else if( ~x68 && ~x24 && x25 && x26 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else if( ~x68 && ~x24 && x25 && ~x26 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && x19 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && x20 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && ~x20 && x21 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && ~x20 && ~x21 && x22 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && ~x20 && ~x21 && ~x22 && x16 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && ~x20 && ~x21 && ~x22 && x16 && ~x11 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && ~x20 && ~x21 && ~x22 && x16 && ~x11 && ~x12 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && ~x20 && ~x21 && ~x22 && x16 && ~x11 && ~x12 && ~x10 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && ~x20 && ~x21 && ~x22 && ~x16 && x17 && x10 && x12 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && ~x20 && ~x21 && ~x22 && ~x16 && x17 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && ~x20 && ~x21 && ~x22 && ~x16 && x17 && ~x10 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x68 && ~x24 && ~x25 && x26 && ~x19 && ~x20 && ~x21 && ~x22 && ~x16 && ~x17 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x68 && ~x24 && ~x25 && ~x26 && x15 && x12 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x68 && ~x24 && ~x25 && ~x26 && x15 && ~x12 && x11 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x68 && ~x24 && ~x25 && ~x26 && x15 && ~x12 && ~x11 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x68 && ~x24 && ~x25 && ~x26 && x15 && ~x12 && ~x11 && ~x10 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x68 && ~x24 && ~x25 && ~x26 && ~x15 && x16 && x10 && x12 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s282;
						end
					else if( ~x68 && ~x24 && ~x25 && ~x26 && ~x15 && x16 && x10 && ~x12 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s392;
						end
					else if( ~x68 && ~x24 && ~x25 && ~x26 && ~x15 && x16 && ~x10 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s282;
						end
					else if( ~x68 && ~x24 && ~x25 && ~x26 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else nx_state = s182;
				s183 : if( x24 && x4 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( x24 && ~x4 && x20 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( x24 && ~x4 && ~x20 && x21 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( x24 && ~x4 && ~x20 && ~x21 && x22 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( x24 && ~x4 && ~x20 && ~x21 && ~x22 && x23 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( x24 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && x16 && x11 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s49;
						end
					else if( x24 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && x16 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x24 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && x13 && x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x24 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && x13 && ~x11 && x12 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( x24 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && x13 && ~x11 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x24 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && ~x13 && x11 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( x24 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && x17 && ~x13 && ~x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( x24 && ~x4 && ~x20 && ~x21 && ~x22 && ~x23 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s51;
						end
					else if( ~x24 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x19 && ~x14 && ~x13 )
						nx_state = s183;
					else if( ~x24 && ~x19 )
						nx_state = s1;
					else nx_state = s183;
				s184 : if( 1'b1 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else nx_state = s184;
				s185 : if( x26 )
						begin
							y14 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x26 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else nx_state = s185;
				s186 : if( x68 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	y22 = 1'b1;	
							nx_state = s401;
						end
					else if( ~x68 && x26 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x68 && ~x26 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s46;
						end
					else nx_state = s186;
				s187 : if( 1'b1 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else nx_state = s187;
				s188 : if( x66 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 && x24 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x66 && ~x24 && x26 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x66 && ~x24 && ~x26 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else nx_state = s188;
				s189 : if( x65 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( ~x65 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s402;
						end
					else nx_state = s189;
				s190 : if( x66 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x66 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s167;
						end
					else nx_state = s190;
				s191 : if( x65 && x66 && x68 && x21 && x20 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s403;
						end
					else if( x65 && x66 && x68 && x21 && ~x20 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( x65 && x66 && x68 && ~x21 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( x65 && x66 && ~x68 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( x65 && ~x66 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x65 && x16 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x65 && ~x16 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else nx_state = s191;
				s192 : if( x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x19 )
						nx_state = s1;
					else nx_state = s192;
				s193 : if( x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( ~x21 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else nx_state = s193;
				s194 : if( x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x21 && ~x20 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x19 )
						nx_state = s1;
					else nx_state = s194;
				s195 : if( x21 && x20 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s194;
						end
					else if( x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x19 )
						nx_state = s1;
					else nx_state = s195;
				s196 : if( x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x21 && ~x20 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x21 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else nx_state = s196;
				s197 : if( x21 && x65 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x65 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x65 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x65 && x20 && ~x17 )
						nx_state = s1;
					else if( x21 && x65 && ~x20 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x21 && ~x65 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && ~x65 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && ~x65 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x65 && ~x18 )
						nx_state = s1;
					else if( ~x21 && x65 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x65 && x22 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x21 && ~x65 && x22 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x21 && ~x65 && x22 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x65 && x22 && x23 && ~x17 )
						nx_state = s1;
					else if( ~x21 && ~x65 && x22 && ~x23 && x18 && x14 )
						nx_state = s40;
					else if( ~x21 && ~x65 && x22 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s40;
					else if( ~x21 && ~x65 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x65 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x21 && ~x65 && ~x22 && x23 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s180;
						end
					else if( ~x21 && ~x65 && ~x22 && ~x23 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s404;
						end
					else nx_state = s197;
				s198 : if( x65 && x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x65 && x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x19 )
						nx_state = s1;
					else if( ~x65 && x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x20 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x65 && ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x65 && ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else nx_state = s198;
				s199 : if( x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x21 && ~x20 && x10 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s302;
						end
					else if( x21 && ~x20 && ~x10 && x11 && x12 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x20 && ~x10 && x11 && x12 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x20 && ~x10 && x11 && x12 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x20 && ~x10 && x11 && x12 && ~x19 )
						nx_state = s1;
					else if( x21 && ~x20 && ~x10 && x11 && ~x12 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s302;
						end
					else if( x21 && ~x20 && ~x10 && ~x11 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x21 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x21 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x21 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x19 )
						nx_state = s1;
					else nx_state = s199;
				s200 : if( 1'b1 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s405;
						end
					else nx_state = s200;
				s201 : if( x20 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x20 && x21 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( ~x20 && ~x21 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else nx_state = s201;
				s202 : if( x10 && x12 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s259;
						end
					else if( x10 && ~x12 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x10 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s259;
						end
					else nx_state = s202;
				s203 : if( x65 && x21 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x65 && x21 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x65 && x21 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x65 && x21 && ~x8 )
						nx_state = s1;
					else if( x65 && ~x21 && x23 && x22 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && x23 && x22 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && x23 && x22 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && ~x21 && x23 && x22 && ~x8 )
						nx_state = s1;
					else if( x65 && ~x21 && x23 && ~x22 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && x23 && ~x22 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && x23 && ~x22 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && ~x21 && x23 && ~x22 && ~x9 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x23 && x8 && x22 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && ~x23 && x8 && x22 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && ~x23 && x8 && x22 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x23 && x8 && ~x22 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && ~x23 && x8 && ~x22 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x21 && ~x23 && x8 && ~x22 && ~x10 && ~x11 )
						nx_state = s1;
					else if( x65 && ~x21 && ~x23 && ~x8 )
						nx_state = s1;
					else if( ~x65 && x66 && x62 && x61 && x13 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && x66 && x62 && x61 && ~x13 && x12 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && x66 && x62 && x61 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x66 && x62 && ~x61 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x62 && x63 && x17 && x13 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && x66 && ~x62 && x63 && x17 && x13 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && x66 && ~x62 && x63 && x17 && ~x13 && x12 && x64 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x65 && x66 && ~x62 && x63 && x17 && ~x13 && x12 && ~x64 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && x66 && ~x62 && x63 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x62 && x63 && ~x17 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x62 && ~x63 && x19 && x13 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && x19 && x13 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && x19 && ~x13 && x12 && x64 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && x19 && ~x13 && x12 && ~x64 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x66 && ~x62 && ~x63 && x19 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x62 && ~x63 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x21 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x65 && ~x66 && ~x21 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else nx_state = s203;
				s204 : if( 1'b1 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else nx_state = s204;
				s205 : if( x21 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && x22 && x23 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && x22 && ~x23 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x21 && ~x22 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s147;
						end
					else nx_state = s205;
				s206 : if( x20 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x20 && ~x15 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else nx_state = s206;
				s207 : if( x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x20 && ~x18 )
						nx_state = s1;
					else if( ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else nx_state = s207;
				s208 : if( x1 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	
							nx_state = s277;
						end
					else if( ~x1 && x17 && x15 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x1 && x17 && ~x15 && x16 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s59;
						end
					else if( ~x1 && x17 && ~x15 && ~x16 )
						begin
							y7 = 1'b1;	y12 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x1 && ~x17 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	y22 = 1'b1;	
							nx_state = s401;
						end
					else nx_state = s208;
				s209 : if( x20 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s393;
						end
					else if( ~x20 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else nx_state = s209;
				s210 : if( x65 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x65 && x66 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x66 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x66 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x65 && x66 && ~x4 )
						nx_state = s1;
					else if( ~x65 && ~x66 && x20 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s393;
						end
					else if( ~x65 && ~x66 && ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x66 && ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x66 && ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x20 && ~x21 && x17 && x13 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x65 && ~x66 && ~x20 && ~x21 && x17 && ~x13 && x12 )
						begin
							y1 = 1'b1;	y10 = 1'b1;	
							nx_state = s148;
						end
					else if( ~x65 && ~x66 && ~x20 && ~x21 && x17 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x66 && ~x20 && ~x21 && ~x17 )
						nx_state = s1;
					else nx_state = s210;
				s211 : if( x66 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x66 && x21 && ~x19 )
						nx_state = s1;
					else if( x66 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x66 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x66 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x66 && ~x21 && ~x20 )
						nx_state = s1;
					else if( ~x66 && x20 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s393;
						end
					else if( ~x66 && ~x20 && x21 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x66 && ~x20 && x21 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x66 && ~x20 && x21 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x66 && ~x20 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x66 && ~x20 && ~x21 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else nx_state = s211;
				s212 : if( x21 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && x22 && x23 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && x22 && ~x23 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x21 && ~x22 && x23 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s147;
						end
					else if( ~x21 && ~x22 && ~x23 && x18 && x14 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && ~x22 && ~x23 && x18 && ~x14 && x13 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( ~x21 && ~x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 && ~x18 )
						nx_state = s1;
					else nx_state = s212;
				s213 : if( x64 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( ~x64 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s152;
						end
					else nx_state = s213;
				s214 : if( x21 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x21 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s308;
						end
					else nx_state = s214;
				s215 : if( 1'b1 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else nx_state = s215;
				s216 : if( x21 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x21 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x21 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x21 && ~x9 )
						nx_state = s1;
					else if( ~x21 && x22 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && ~x22 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s216;
				s217 : if( x21 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x21 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x21 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x21 && ~x9 )
						nx_state = s1;
					else if( ~x21 && x22 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x21 && x22 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x21 && x22 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x7 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s217;
				s218 : if( x21 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x21 && x22 && x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s219;
						end
					else if( ~x21 && x22 && ~x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s28;
						end
					else if( ~x21 && ~x22 && x8 && x16 && x15 && x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s219;
						end
					else if( ~x21 && ~x22 && x8 && x16 && x15 && ~x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s309;
						end
					else if( ~x21 && ~x22 && x8 && x16 && ~x15 && x10 )
						begin
							y2 = 1'b1;	y16 = 1'b1;	y24 = 1'b1;	
							nx_state = s124;
						end
					else if( ~x21 && ~x22 && x8 && x16 && ~x15 && ~x10 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s310;
						end
					else if( ~x21 && ~x22 && x8 && ~x16 && x17 && x10 && x15 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s219;
						end
					else if( ~x21 && ~x22 && x8 && ~x16 && x17 && x10 && ~x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s308;
						end
					else if( ~x21 && ~x22 && x8 && ~x16 && x17 && ~x10 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s79;
						end
					else if( ~x21 && ~x22 && x8 && ~x16 && ~x17 && x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s219;
						end
					else if( ~x21 && ~x22 && x8 && ~x16 && ~x17 && ~x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s311;
						end
					else if( ~x21 && ~x22 && ~x8 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else nx_state = s218;
				s219 : if( 1'b1 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else nx_state = s219;
				s220 : if( x21 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s311;
						end
					else if( ~x21 && x22 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && ~x22 && x3 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s218;
						end
					else if( ~x21 && ~x22 && ~x3 && x8 && x16 && x15 && x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s219;
						end
					else if( ~x21 && ~x22 && ~x3 && x8 && x16 && x15 && ~x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s309;
						end
					else if( ~x21 && ~x22 && ~x3 && x8 && x16 && ~x15 && x10 )
						begin
							y2 = 1'b1;	y16 = 1'b1;	y24 = 1'b1;	
							nx_state = s124;
						end
					else if( ~x21 && ~x22 && ~x3 && x8 && x16 && ~x15 && ~x10 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s310;
						end
					else if( ~x21 && ~x22 && ~x3 && x8 && ~x16 && x17 && x10 && x15 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s219;
						end
					else if( ~x21 && ~x22 && ~x3 && x8 && ~x16 && x17 && x10 && ~x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s308;
						end
					else if( ~x21 && ~x22 && ~x3 && x8 && ~x16 && x17 && ~x10 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s79;
						end
					else if( ~x21 && ~x22 && ~x3 && x8 && ~x16 && ~x17 && x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s219;
						end
					else if( ~x21 && ~x22 && ~x3 && x8 && ~x16 && ~x17 && ~x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s311;
						end
					else if( ~x21 && ~x22 && ~x3 && ~x8 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else nx_state = s220;
				s221 : if( x21 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x21 && x22 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && ~x22 )
						begin
							y2 = 1'b1;	y16 = 1'b1;	y24 = 1'b1;	
							nx_state = s124;
						end
					else nx_state = s221;
				s222 : if( 1'b1 )
						begin
							y17 = 1'b1;	
							nx_state = s17;
						end
					else nx_state = s222;
				s223 : if( x21 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s161;
						end
					else if( ~x21 && x22 && x8 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x8 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x12 && x23 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x21 && ~x22 && x12 && ~x23 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x21 && ~x22 && ~x12 && x23 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && ~x12 && x23 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && ~x12 && x23 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x12 && x23 && ~x9 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x12 && ~x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && ~x12 && ~x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && ~x12 && ~x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x12 && ~x23 && ~x8 )
						nx_state = s1;
					else nx_state = s223;
				s224 : if( x66 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( ~x66 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else nx_state = s224;
				s225 : if( 1'b1 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s123;
						end
					else nx_state = s225;
				s226 : if( x21 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && x22 && x17 && x10 && x15 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x21 && x22 && x17 && x10 && ~x15 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x21 && x22 && x17 && ~x10 )
						begin
							y13 = 1'b1;	y16 = 1'b1;	
							nx_state = s284;
						end
					else if( ~x21 && x22 && ~x17 && x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s219;
						end
					else if( ~x21 && x22 && ~x17 && ~x10 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	
							nx_state = s217;
						end
					else if( ~x21 && ~x22 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s226;
				s227 : if( x21 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x23 && x22 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x23 && x22 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x23 && x22 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x23 && x22 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x23 && ~x22 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x23 && ~x22 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x23 && ~x22 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x23 && ~x22 && ~x9 )
						nx_state = s1;
					else if( ~x21 && ~x23 && x8 && x22 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x23 && x8 && x22 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x23 && x8 && x22 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && ~x23 && x8 && ~x22 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x23 && x8 && ~x22 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x23 && x8 && ~x22 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x23 && ~x8 )
						nx_state = s1;
					else nx_state = s227;
				s228 : if( x21 && x18 )
						begin
							y14 = 1'b1;	y19 = 1'b1;	
							nx_state = s116;
						end
					else if( x21 && ~x18 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s117;
						end
					else if( ~x21 && x22 && x23 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x21 && x22 && x23 && ~x12 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x23 && ~x12 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x23 && ~x12 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x12 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s243;
						end
					else if( ~x21 && ~x22 )
						begin
							y14 = 1'b1;	y19 = 1'b1;	
							nx_state = s116;
						end
					else nx_state = s228;
				s229 : if( x21 && x18 && x4 && x15 && x17 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x21 && x18 && x4 && x15 && ~x17 )
						begin
							y12 = 1'b1;	
							nx_state = s231;
						end
					else if( x21 && x18 && x4 && ~x15 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s235;
						end
					else if( x21 && x18 && ~x4 )
						begin
							y12 = 1'b1;	
							nx_state = s231;
						end
					else if( x21 && ~x18 && x19 && x15 && x4 && x17 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x21 && ~x18 && x19 && x15 && x4 && ~x17 )
						begin
							y12 = 1'b1;	
							nx_state = s231;
						end
					else if( x21 && ~x18 && x19 && x15 && ~x4 )
						begin
							y12 = 1'b1;	
							nx_state = s231;
						end
					else if( x21 && ~x18 && x19 && ~x15 && x16 && x14 )
						begin
							y12 = 1'b1;	
							nx_state = s231;
						end
					else if( x21 && ~x18 && x19 && ~x15 && x16 && ~x14 && x17 )
						begin
							y12 = 1'b1;	
							nx_state = s231;
						end
					else if( x21 && ~x18 && x19 && ~x15 && x16 && ~x14 && ~x17 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && ~x18 && x19 && ~x15 && x16 && ~x14 && ~x17 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && ~x18 && x19 && ~x15 && x16 && ~x14 && ~x17 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x18 && x19 && ~x15 && x16 && ~x14 && ~x17 && ~x8 )
						nx_state = s1;
					else if( x21 && ~x18 && x19 && ~x15 && ~x16 && x17 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s231;
						end
					else if( x21 && ~x18 && x19 && ~x15 && ~x16 && x17 && ~x12 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && ~x18 && x19 && ~x15 && ~x16 && x17 && ~x12 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && ~x18 && x19 && ~x15 && ~x16 && x17 && ~x12 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x18 && x19 && ~x15 && ~x16 && x17 && ~x12 && ~x8 )
						nx_state = s1;
					else if( x21 && ~x18 && x19 && ~x15 && ~x16 && ~x17 && x13 )
						begin
							y12 = 1'b1;	
							nx_state = s231;
						end
					else if( x21 && ~x18 && x19 && ~x15 && ~x16 && ~x17 && ~x13 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && ~x18 && x19 && ~x15 && ~x16 && ~x17 && ~x13 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && ~x18 && x19 && ~x15 && ~x16 && ~x17 && ~x13 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x18 && x19 && ~x15 && ~x16 && ~x17 && ~x13 && ~x8 )
						nx_state = s1;
					else if( x21 && ~x18 && ~x19 && x4 )
						begin
							y15 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s36;
						end
					else if( x21 && ~x18 && ~x19 && ~x4 )
						begin
							y12 = 1'b1;	
							nx_state = s231;
						end
					else if( ~x21 && x23 && x22 && x6 )
						begin
							y12 = 1'b1;	
							nx_state = s231;
						end
					else if( ~x21 && x23 && x22 && ~x6 && x7 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( ~x21 && x23 && x22 && ~x6 && x7 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x21 && x23 && x22 && ~x6 && x7 && ~x18 && x19 && x15 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x21 && x23 && x22 && ~x6 && x7 && ~x18 && x19 && ~x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( ~x21 && x23 && x22 && ~x6 && x7 && ~x18 && ~x19 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s33;
						end
					else if( ~x21 && x23 && x22 && ~x6 && ~x7 )
						begin
							y3 = 1'b1;	y12 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x21 && x23 && ~x22 )
						begin
							y12 = 1'b1;	y19 = 1'b1;	
							nx_state = s230;
						end
					else if( ~x21 && ~x23 && x22 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s161;
						end
					else if( ~x21 && ~x23 && ~x22 && x6 )
						begin
							y12 = 1'b1;	
							nx_state = s231;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x6 && x7 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x6 && x7 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x6 && x7 && ~x18 && x19 && x15 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x6 && x7 && ~x18 && x19 && ~x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x6 && x7 && ~x18 && ~x19 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s33;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x6 && ~x7 )
						begin
							y3 = 1'b1;	y12 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s34;
						end
					else nx_state = s229;
				s230 : if( x21 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( ~x21 && x22 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x21 && x22 && ~x18 && x19 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x21 && x22 && ~x18 && x19 && ~x15 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x21 && x22 && ~x18 && ~x19 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x16 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x16 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && x16 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s228;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && ~x20 )
						begin
							y12 = 1'b1;	
							nx_state = s231;
						end
					else if( ~x21 && ~x22 && ~x23 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( ~x21 && ~x22 && ~x23 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x21 && ~x22 && ~x23 && ~x18 && x19 && x15 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( ~x21 && ~x22 && ~x23 && ~x18 && ~x19 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s33;
						end
					else nx_state = s230;
				s231 : if( x65 && x66 )
						nx_state = s40;
					else if( x65 && ~x66 && x21 && x5 )
						begin
							y3 = 1'b1;	y12 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s34;
						end
					else if( x65 && ~x66 && x21 && ~x5 && x6 && x18 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && ~x66 && x21 && ~x5 && x6 && x18 && x15 && ~x17 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	
							nx_state = s244;
						end
					else if( x65 && ~x66 && x21 && ~x5 && x6 && x18 && ~x15 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x65 && ~x66 && x21 && ~x5 && x6 && ~x18 && x19 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && ~x66 && x21 && ~x5 && x6 && ~x18 && x19 && x15 && ~x17 )
						begin
							y8 = 1'b1;	
							nx_state = s246;
						end
					else if( x65 && ~x66 && x21 && ~x5 && x6 && ~x18 && x19 && ~x15 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s227;
						end
					else if( x65 && ~x66 && x21 && ~x5 && x6 && ~x18 && ~x19 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s31;
						end
					else if( x65 && ~x66 && x21 && ~x5 && ~x6 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s247;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x23 && x7 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x23 && x7 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x23 && x7 && ~x18 && x19 && x15 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s247;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x23 && x7 && ~x18 && x19 && ~x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x23 && x7 && ~x18 && ~x19 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s33;
						end
					else if( x65 && ~x66 && ~x21 && x22 && x23 && ~x7 )
						begin
							y3 = 1'b1;	y12 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s34;
						end
					else if( x65 && ~x66 && ~x21 && x22 && ~x23 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s161;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && x23 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s161;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x23 && x7 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x23 && x7 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x23 && x7 && ~x18 && x19 && x15 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s247;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x23 && x7 && ~x18 && x19 && ~x15 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x23 && x7 && ~x18 && ~x19 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s33;
						end
					else if( x65 && ~x66 && ~x21 && ~x22 && ~x23 && ~x7 )
						begin
							y3 = 1'b1;	y12 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s34;
						end
					else if( ~x65 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else nx_state = s231;
				s232 : if( x21 )
						nx_state = s1;
					else if( ~x21 && x22 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x21 && ~x22 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s322;
						end
					else nx_state = s232;
				s233 : if( x21 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s161;
						end
					else if( ~x21 && ~x22 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s161;
						end
					else nx_state = s233;
				s234 : if( x21 && x65 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && x65 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && x65 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && x65 && ~x8 )
						nx_state = s1;
					else if( x21 && ~x65 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x21 && x65 && x23 && x22 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x65 && x23 && x22 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x65 && x23 && x22 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x65 && x23 && x22 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x65 && x23 && ~x22 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x65 && x23 && ~x22 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x65 && x23 && ~x22 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x65 && x23 && ~x22 && ~x9 )
						nx_state = s1;
					else if( ~x21 && x65 && ~x23 && x8 && x22 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x65 && ~x23 && x8 && x22 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x65 && ~x23 && x8 && x22 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && x65 && ~x23 && x8 && ~x22 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x65 && ~x23 && x8 && ~x22 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x65 && ~x23 && x8 && ~x22 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x65 && ~x23 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x65 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else nx_state = s234;
				s235 : if( x21 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s161;
						end
					else if( ~x21 && ~x22 && x23 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s161;
						end
					else if( ~x21 && ~x22 && ~x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && ~x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && ~x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 && ~x8 )
						nx_state = s1;
					else nx_state = s235;
				s236 : if( 1'b1 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s28;
						end
					else nx_state = s236;
				s237 : if( x21 && x18 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && x18 && x15 && ~x17 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	
							nx_state = s244;
						end
					else if( x21 && x18 && ~x15 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x21 && ~x18 && x19 && x15 && x17 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x18 && x19 && x15 && ~x17 )
						begin
							y8 = 1'b1;	
							nx_state = s246;
						end
					else if( x21 && ~x18 && x19 && ~x15 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s157;
						end
					else if( x21 && ~x18 && ~x19 )
						begin
							y1 = 1'b1;	y3 = 1'b1;	y4 = 1'b1;	
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s31;
						end
					else if( ~x21 && x22 && x23 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( ~x21 && x22 && x23 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x21 && x22 && x23 && ~x18 && x19 && x15 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x21 && x22 && x23 && ~x18 && x19 && ~x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x21 && x22 && x23 && ~x18 && ~x19 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s33;
						end
					else if( ~x21 && x22 && ~x23 )
						begin
							y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s161;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x16 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x16 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && x16 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s228;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && x18 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x18 && x17 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x18 && ~x17 && x5 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s283;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x18 && ~x17 && ~x5 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && ~x20 )
						begin
							y12 = 1'b1;	
							nx_state = s231;
						end
					else if( ~x21 && ~x22 && ~x23 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( ~x21 && ~x22 && ~x23 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x21 && ~x22 && ~x23 && ~x18 && x19 && x15 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x21 && ~x22 && ~x23 && ~x18 && x19 && ~x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x21 && ~x22 && ~x23 && ~x18 && ~x19 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s33;
						end
					else nx_state = s237;
				s238 : if( x21 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s33;
						end
					else if( ~x21 && x22 && x23 && x15 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s240;
						end
					else if( ~x21 && x22 && x23 && ~x15 && x19 && x18 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s240;
						end
					else if( ~x21 && x22 && x23 && ~x15 && x19 && ~x18 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x23 && ~x15 && x19 && ~x18 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x23 && ~x15 && x19 && ~x18 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x15 && x19 && ~x18 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x15 && ~x19 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s240;
						end
					else if( ~x21 && x22 && ~x23 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 && x15 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s240;
						end
					else if( ~x21 && ~x22 && ~x23 && ~x15 && x19 && x18 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s240;
						end
					else if( ~x21 && ~x22 && ~x23 && ~x15 && x19 && ~x18 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && ~x23 && ~x15 && x19 && ~x18 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && ~x23 && ~x15 && x19 && ~x18 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 && ~x15 && x19 && ~x18 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 && ~x15 && ~x19 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s240;
						end
					else nx_state = s238;
				s239 : if( x26 )
						begin
							y6 = 1'b1;	y13 = 1'b1;	
							nx_state = s165;
						end
					else if( ~x26 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s25;
						end
					else nx_state = s239;
				s240 : if( x21 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x21 && x22 && x23 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && x6 && x18 && x15 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( ~x21 && x22 && ~x23 && x6 && x18 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x21 && x22 && ~x23 && x6 && ~x18 && x19 && x15 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x21 && x22 && ~x23 && x6 && ~x18 && x19 && ~x15 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x21 && x22 && ~x23 && x6 && ~x18 && ~x19 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s229;
						end
					else if( ~x21 && x22 && ~x23 && ~x6 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s28;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x20 && x16 && x18 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x20 && x16 && ~x18 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x20 && ~x16 && x17 && x18 )
						begin
							y24 = 1'b1;	y25 = 1'b1;	
							nx_state = s157;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x20 && ~x16 && x17 && ~x18 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	y20 = 1'b1;	
							y26 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x20 && ~x16 && ~x17 && x18 && x11 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x20 && ~x16 && ~x17 && x18 && ~x11 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x20 && ~x16 && ~x17 && x18 && ~x11 && x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && x19 && x20 && ~x16 && ~x17 && x18 && ~x11 && ~x9 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && x19 && x20 && ~x16 && ~x17 && ~x18 && x10 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x20 && ~x16 && ~x17 && ~x18 && ~x10 && x9 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x20 && ~x16 && ~x17 && ~x18 && ~x10 && x9 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && x19 && x20 && ~x16 && ~x17 && ~x18 && ~x10 && ~x9 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && x19 && ~x20 && x17 && x16 )
						begin
							y18 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x20 && x17 && ~x16 && x18 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x20 && x17 && ~x16 && ~x18 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s233;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x20 && ~x17 && x18 && x16 )
						begin
							y18 = 1'b1;	
							nx_state = s234;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x20 && ~x17 && x18 && ~x16 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	y20 = 1'b1;	
							nx_state = s235;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x20 && ~x17 && ~x18 && x3 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x20 && ~x17 && ~x18 && ~x3 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x20 && ~x17 && ~x18 && ~x3 && ~x5 && x16 )
						begin
							y5 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x20 && ~x17 && ~x18 && ~x3 && ~x5 && ~x16 )
						begin
							y16 = 1'b1;	y20 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && x16 && x3 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && x16 && ~x3 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && x16 && ~x3 && ~x5 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && x17 && x18 && x3 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && x17 && x18 && ~x3 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && x17 && x18 && ~x3 && ~x5 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && x17 && ~x18 && x15 && x3 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && x17 && ~x18 && x15 && ~x3 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && x17 && ~x18 && x15 && ~x3 && ~x5 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && x17 && ~x18 && ~x15 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x17 && x18 && x13 && x3 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x17 && x18 && x13 && ~x3 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x17 && x18 && x13 && ~x3 && ~x5 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s227;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x17 && x18 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x17 && ~x18 && x12 && x3 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x17 && ~x18 && x12 && ~x3 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x17 && ~x18 && ~x12 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x17 && ~x18 && ~x12 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x17 && ~x18 && ~x12 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x19 && x20 && ~x16 && ~x17 && ~x18 && ~x12 && ~x9 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x19 && ~x20 && x3 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && ~x20 && ~x3 && x5 )
						begin
							y12 = 1'b1;	y16 = 1'b1;	
							nx_state = s237;
						end
					else if( ~x21 && ~x22 && x23 && ~x19 && ~x20 && ~x3 && ~x5 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( ~x21 && ~x22 && ~x23 )
						nx_state = s1;
					else nx_state = s240;
				s241 : if( 1'b1 )
						begin
							y7 = 1'b1;	
							nx_state = s338;
						end
					else nx_state = s241;
				s242 : if( x65 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( ~x65 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s51;
						end
					else nx_state = s242;
				s243 : if( x21 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x21 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x21 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	y21 = 1'b1;	
							nx_state = s117;
						end
					else if( ~x21 && x22 && ~x12 && x8 && x9 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && ~x12 && x8 && ~x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && ~x12 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x12 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x12 && x23 )
						begin
							y6 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s247;
						end
					else if( ~x21 && ~x22 && x12 && ~x23 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x21 && ~x22 && ~x12 && x23 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && ~x12 && x23 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && ~x12 && x23 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x12 && x23 && ~x9 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x12 && ~x23 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && ~x12 && ~x23 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && ~x12 && ~x23 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x12 && ~x23 && ~x8 )
						nx_state = s1;
					else nx_state = s243;
				s244 : if( x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x8 )
						nx_state = s1;
					else nx_state = s244;
				s245 : if( 1'b1 )
						begin
							y3 = 1'b1;	y12 = 1'b1;	y16 = 1'b1;	
							y17 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s406;
						end
					else nx_state = s245;
				s246 : if( x65 && x67 )
						begin
							y8 = 1'b1;	y16 = 1'b1;	
							nx_state = s407;
						end
					else if( x65 && ~x67 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x65 && x21 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x65 && x21 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x65 && x21 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x65 && x21 && ~x3 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 )
						nx_state = s1;
					else if( ~x65 && ~x21 && ~x22 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && ~x21 && ~x22 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && ~x21 && ~x22 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x65 && ~x21 && ~x22 && ~x8 )
						nx_state = s1;
					else nx_state = s246;
				s247 : if( x21 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	y8 = 1'b1;	
							nx_state = s238;
						end
					else if( ~x21 && x22 && x23 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x21 && x22 && x23 && ~x12 && x8 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x23 && ~x12 && x8 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && x22 && x23 && ~x12 && x8 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x12 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 )
						begin
							y14 = 1'b1;	y19 = 1'b1;	
							nx_state = s116;
						end
					else if( ~x21 && ~x22 && x23 && x9 && x10 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && x23 && x9 && ~x10 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x22 && x23 && x9 && ~x10 && ~x11 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x9 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 )
						begin
							y6 = 1'b1;	y19 = 1'b1;	
							nx_state = s223;
						end
					else nx_state = s247;
				s248 : if( x22 && x21 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( x22 && ~x21 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s409;
						end
					else if( ~x22 && x19 && x21 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( ~x22 && x19 && ~x21 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s409;
						end
					else if( ~x22 && ~x19 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else nx_state = s248;
				s249 : if( x21 && x18 && x16 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( x21 && x18 && ~x16 && x13 && x15 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( x21 && x18 && ~x16 && x13 && ~x15 && x17 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s409;
						end
					else if( x21 && x18 && ~x16 && x13 && ~x15 && ~x17 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( x21 && x18 && ~x16 && ~x13 && x17 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s409;
						end
					else if( x21 && x18 && ~x16 && ~x13 && ~x17 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( x21 && ~x18 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s409;
						end
					else if( ~x21 && x19 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( ~x21 && ~x19 && x22 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( ~x21 && ~x19 && ~x22 && x20 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s409;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x20 && x16 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && x15 && x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && x15 && ~x13 && x17 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s409;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && x15 && ~x13 && ~x17 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && ~x15 && x17 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s409;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && ~x15 && ~x17 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else nx_state = s249;
				s250 : if( x65 && x60 && x61 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s68;
						end
					else if( x65 && x60 && ~x61 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( x65 && ~x60 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x65 && x23 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s410;
						end
					else if( ~x65 && ~x23 && x19 )
						begin
							y14 = 1'b1;	
							nx_state = s285;
						end
					else if( ~x65 && ~x23 && ~x19 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s84;
						end
					else nx_state = s250;
				s251 : if( x60 && x61 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s256;
						end
					else if( x60 && ~x61 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x60 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else nx_state = s251;
				s252 : if( x60 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x60 && ~x7 && x61 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x60 && ~x7 && x61 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x60 && ~x7 && x61 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x60 && ~x7 && x61 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x60 && ~x7 && ~x61 )
						nx_state = s39;
					else if( ~x60 && x61 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x60 && x61 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x60 && x61 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( ~x60 && x61 && x62 && ~x18 )
						nx_state = s1;
					else if( ~x60 && x61 && ~x62 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( ~x60 && x61 && ~x62 && ~x7 )
						nx_state = s39;
					else if( ~x60 && ~x61 && x62 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x60 && ~x61 && ~x62 )
						nx_state = s40;
					else nx_state = s252;
				s253 : if( x60 && x61 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s257;
						end
					else if( x60 && ~x61 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x60 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else nx_state = s253;
				s254 : if( x65 && x60 && x61 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x60 && x61 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x60 && x61 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x60 && x61 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x60 && ~x61 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x60 && ~x61 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x60 && ~x61 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x65 && x60 && ~x61 && ~x18 )
						nx_state = s39;
					else if( x65 && ~x60 && x61 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && ~x60 && x61 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && ~x60 && x61 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x65 && ~x60 && x61 && x62 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x60 && x61 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x60 && x61 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x60 && x61 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x65 && ~x60 && x61 && ~x62 && ~x18 )
						nx_state = s39;
					else if( x65 && ~x60 && ~x61 )
						nx_state = s40;
					else if( ~x65 && x20 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && ~x20 && x18 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x20 && x18 && ~x13 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x65 && ~x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( ~x65 && ~x20 && ~x18 )
						nx_state = s1;
					else nx_state = s254;
				s255 : if( x67 && x22 && x4 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x67 && x22 && ~x4 && x20 && x15 && x8 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x67 && x22 && ~x4 && x20 && x15 && ~x8 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x67 && x22 && ~x4 && x20 && ~x15 && x16 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s302;
						end
					else if( x67 && x22 && ~x4 && x20 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s122;
						end
					else if( x67 && x22 && ~x4 && ~x20 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							y25 = 1'b1;	
							nx_state = s368;
						end
					else if( x67 && ~x22 && x23 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x67 && ~x22 && ~x23 )
						nx_state = s1;
					else if( ~x67 && x61 && x60 && x3 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s118;
						end
					else if( ~x67 && x61 && x60 && ~x3 && x18 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s38;
						end
					else if( ~x67 && x61 && x60 && ~x3 && ~x18 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s319;
						end
					else if( ~x67 && x61 && ~x60 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x67 && x61 && ~x60 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x67 && x61 && ~x60 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( ~x67 && x61 && ~x60 && x62 && ~x18 )
						nx_state = s1;
					else if( ~x67 && x61 && ~x60 && ~x62 && x19 && x15 )
						nx_state = s73;
					else if( ~x67 && x61 && ~x60 && ~x62 && x19 && ~x15 && x16 )
						begin
							y12 = 1'b1;	
							nx_state = s291;
						end
					else if( ~x67 && x61 && ~x60 && ~x62 && x19 && ~x15 && ~x16 )
						nx_state = s73;
					else if( ~x67 && x61 && ~x60 && ~x62 && ~x19 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y24 = 1'b1;	
							nx_state = s64;
						end
					else if( ~x67 && ~x61 && x60 && x19 && x15 )
						nx_state = s73;
					else if( ~x67 && ~x61 && x60 && x19 && ~x15 && x16 )
						begin
							y12 = 1'b1;	
							nx_state = s291;
						end
					else if( ~x67 && ~x61 && x60 && x19 && ~x15 && ~x16 )
						nx_state = s73;
					else if( ~x67 && ~x61 && x60 && ~x19 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y24 = 1'b1;	
							nx_state = s64;
						end
					else if( ~x67 && ~x61 && ~x60 && x62 )
						nx_state = s1;
					else if( ~x67 && ~x61 && ~x60 && ~x62 && x18 && x15 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x67 && ~x61 && ~x60 && ~x62 && x18 && x15 && ~x7 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x67 && ~x61 && ~x60 && ~x62 && x18 && x15 && ~x7 && ~x11 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && x4 )
						nx_state = s40;
					else if( ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && ~x4 && x11 && x9 )
						nx_state = s40;
					else if( ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && ~x4 && x11 && ~x9 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && ~x4 && x11 && ~x9 && ~x7 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s118;
						end
					else if( ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && ~x4 && ~x11 && x9 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && ~x4 && ~x11 && x9 && ~x7 && x10 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && ~x4 && ~x11 && x9 && ~x7 && ~x10 )
						nx_state = s40;
					else if( ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && x7 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && x7 && ~x8 )
						nx_state = s40;
					else if( ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && ~x7 && x12 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && ~x7 && ~x12 )
						nx_state = s40;
					else if( ~x67 && ~x61 && ~x60 && ~x62 && x18 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x67 && ~x61 && ~x60 && ~x62 && ~x18 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y24 = 1'b1;	
							nx_state = s64;
						end
					else nx_state = s255;
				s256 : if( x60 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s68;
						end
					else if( ~x60 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else nx_state = s256;
				s257 : if( 1'b1 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s68;
						end
					else nx_state = s257;
				s258 : if( x60 && x61 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( x60 && ~x61 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x60 && ~x61 && ~x2 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x60 && x61 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x60 && x61 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x60 && x61 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( ~x60 && x61 && x62 && ~x18 )
						nx_state = s1;
					else if( ~x60 && x61 && ~x62 && x2 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x60 && x61 && ~x62 && ~x2 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x60 && ~x61 && x62 && x7 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x60 && ~x61 && x62 && ~x7 )
						nx_state = s40;
					else if( ~x60 && ~x61 && ~x62 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else nx_state = s258;
				s259 : if( x21 && x20 && x10 && x12 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x20 && x10 && x12 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x20 && x10 && x12 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x20 && x10 && x12 && ~x17 )
						nx_state = s1;
					else if( x21 && x20 && x10 && ~x12 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s302;
						end
					else if( x21 && x20 && ~x10 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x20 && ~x10 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x20 && ~x10 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x20 && ~x10 && ~x17 )
						nx_state = s1;
					else if( x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( ~x21 && x10 && x12 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x21 && x10 && x12 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x21 && x10 && x12 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x10 && x12 && ~x19 )
						nx_state = s1;
					else if( ~x21 && x10 && ~x12 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x21 && ~x10 && x19 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x21 && ~x10 && x19 && ~x14 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x21 && ~x10 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x10 && ~x19 )
						nx_state = s1;
					else nx_state = s259;
				s260 : if( x60 && x61 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x60 && x61 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x60 && x61 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x60 && x61 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x60 && ~x61 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x60 && ~x61 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x60 && ~x61 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x60 && ~x61 && ~x18 )
						nx_state = s39;
					else if( ~x60 && x61 && x62 )
						nx_state = s1;
					else if( ~x60 && x61 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x60 && x61 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x60 && x61 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( ~x60 && x61 && ~x62 && ~x18 )
						nx_state = s39;
					else if( ~x60 && ~x61 )
						nx_state = s40;
					else nx_state = s260;
				s261 : if( x61 && x60 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x61 && x60 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x61 && x60 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x61 && x60 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x61 && ~x60 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x61 && ~x60 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x61 && ~x60 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x61 && ~x60 && x62 && ~x18 )
						nx_state = s1;
					else if( x61 && ~x60 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x61 && ~x60 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x61 && ~x60 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x61 && ~x60 && ~x62 && ~x18 )
						nx_state = s39;
					else if( ~x61 && x60 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x61 && x60 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x61 && x60 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( ~x61 && x60 && ~x18 )
						nx_state = s39;
					else if( ~x61 && ~x60 && x62 && x19 && x15 && x12 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x61 && ~x60 && x62 && x19 && x15 && x12 && ~x7 )
						begin
							y12 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x61 && ~x60 && x62 && x19 && x15 && ~x12 && x7 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x61 && ~x60 && x62 && x19 && x15 && ~x12 && ~x7 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s263;
						end
					else if( ~x61 && ~x60 && x62 && x19 && ~x15 && x16 && x7 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x61 && ~x60 && x62 && x19 && ~x15 && x16 && x7 && ~x12 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s262;
						end
					else if( ~x61 && ~x60 && x62 && x19 && ~x15 && x16 && ~x7 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s258;
						end
					else if( ~x61 && ~x60 && x62 && x19 && ~x15 && ~x16 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x61 && ~x60 && x62 && x19 && ~x15 && ~x16 && ~x7 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x61 && ~x60 && x62 && ~x19 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y23 = 1'b1;	
							nx_state = s411;
						end
					else if( ~x61 && ~x60 && ~x62 )
						nx_state = s40;
					else nx_state = s261;
				s262 : if( x65 && x61 && x60 && x19 && x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x61 && x60 && x19 && ~x13 && x14 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x65 && x61 && x60 && x19 && ~x13 && ~x14 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x61 && x60 && ~x19 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && x61 && ~x60 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x61 && ~x60 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x65 && x61 && ~x60 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x65 && x61 && ~x60 && x62 && ~x18 )
						nx_state = s1;
					else if( x65 && x61 && ~x60 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x65 && x61 && ~x60 && ~x62 && ~x18 )
						nx_state = s39;
					else if( x65 && ~x61 && x60 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x61 && x60 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x61 && x60 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x65 && ~x61 && x60 && ~x18 )
						nx_state = s39;
					else if( x65 && ~x61 && ~x60 && x62 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s258;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 )
						nx_state = s40;
					else if( ~x65 && x21 && x10 && x5 && x16 && x15 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s399;
						end
					else if( ~x65 && x21 && x10 && x5 && x16 && ~x15 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x21 && x10 && x5 && ~x16 && x17 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s215;
						end
					else if( ~x65 && x21 && x10 && x5 && ~x16 && ~x17 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s215;
						end
					else if( ~x65 && x21 && x10 && ~x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x21 && ~x10 && x16 && x5 && x15 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s215;
						end
					else if( ~x65 && x21 && ~x10 && x16 && x5 && ~x15 )
						begin
							y13 = 1'b1;	y16 = 1'b1;	
							nx_state = s284;
						end
					else if( ~x65 && x21 && ~x10 && x16 && ~x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && x14 && x13 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && x14 && ~x13 && x15 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && x14 && ~x13 && ~x15 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && x14 && ~x13 && ~x15 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && x14 && ~x13 && ~x15 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && x14 && ~x13 && ~x15 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && ~x14 && x15 && x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && ~x14 && x15 && ~x12 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && ~x14 && x15 && ~x12 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && ~x14 && x15 && ~x12 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && ~x14 && x15 && ~x12 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && ~x14 && ~x15 && x11 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && ~x14 && ~x15 && ~x11 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && ~x14 && ~x15 && ~x11 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && ~x14 && ~x15 && ~x11 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && x21 && ~x10 && ~x16 && x17 && ~x14 && ~x15 && ~x11 && ~x9 )
						nx_state = s1;
					else if( ~x65 && x21 && ~x10 && ~x16 && ~x17 && x5 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else if( ~x65 && x21 && ~x10 && ~x16 && ~x17 && ~x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && ~x21 && x22 && x17 && x18 && x10 && x15 )
						begin
							y20 = 1'b1;	
							nx_state = s363;
						end
					else if( ~x65 && ~x21 && x22 && x17 && x18 && x10 && ~x15 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && x14 && x15 && x9 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y16 = 1'b1;	
							y23 = 1'b1;	
							nx_state = s310;
						end
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && x14 && x15 && ~x9 && x7 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && x14 && x15 && ~x9 && ~x7 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && x14 && ~x15 && x8 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && x14 && ~x15 && ~x8 && x7 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && x14 && ~x15 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && ~x14 && x15 && x9 )
						begin
							y6 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && ~x14 && x15 && ~x9 && x8 && x7 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && ~x14 && x15 && ~x9 && x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && ~x14 && x15 && ~x9 && ~x8 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && ~x14 && ~x15 && x8 )
						begin
							y6 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x65 && ~x21 && x22 && x17 && x18 && ~x10 && ~x14 && ~x15 && ~x8 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && ~x21 && x22 && x17 && ~x18 && x14 && x10 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s335;
						end
					else if( ~x65 && ~x21 && x22 && x17 && ~x18 && x14 && ~x10 && x15 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s410;
						end
					else if( ~x65 && ~x21 && x22 && x17 && ~x18 && x14 && ~x10 && ~x15 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && ~x21 && x22 && x17 && ~x18 && ~x14 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( ~x65 && ~x21 && x22 && x17 && ~x18 && ~x14 && ~x2 && x5 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s226;
						end
					else if( ~x65 && ~x21 && x22 && x17 && ~x18 && ~x14 && ~x2 && ~x5 && x15 && x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s219;
						end
					else if( ~x65 && ~x21 && x22 && x17 && ~x18 && ~x14 && ~x2 && ~x5 && x15 && ~x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s309;
						end
					else if( ~x65 && ~x21 && x22 && x17 && ~x18 && ~x14 && ~x2 && ~x5 && ~x15 && x10 )
						begin
							y2 = 1'b1;	y16 = 1'b1;	y24 = 1'b1;	
							nx_state = s124;
						end
					else if( ~x65 && ~x21 && x22 && x17 && ~x18 && ~x14 && ~x2 && ~x5 && ~x15 && ~x10 )
						begin
							y14 = 1'b1;	y16 = 1'b1;	
							nx_state = s216;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && x2 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && x10 && x5 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s226;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && x10 && ~x5 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s219;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && x14 && x15 && x5 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s226;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && x14 && x15 && ~x5 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && x14 && ~x15 && x13 && x5 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s226;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && x14 && ~x15 && x13 && ~x5 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && x14 && ~x15 && ~x13 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && x14 && ~x15 && ~x13 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && x14 && ~x15 && ~x13 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && x14 && ~x15 && ~x13 && ~x7 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && x15 && x12 && x5 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s226;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && x15 && x12 && ~x5 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && x15 && ~x12 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && x15 && ~x12 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && x15 && ~x12 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && x15 && ~x12 && ~x7 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && ~x15 && x11 && x5 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s226;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && ~x15 && x11 && ~x5 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && ~x15 && ~x11 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && ~x15 && ~x11 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && ~x15 && ~x11 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && x18 && ~x10 && ~x14 && ~x15 && ~x11 && ~x7 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && ~x18 && x5 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && ~x18 && ~x5 && x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s219;
						end
					else if( ~x65 && ~x21 && x22 && ~x17 && ~x2 && ~x18 && ~x5 && ~x10 )
						begin
							y9 = 1'b1;	y15 = 1'b1;	
							nx_state = s311;
						end
					else if( ~x65 && ~x21 && ~x22 )
						nx_state = s1;
					else nx_state = s262;
				s263 : if( x60 && x61 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x60 && ~x61 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x60 && ~x61 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x60 && ~x61 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( x60 && ~x61 && ~x18 )
						nx_state = s39;
					else if( ~x60 && x61 && x62 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x60 && x61 && x62 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x60 && x61 && x62 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( ~x60 && x61 && x62 && ~x18 )
						nx_state = s1;
					else if( ~x60 && x61 && ~x62 && x18 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x60 && x61 && ~x62 && x18 && ~x13 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x60 && x61 && ~x62 && x18 && ~x13 && ~x14 )
						nx_state = s39;
					else if( ~x60 && x61 && ~x62 && ~x18 )
						nx_state = s39;
					else if( ~x60 && ~x61 )
						nx_state = s40;
					else nx_state = s263;
				s264 : if( x65 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s68;
						end
					else if( ~x65 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s370;
						end
					else nx_state = s264;
				s265 : if( x21 )
						nx_state = s1;
					else if( ~x21 && x22 && x12 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x21 && x22 && ~x12 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x21 && x22 && ~x12 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x21 && x22 && ~x12 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x12 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x7 && x18 && x15 )
						begin
							y8 = 1'b1;	y18 = 1'b1;	
							nx_state = s82;
						end
					else if( ~x21 && ~x22 && x7 && x18 && ~x15 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s374;
						end
					else if( ~x21 && ~x22 && x7 && ~x18 && x19 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s320;
						end
					else if( ~x21 && ~x22 && x7 && ~x18 && x19 && ~x15 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x21 && ~x22 && x7 && ~x18 && ~x19 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x21 && ~x22 && ~x7 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s385;
						end
					else nx_state = s265;
				s266 : if( x21 )
						nx_state = s1;
					else if( ~x21 && x22 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x21 && x22 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x21 && x22 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && ~x22 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && ~x22 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x8 )
						nx_state = s1;
					else nx_state = s266;
				s267 : if( x65 && x2 && x18 && x19 && x14 && x17 && x20 && x16 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x65 && x2 && x18 && x19 && x14 && x17 && x20 && ~x16 )
						begin
							y24 = 1'b1;	
							nx_state = s346;
						end
					else if( x65 && x2 && x18 && x19 && x14 && x17 && ~x20 && x16 )
						begin
							y13 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	y29 = 1'b1;	y30 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s347;
						end
					else if( x65 && x2 && x18 && x19 && x14 && x17 && ~x20 && ~x16 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x65 && x2 && x18 && x19 && x14 && ~x17 && x20 && x8 && x16 )
						begin
							y13 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	y29 = 1'b1;	y30 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s347;
						end
					else if( x65 && x2 && x18 && x19 && x14 && ~x17 && x20 && x8 && ~x16 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && x18 && x19 && x14 && ~x17 && x20 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && x18 && x19 && x14 && ~x17 && ~x20 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && x15 && x17 && x20 && x16 )
						begin
							y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && x15 && x17 && x20 && ~x16 )
						begin
							y4 = 1'b1;	y12 = 1'b1;	y27 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && x15 && x17 && ~x20 && x16 )
						begin
							y24 = 1'b1;	
							nx_state = s346;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && x15 && x17 && ~x20 && ~x16 )
						begin
							y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && x15 && ~x17 && x16 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && x15 && ~x17 && ~x16 && x13 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && x15 && ~x17 && ~x16 && ~x13 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && x15 && ~x17 && ~x16 && ~x13 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && x15 && ~x17 && ~x16 && ~x13 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && x18 && x19 && ~x14 && x15 && ~x17 && ~x16 && ~x13 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && x17 && x16 && x7 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && x17 && x16 && ~x7 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && x17 && x16 && ~x7 && x5 && ~x6 )
						nx_state = s1;
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && x17 && x16 && ~x7 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && x17 && ~x16 && x6 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && x17 && ~x16 && ~x6 && x5 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && x17 && ~x16 && ~x6 && x5 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && x17 && ~x16 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && ~x17 && x16 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && ~x17 && x16 && ~x12 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && ~x17 && x16 && ~x12 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && ~x17 && x16 && ~x12 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && ~x17 && x16 && ~x12 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && ~x17 && ~x16 && x11 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && ~x17 && ~x16 && ~x11 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && ~x17 && ~x16 && ~x11 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && ~x17 && ~x16 && ~x11 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && x18 && x19 && ~x14 && ~x15 && ~x17 && ~x16 && ~x11 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && x17 && x20 && x14 && x13 )
						begin
							y10 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s349;
						end
					else if( x65 && x2 && x18 && ~x19 && x17 && x20 && x14 && ~x13 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x65 && x2 && x18 && ~x19 && x17 && x20 && ~x14 && x13 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	y19 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s349;
						end
					else if( x65 && x2 && x18 && ~x19 && x17 && x20 && ~x14 && ~x13 && x6 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s102;
						end
					else if( x65 && x2 && x18 && ~x19 && x17 && x20 && ~x14 && ~x13 && ~x6 && x5 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && x18 && ~x19 && x17 && x20 && ~x14 && ~x13 && ~x6 && x5 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && x17 && x20 && ~x14 && ~x13 && ~x6 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && x17 && ~x20 && x15 && x14 )
						begin
							y10 = 1'b1;	y19 = 1'b1;	y21 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s349;
						end
					else if( x65 && x2 && x18 && ~x19 && x17 && ~x20 && x15 && ~x14 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s102;
						end
					else if( x65 && x2 && x18 && ~x19 && x17 && ~x20 && ~x15 && x14 )
						begin
							y15 = 1'b1;	y28 = 1'b1;	
							nx_state = s350;
						end
					else if( x65 && x2 && x18 && ~x19 && x17 && ~x20 && ~x15 && ~x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && x13 && x12 && x14 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && x13 && x12 && ~x14 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && x13 && x12 && ~x14 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && x13 && x12 && ~x14 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && x13 && x12 && ~x14 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && x13 && ~x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && ~x13 && x11 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && ~x13 && x11 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && ~x13 && x11 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && ~x13 && x11 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && ~x17 && x20 && ~x13 && ~x11 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && x15 && x12 && x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s241;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && x15 && x12 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && x15 && ~x12 && x14 && x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s241;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && x15 && ~x12 && x14 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && x15 && ~x12 && ~x14 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && x15 && ~x12 && ~x14 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && x15 && ~x12 && ~x14 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && x15 && ~x12 && ~x14 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && x14 && x13 && x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s241;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && x14 && x13 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && x14 && ~x13 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && x14 && ~x13 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && x14 && ~x13 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && x14 && ~x13 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && ~x14 && x11 && x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s241;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && ~x14 && x11 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && ~x14 && ~x11 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && ~x14 && ~x11 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && ~x14 && ~x11 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && x18 && ~x19 && ~x17 && ~x20 && ~x15 && ~x14 && ~x11 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && ~x18 && x17 && x19 && x15 && x14 && x20 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && x15 && x14 && ~x20 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && x15 && ~x14 && x16 && x20 && x13 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && x15 && ~x14 && x16 && x20 && ~x13 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	y32 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && x15 && ~x14 && x16 && ~x20 && x13 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && x15 && ~x14 && x16 && ~x20 && ~x13 )
						begin
							y4 = 1'b1;	y29 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && x15 && ~x14 && ~x16 && x20 )
						begin
							y4 = 1'b1;	y29 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && x15 && ~x14 && ~x16 && ~x20 && x4 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	y28 = 1'b1;	
							nx_state = s348;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && x15 && ~x14 && ~x16 && ~x20 && ~x4 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && ~x15 && x14 && x16 && x20 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && ~x15 && x14 && x16 && ~x20 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && ~x15 && x14 && ~x16 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && ~x15 && ~x14 && x20 && x8 && x16 )
						begin
							y4 = 1'b1;	y18 = 1'b1;	y29 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && ~x15 && ~x14 && x20 && x8 && ~x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && ~x15 && ~x14 && x20 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && ~x15 && ~x14 && ~x20 && x8 && x16 )
						begin
							y4 = 1'b1;	y17 = 1'b1;	y29 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && ~x15 && ~x14 && ~x20 && x8 && ~x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	y21 = 1'b1;	y28 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && x19 && ~x15 && ~x14 && ~x20 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && x16 && x14 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	y21 = 1'b1;	y28 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && x16 && ~x14 && x15 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && x16 && ~x14 && x15 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && x16 && ~x14 && x15 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && x16 && ~x14 && x15 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && x16 && ~x14 && ~x15 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && ~x16 && x13 && x14 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	y21 = 1'b1;	y28 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && ~x16 && x13 && x14 && ~x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && ~x16 && x13 && ~x14 && x4 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && ~x16 && x13 && ~x14 && ~x4 )
						begin
							y4 = 1'b1;	y12 = 1'b1;	y27 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && ~x16 && ~x13 && x8 )
						begin
							y13 = 1'b1;	y20 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	y29 = 1'b1;	y30 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s347;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && x20 && ~x16 && ~x13 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && x14 && x16 )
						begin
							y24 = 1'b1;	
							nx_state = s346;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && x14 && ~x16 && x15 && x13 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && x14 && ~x16 && x15 && ~x13 )
						begin
							y4 = 1'b1;	y12 = 1'b1;	y27 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && x14 && ~x16 && ~x15 )
						begin
							y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && ~x14 && x15 && x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && ~x14 && x15 && ~x16 && x8 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							y19 = 1'b1;	y21 = 1'b1;	y28 = 1'b1;	
							nx_state = s351;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && ~x14 && x15 && ~x16 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && ~x14 && ~x15 && x8 && x16 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && ~x14 && ~x15 && x8 && x16 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && ~x14 && ~x15 && x8 && x16 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && ~x14 && ~x15 && x8 && x16 && ~x5 )
						nx_state = s1;
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && ~x14 && ~x15 && x8 && ~x16 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	y19 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s349;
						end
					else if( x65 && x2 && ~x18 && x17 && ~x19 && ~x20 && ~x14 && ~x15 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && x2 && ~x18 && ~x17 && x8 )
						begin
							y4 = 1'b1;	y18 = 1'b1;	
							nx_state = s395;
						end
					else if( x65 && x2 && ~x18 && ~x17 && ~x8 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y28 = 1'b1;	
							nx_state = s412;
						end
					else if( x65 && ~x2 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x65 && x21 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x65 && x21 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x65 && x21 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x65 && ~x21 && x22 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x65 && ~x21 && x22 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x21 && ~x22 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && ~x21 && ~x22 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x65 && ~x21 && ~x22 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x65 && ~x21 && ~x22 && ~x8 )
						nx_state = s1;
					else nx_state = s267;
				s268 : if( 1'b1 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else nx_state = s268;
				s269 : if( x21 && x66 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x21 && x66 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x21 && x66 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x21 && x66 && ~x19 )
						nx_state = s1;
					else if( x21 && ~x66 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( x21 && ~x66 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( x21 && ~x66 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x21 && ~x66 && ~x3 )
						nx_state = s1;
					else if( ~x21 && x66 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x21 && x66 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x21 && x66 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x21 && x66 && ~x20 )
						nx_state = s1;
					else if( ~x21 && ~x66 && x22 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x21 && ~x66 && x22 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x21 && ~x66 && x22 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x66 && x22 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x66 && ~x22 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && ~x66 && ~x22 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && ~x66 && ~x22 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && ~x66 && ~x22 && ~x8 )
						nx_state = s1;
					else nx_state = s269;
				s270 : if( x21 )
						begin
							y18 = 1'b1;	
							nx_state = s394;
						end
					else if( ~x21 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x21 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x21 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x6 )
						nx_state = s1;
					else nx_state = s270;
				s271 : if( 1'b1 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else nx_state = s271;
				s272 : if( x21 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x21 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else nx_state = s272;
				s273 : if( x21 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( x21 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( x21 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( x21 && ~x3 )
						nx_state = s1;
					else if( ~x21 && x22 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x21 && x22 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x21 && x22 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && ~x22 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && ~x22 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x8 )
						nx_state = s1;
					else nx_state = s273;
				s274 : if( x21 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x21 && x22 && x5 && x18 && x17 && x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x21 && x22 && x5 && x18 && x17 && ~x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x21 && x22 && x5 && x18 && ~x17 && x12 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s386;
						end
					else if( ~x21 && x22 && x5 && x18 && ~x17 && ~x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s374;
						end
					else if( ~x21 && x22 && x5 && ~x18 && x19 && x12 && x17 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x21 && x22 && x5 && ~x18 && x19 && x12 && ~x17 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x21 && x22 && x5 && ~x18 && x19 && ~x12 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x21 && x22 && x5 && ~x18 && ~x19 && x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x21 && x22 && x5 && ~x18 && ~x19 && ~x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && x22 && ~x5 )
						begin
							y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s376;
						end
					else if( ~x21 && ~x22 && x18 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && ~x22 && x18 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && ~x22 && x18 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x18 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x18 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else nx_state = s274;
				s275 : if( x21 && x19 && x18 && x17 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s272;
						end
					else if( x21 && x19 && x18 && x17 && ~x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s272;
						end
					else if( x21 && x19 && x18 && ~x17 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x21 && x19 && x18 && ~x17 && ~x12 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x21 && x19 && ~x18 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s274;
						end
					else if( x21 && ~x19 && x9 && x20 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s272;
						end
					else if( x21 && ~x19 && x9 && x20 && ~x12 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s105;
						end
					else if( x21 && ~x19 && x9 && ~x20 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s270;
						end
					else if( x21 && ~x19 && x9 && ~x20 && ~x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s109;
						end
					else if( x21 && ~x19 && ~x9 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s274;
						end
					else if( ~x21 && x22 && x3 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s274;
						end
					else if( ~x21 && x22 && ~x3 && x5 && x18 && x17 && x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x21 && x22 && ~x3 && x5 && x18 && x17 && ~x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x21 && x22 && ~x3 && x5 && x18 && ~x17 && x12 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s386;
						end
					else if( ~x21 && x22 && ~x3 && x5 && x18 && ~x17 && ~x12 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s374;
						end
					else if( ~x21 && x22 && ~x3 && x5 && ~x18 && x19 && x12 && x17 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x21 && x22 && ~x3 && x5 && ~x18 && x19 && x12 && ~x17 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s388;
						end
					else if( ~x21 && x22 && ~x3 && x5 && ~x18 && x19 && ~x12 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x21 && x22 && ~x3 && x5 && ~x18 && ~x19 && x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s271;
						end
					else if( ~x21 && x22 && ~x3 && x5 && ~x18 && ~x19 && ~x12 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x21 && x22 && ~x3 && ~x5 )
						begin
							y14 = 1'b1;	y18 = 1'b1;	
							nx_state = s376;
						end
					else if( ~x21 && ~x22 && x18 && x15 )
						begin
							y8 = 1'b1;	y18 = 1'b1;	
							nx_state = s82;
						end
					else if( ~x21 && ~x22 && x18 && ~x15 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s374;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && x15 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s413;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && x15 && ~x5 )
						begin
							y3 = 1'b1;	
							nx_state = s320;
						end
					else if( ~x21 && ~x22 && ~x18 && x19 && ~x15 )
						begin
							y4 = 1'b1;	y21 = 1'b1;	
							nx_state = s273;
						end
					else if( ~x21 && ~x22 && ~x18 && ~x19 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else nx_state = s275;
				s276 : if( x16 && x15 && x10 && x12 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x16 && x15 && x10 && ~x12 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( x16 && x15 && ~x10 && x11 && x12 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s126;
						end
					else if( x16 && x15 && ~x10 && x11 && ~x12 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s192;
						end
					else if( x16 && x15 && ~x10 && ~x11 && x12 && x13 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s125;
						end
					else if( x16 && x15 && ~x10 && ~x11 && x12 && ~x13 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x16 && x15 && ~x10 && ~x11 && x12 && ~x13 && x17 && ~x14 )
						nx_state = s1;
					else if( x16 && x15 && ~x10 && ~x11 && x12 && ~x13 && ~x17 )
						nx_state = s1;
					else if( x16 && x15 && ~x10 && ~x11 && ~x12 && x14 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s125;
						end
					else if( x16 && x15 && ~x10 && ~x11 && ~x12 && ~x14 && x17 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x16 && x15 && ~x10 && ~x11 && ~x12 && ~x14 && x17 && ~x13 )
						nx_state = s1;
					else if( x16 && x15 && ~x10 && ~x11 && ~x12 && ~x14 && ~x17 )
						nx_state = s1;
					else if( x16 && ~x15 && x12 && x10 && x8 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x16 && ~x15 && x12 && x10 && x8 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x16 && ~x15 && x12 && x10 && x8 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x16 && ~x15 && x12 && x10 && x8 && ~x17 )
						nx_state = s1;
					else if( x16 && ~x15 && x12 && x10 && ~x8 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x16 && ~x15 && x12 && x10 && ~x8 && ~x5 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s132;
						end
					else if( x16 && ~x15 && x12 && x10 && ~x8 && ~x5 && ~x2 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s199;
						end
					else if( x16 && ~x15 && x12 && ~x10 && x11 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x16 && ~x15 && x12 && ~x10 && x11 && ~x5 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s132;
						end
					else if( x16 && ~x15 && x12 && ~x10 && x11 && ~x5 && ~x2 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s199;
						end
					else if( x16 && ~x15 && x12 && ~x10 && ~x11 && x7 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x16 && ~x15 && x12 && ~x10 && ~x11 && x7 && ~x5 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s132;
						end
					else if( x16 && ~x15 && x12 && ~x10 && ~x11 && x7 && ~x5 && ~x2 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s199;
						end
					else if( x16 && ~x15 && x12 && ~x10 && ~x11 && ~x7 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x16 && ~x15 && x12 && ~x10 && ~x11 && ~x7 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x16 && ~x15 && x12 && ~x10 && ~x11 && ~x7 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x16 && ~x15 && x12 && ~x10 && ~x11 && ~x7 && ~x17 )
						nx_state = s1;
					else if( x16 && ~x15 && ~x12 && x10 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x16 && ~x15 && ~x12 && x10 && ~x5 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s200;
						end
					else if( x16 && ~x15 && ~x12 && x10 && ~x5 && ~x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s132;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && x11 && x9 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && x11 && x9 && ~x5 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s132;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && x11 && x9 && ~x5 && ~x2 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s199;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x16 && ~x15 && ~x12 && ~x10 && x11 && ~x9 && ~x17 )
						nx_state = s1;
					else if( x16 && ~x15 && ~x12 && ~x10 && ~x11 && x8 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && ~x11 && x8 && ~x5 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s132;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && ~x11 && x8 && ~x5 && ~x2 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s199;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x16 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x16 && ~x15 && ~x12 && ~x10 && ~x11 && ~x8 && ~x17 )
						nx_state = s1;
					else if( ~x16 && x15 && x10 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x16 && x15 && x10 && ~x5 && x11 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s132;
						end
					else if( ~x16 && x15 && x10 && ~x5 && x11 && ~x2 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x16 && x15 && x10 && ~x5 && ~x11 && x12 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s132;
						end
					else if( ~x16 && x15 && x10 && ~x5 && ~x11 && x12 && ~x2 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s193;
						end
					else if( ~x16 && x15 && x10 && ~x5 && ~x11 && ~x12 && x2 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s195;
						end
					else if( ~x16 && x15 && x10 && ~x5 && ~x11 && ~x12 && ~x2 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y13 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x16 && x15 && ~x10 && x11 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x16 && x15 && ~x10 && ~x11 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x16 && x15 && ~x10 && ~x11 && ~x5 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s132;
						end
					else if( ~x16 && x15 && ~x10 && ~x11 && ~x5 && ~x2 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x16 && x15 && ~x10 && ~x11 && ~x5 && ~x2 && ~x12 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x16 && ~x15 && x5 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	
							nx_state = s10;
						end
					else if( ~x16 && ~x15 && ~x5 && x2 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s132;
						end
					else if( ~x16 && ~x15 && ~x5 && ~x2 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s390;
						end
					else nx_state = s276;
				s277 : if( x20 && x17 && x15 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s198;
						end
					else if( x20 && x17 && ~x15 && x16 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s59;
						end
					else if( x20 && x17 && ~x15 && ~x16 )
						begin
							y7 = 1'b1;	y12 = 1'b1;	
							nx_state = s211;
						end
					else if( x20 && ~x17 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	y22 = 1'b1;	
							nx_state = s401;
						end
					else if( ~x20 && x21 )
						begin
							y12 = 1'b1;	y15 = 1'b1;	y22 = 1'b1;	
							nx_state = s401;
						end
					else if( ~x20 && ~x21 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s186;
						end
					else nx_state = s277;
				s278 : if( x65 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x4 )
						nx_state = s1;
					else if( ~x65 && x67 && x24 && x26 )
						nx_state = s1;
					else if( ~x65 && x67 && x24 && ~x26 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && x67 && x24 && ~x26 && ~x4 && x19 && x16 && x11 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s188;
						end
					else if( ~x65 && x67 && x24 && ~x26 && ~x4 && x19 && x16 && x11 && ~x12 && x13 )
						begin
							y6 = 1'b1;	
							nx_state = s172;
						end
					else if( ~x65 && x67 && x24 && ~x26 && ~x4 && x19 && x16 && x11 && ~x12 && ~x13 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x65 && x67 && x24 && ~x26 && ~x4 && x19 && x16 && ~x11 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x65 && x67 && x24 && ~x26 && ~x4 && x19 && ~x16 && x17 && x11 && x13 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else if( ~x65 && x67 && x24 && ~x26 && ~x4 && x19 && ~x16 && x17 && x11 && ~x13 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s46;
						end
					else if( ~x65 && x67 && x24 && ~x26 && ~x4 && x19 && ~x16 && x17 && ~x11 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else if( ~x65 && x67 && x24 && ~x26 && ~x4 && x19 && ~x16 && ~x17 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x65 && x67 && x24 && ~x26 && ~x4 && ~x19 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && x67 && ~x24 && x25 && x26 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( ~x65 && x67 && ~x24 && x25 && ~x26 && x15 && x10 && x11 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s187;
						end
					else if( ~x65 && x67 && ~x24 && x25 && ~x26 && x15 && x10 && ~x11 && x12 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s185;
						end
					else if( ~x65 && x67 && ~x24 && x25 && ~x26 && x15 && x10 && ~x11 && ~x12 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s160;
						end
					else if( ~x65 && x67 && ~x24 && x25 && ~x26 && x15 && ~x10 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x65 && x67 && ~x24 && x25 && ~x26 && ~x15 && x16 && x10 && x12 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x65 && x67 && ~x24 && x25 && ~x26 && ~x15 && x16 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && x67 && ~x24 && x25 && ~x26 && ~x15 && x16 && ~x10 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x65 && x67 && ~x24 && x25 && ~x26 && ~x15 && ~x16 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x65 && x67 && ~x24 && ~x25 )
						nx_state = s1;
					else if( ~x65 && ~x67 && x21 && x9 && x3 )
						nx_state = s40;
					else if( ~x65 && ~x67 && x21 && x9 && ~x3 && x4 )
						nx_state = s40;
					else if( ~x65 && ~x67 && x21 && x9 && ~x3 && ~x4 )
						nx_state = s1;
					else if( ~x65 && ~x67 && x21 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && x22 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 && ~x67 && ~x21 && x22 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && x22 && ~x5 )
						nx_state = s1;
					else if( ~x65 && ~x67 && ~x21 && ~x22 )
						nx_state = s1;
					else nx_state = s278;
				s279 : if( x66 && x21 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( x66 && ~x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s344;
						end
					else if( ~x66 && x68 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x66 && ~x68 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s402;
						end
					else nx_state = s279;
				s280 : if( 1'b1 )
						begin
							y8 = 1'b1;	y17 = 1'b1;	y23 = 1'b1;	
							nx_state = s164;
						end
					else nx_state = s280;
				s281 : if( x24 && x26 )
						begin
							y17 = 1'b1;	
							nx_state = s150;
						end
					else if( x24 && ~x26 && x16 && x11 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s188;
						end
					else if( x24 && ~x26 && x16 && x11 && ~x12 && x13 )
						begin
							y6 = 1'b1;	
							nx_state = s172;
						end
					else if( x24 && ~x26 && x16 && x11 && ~x12 && ~x13 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x24 && ~x26 && x16 && ~x11 )
						begin
							y5 = 1'b1;	y14 = 1'b1;	y22 = 1'b1;	
							nx_state = s160;
						end
					else if( x24 && ~x26 && ~x16 && x17 && x11 && x13 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else if( x24 && ~x26 && ~x16 && x17 && x11 && ~x13 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s46;
						end
					else if( x24 && ~x26 && ~x16 && x17 && ~x11 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else if( x24 && ~x26 && ~x16 && ~x17 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x24 && x25 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else if( ~x24 && ~x25 && x26 && x16 && x11 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x24 && ~x25 && x26 && x16 && ~x11 && x12 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x24 && ~x25 && x26 && x16 && ~x11 && ~x12 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x24 && ~x25 && x26 && x16 && ~x11 && ~x12 && ~x10 )
						begin
							y12 = 1'b1;	y14 = 1'b1;	
							nx_state = s49;
						end
					else if( ~x24 && ~x25 && x26 && ~x16 && x17 && x10 && x12 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x24 && ~x25 && x26 && ~x16 && x17 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x24 && ~x25 && x26 && ~x16 && x17 && ~x10 )
						begin
							y13 = 1'b1;	y15 = 1'b1;	
							nx_state = s166;
						end
					else if( ~x24 && ~x25 && x26 && ~x16 && ~x17 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x24 && ~x25 && ~x26 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else nx_state = s281;
				s282 : if( x24 && x26 && x18 && x15 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( x24 && x26 && x18 && ~x15 && x14 )
						begin
							y6 = 1'b1;	y12 = 1'b1;	
							nx_state = s162;
						end
					else if( x24 && x26 && x18 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x24 && x26 && ~x18 )
						nx_state = s1;
					else if( x24 && ~x26 && x20 && x15 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( x24 && ~x26 && x20 && ~x15 && x14 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( x24 && ~x26 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x24 && ~x26 && ~x20 )
						nx_state = s1;
					else if( ~x24 && x25 && x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x25 && x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( ~x24 && x25 && x19 && ~x14 && ~x13 && x26 )
						nx_state = s282;
					else if( ~x24 && x25 && x19 && ~x14 && ~x13 && ~x26 )
						nx_state = s1;
					else if( ~x24 && x25 && ~x19 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && x18 && x14 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && x13 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x24 && ~x25 && x26 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && x26 && ~x18 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && x10 && x12 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x24 && ~x25 && ~x26 && x10 && x12 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x24 && ~x25 && ~x26 && x10 && x12 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && x10 && x12 && ~x17 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && x10 && ~x12 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x10 && x17 && x14 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x10 && x17 && ~x14 && x13 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x24 && ~x25 && ~x26 && ~x10 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x24 && ~x25 && ~x26 && ~x10 && ~x17 )
						nx_state = s1;
					else nx_state = s282;
				s283 : if( x65 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s54;
						end
					else if( ~x65 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else nx_state = s283;
				s284 : if( x21 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x21 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x21 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x21 && ~x9 )
						nx_state = s1;
					else if( ~x21 && x22 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && ~x22 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else nx_state = s284;
				s285 : if( x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x18 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x21 && x22 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x21 && x22 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x17 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && x18 && x14 )
						nx_state = s40;
					else if( ~x21 && x22 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s40;
					else if( ~x21 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x21 && ~x22 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s180;
						end
					else nx_state = s285;
				s286 : if( x65 && x60 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s314;
						end
					else if( x65 && ~x60 )
						begin
							y11 = 1'b1;	
							nx_state = s356;
						end
					else if( ~x65 && x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x65 && x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x65 && x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x23 && x10 && x12 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x21 && x22 && x23 && x10 && x12 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x21 && x22 && x23 && x10 && x12 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x23 && x10 && x12 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x23 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s341;
						end
					else if( ~x65 && ~x21 && x22 && x23 && ~x10 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x21 && x22 && x23 && ~x10 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x65 && ~x21 && x22 && x23 && ~x10 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && x23 && ~x10 && ~x17 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x23 && x18 && x14 )
						nx_state = s40;
					else if( ~x65 && ~x21 && x22 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s40;
					else if( ~x65 && ~x21 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x65 && ~x21 && ~x22 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s180;
						end
					else nx_state = s286;
				s287 : if( 1'b1 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y19 = 1'b1;	
							nx_state = s226;
						end
					else nx_state = s287;
				s288 : if( x65 && x22 && x21 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x22 && x21 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x22 && x21 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && x22 && x21 && ~x4 )
						nx_state = s1;
					else if( x65 && x22 && ~x21 && x18 && x19 )
						nx_state = s1;
					else if( x65 && x22 && ~x21 && x18 && ~x19 && x10 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( x65 && x22 && ~x21 && x18 && ~x19 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x22 && ~x21 && x18 && ~x19 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x22 && ~x21 && x18 && ~x19 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && x22 && ~x21 && x18 && ~x19 && ~x10 && ~x4 )
						nx_state = s1;
					else if( x65 && x22 && ~x21 && ~x18 && x19 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x22 && ~x21 && ~x18 && x19 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x22 && ~x21 && ~x18 && x19 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && x22 && ~x21 && ~x18 && ~x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x22 && ~x21 && ~x18 && ~x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x22 && ~x21 && ~x18 && ~x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && x22 && ~x21 && ~x18 && ~x19 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x22 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x22 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && ~x22 && ~x4 )
						nx_state = s1;
					else if( ~x65 && x21 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x21 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x21 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( ~x65 && x21 && ~x9 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x22 )
						nx_state = s1;
					else if( ~x65 && ~x21 && ~x22 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x65 && ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x65 && ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s288;
				s289 : if( 1'b1 )
						begin
							y12 = 1'b1;	
							nx_state = s210;
						end
					else nx_state = s289;
				s290 : if( x65 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x65 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else nx_state = s290;
				s291 : if( x65 && x60 )
						nx_state = s73;
					else if( x65 && ~x60 && x61 )
						nx_state = s73;
					else if( x65 && ~x60 && ~x61 )
						nx_state = s40;
					else if( ~x65 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else nx_state = s291;
				s292 : if( x65 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x65 )
						begin
							y17 = 1'b1;	
							nx_state = s17;
						end
					else nx_state = s292;
				s293 : if( x66 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x66 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else nx_state = s293;
				s294 : if( x21 )
						begin
							y35 = 1'b1;	
							nx_state = s26;
						end
					else if( ~x21 && x23 && x22 )
						begin
							y20 = 1'b1;	
							nx_state = s363;
						end
					else if( ~x21 && x23 && ~x22 )
						begin
							y35 = 1'b1;	
							nx_state = s26;
						end
					else if( ~x21 && ~x23 && x22 && x17 && x15 && x9 )
						begin
							y4 = 1'b1;	y7 = 1'b1;	
							nx_state = s119;
						end
					else if( ~x21 && ~x23 && x22 && x17 && x15 && ~x9 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( ~x21 && ~x23 && x22 && x17 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( ~x21 && ~x23 && x22 && x17 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x21 && ~x23 && x22 && ~x17 )
						begin
							y35 = 1'b1;	
							nx_state = s26;
						end
					else if( ~x21 && ~x23 && ~x22 && x2 )
						begin
							y35 = 1'b1;	
							nx_state = s26;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x2 && x17 && x15 && x9 )
						begin
							y6 = 1'b1;	
							nx_state = s91;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x2 && x17 && x15 && ~x9 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x2 && x17 && ~x15 && x16 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x2 && x17 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							y30 = 1'b1;	
							nx_state = s205;
						end
					else if( ~x21 && ~x23 && ~x22 && ~x2 && ~x17 )
						begin
							y36 = 1'b1;	
							nx_state = s55;
						end
					else nx_state = s294;
				s295 : if( 1'b1 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	y11 = 1'b1;	
							nx_state = s240;
						end
					else nx_state = s295;
				s296 : if( x66 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x66 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else nx_state = s296;
				s297 : if( x66 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x66 && x24 )
						begin
							y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s182;
						end
					else if( ~x66 && ~x24 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else nx_state = s297;
				s298 : if( x65 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	y24 = 1'b1;	
							nx_state = s99;
						end
					else if( ~x65 && x63 && x1 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y28 = 1'b1;	
							nx_state = s156;
						end
					else if( ~x65 && x63 && ~x1 && x18 && x15 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x65 && x63 && ~x1 && x18 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x65 && x63 && ~x1 && x18 && ~x15 && x16 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( ~x65 && x63 && ~x1 && x18 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x65 && x63 && ~x1 && ~x18 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	y14 = 1'b1;	
							y29 = 1'b1;	
							nx_state = s152;
						end
					else if( ~x65 && ~x63 )
						begin
							y3 = 1'b1;	y22 = 1'b1;	y37 = 1'b1;	
							nx_state = s397;
						end
					else nx_state = s298;
				s299 : if( 1'b1 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	
							nx_state = s345;
						end
					else nx_state = s299;
				s300 : if( x21 && x66 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x66 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x21 && x66 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && x66 && x20 && ~x17 )
						nx_state = s1;
					else if( x21 && x66 && ~x20 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x21 && ~x66 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x21 && ~x66 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x21 && ~x66 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x21 && ~x66 && ~x4 )
						nx_state = s1;
					else if( ~x21 && x66 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x66 && x22 && x18 && x19 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x66 && x22 && x18 && x19 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x66 && x22 && x18 && x19 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x66 && x22 && x18 && ~x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x66 && x22 && x18 && ~x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x66 && x22 && x18 && ~x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x66 && x22 && x18 && ~x19 && ~x4 )
						nx_state = s1;
					else if( ~x21 && ~x66 && x22 && ~x18 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x66 && x22 && ~x18 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x66 && x22 && ~x18 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x66 && x22 && ~x18 && ~x4 )
						nx_state = s1;
					else if( ~x21 && ~x66 && ~x22 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x66 && ~x22 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x66 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x66 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s300;
				s301 : if( x65 && x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x65 && x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x21 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x65 && x19 )
						begin
							y4 = 1'b1;	y14 = 1'b1;	
							nx_state = s304;
						end
					else if( ~x65 && ~x19 && x20 && x15 && x10 && x11 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s334;
						end
					else if( ~x65 && ~x19 && x20 && x15 && x10 && ~x11 && x12 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s334;
						end
					else if( ~x65 && ~x19 && x20 && x15 && x10 && ~x11 && ~x12 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x65 && ~x19 && x20 && x15 && ~x10 && x12 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x65 && ~x19 && x20 && x15 && ~x10 && x12 && ~x11 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x65 && ~x19 && x20 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x65 && ~x19 && x20 && ~x15 && x16 && x10 && x12 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && ~x19 && x20 && ~x15 && x16 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s341;
						end
					else if( ~x65 && ~x19 && x20 && ~x15 && x16 && ~x10 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && ~x19 && x20 && ~x15 && ~x16 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s81;
						end
					else if( ~x65 && ~x19 && ~x20 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else nx_state = s301;
				s302 : if( x65 && x67 && x22 && x17 && x18 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && x22 && x17 && ~x18 && x19 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && x67 && x22 && x17 && ~x18 && ~x19 )
						nx_state = s1;
					else if( x65 && x67 && x22 && ~x17 )
						nx_state = s1;
					else if( x65 && x67 && ~x22 && x18 && x13 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && x67 && ~x22 && x18 && x13 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x67 && ~x22 && x18 && ~x13 && x12 && x23 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && x67 && ~x22 && x18 && ~x13 && x12 && ~x23 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && x67 && ~x22 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x65 && x67 && ~x22 && ~x18 )
						nx_state = s1;
					else if( x65 && ~x67 && x21 && x20 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x67 && x21 && x20 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x67 && x21 && x20 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && x21 && x20 && ~x17 )
						nx_state = s1;
					else if( x65 && ~x67 && x21 && ~x20 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && ~x67 && x21 && ~x20 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x65 && ~x67 && x21 && ~x20 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x65 && ~x67 && x21 && ~x20 && ~x19 )
						nx_state = s1;
					else if( x65 && ~x67 && ~x21 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s259;
						end
					else if( ~x65 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	y21 = 1'b1;	
							nx_state = s45;
						end
					else nx_state = s302;
				s303 : if( x20 && x21 && x17 && x14 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x20 && x21 && x17 && ~x14 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x20 && x21 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x20 && x21 && ~x17 )
						nx_state = s1;
					else if( x20 && ~x21 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x20 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else nx_state = s303;
				s304 : if( x21 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x21 && x20 && x15 && x10 && x11 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s334;
						end
					else if( ~x21 && x20 && x15 && x10 && ~x11 && x12 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s334;
						end
					else if( ~x21 && x20 && x15 && x10 && ~x11 && ~x12 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x21 && x20 && x15 && ~x10 && x12 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x21 && x20 && x15 && ~x10 && x12 && ~x11 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && x20 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x21 && x20 && ~x15 && x16 && x10 && x12 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x21 && x20 && ~x15 && x16 && x10 && ~x12 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s341;
						end
					else if( ~x21 && x20 && ~x15 && x16 && ~x10 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x21 && x20 && ~x15 && ~x16 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s81;
						end
					else if( ~x21 && ~x20 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else nx_state = s304;
				s305 : if( x68 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x68 && x21 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x68 && ~x21 && x22 && x23 && x15 && x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x68 && ~x21 && x22 && x23 && x15 && ~x10 && x12 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x68 && ~x21 && x22 && x23 && x15 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s285;
						end
					else if( ~x68 && ~x21 && x22 && x23 && ~x15 && x16 && x10 && x12 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x68 && ~x21 && x22 && x23 && ~x15 && x16 && x10 && ~x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x68 && ~x21 && x22 && x23 && ~x15 && x16 && ~x10 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x68 && ~x21 && x22 && x23 && ~x15 && ~x16 )
						nx_state = s40;
					else if( ~x68 && ~x21 && x22 && ~x23 && x6 && x15 && x11 && x10 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s334;
						end
					else if( ~x68 && ~x21 && x22 && ~x23 && x6 && x15 && x11 && ~x10 )
						begin
							y14 = 1'b1;	
							nx_state = s285;
						end
					else if( ~x68 && ~x21 && x22 && ~x23 && x6 && x15 && ~x11 && x12 && x10 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s334;
						end
					else if( ~x68 && ~x21 && x22 && ~x23 && x6 && x15 && ~x11 && x12 && ~x10 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x68 && ~x21 && x22 && ~x23 && x6 && x15 && ~x11 && ~x12 && x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x68 && ~x21 && x22 && ~x23 && x6 && x15 && ~x11 && ~x12 && ~x10 )
						begin
							y14 = 1'b1;	
							nx_state = s285;
						end
					else if( ~x68 && ~x21 && x22 && ~x23 && x6 && ~x15 && x16 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x68 && ~x21 && x22 && ~x23 && x6 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s180;
						end
					else if( ~x68 && ~x21 && x22 && ~x23 && ~x6 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x68 && ~x21 && ~x22 && x23 && x15 && x7 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s81;
						end
					else if( ~x68 && ~x21 && ~x22 && x23 && x15 && ~x7 && x9 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x68 && ~x21 && ~x22 && x23 && x15 && ~x7 && ~x9 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x68 && ~x21 && ~x22 && x23 && ~x15 && x16 && x7 && x9 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x68 && ~x21 && ~x22 && x23 && ~x15 && x16 && x7 && ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x68 && ~x21 && ~x22 && x23 && ~x15 && x16 && ~x7 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x68 && ~x21 && ~x22 && x23 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x68 && ~x21 && ~x22 && ~x23 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s81;
						end
					else nx_state = s305;
				s306 : if( x21 && x20 && x18 && x15 && x10 && x11 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s192;
						end
					else if( x21 && x20 && x18 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s193;
						end
					else if( x21 && x20 && x18 && x15 && x10 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s194;
						end
					else if( x21 && x20 && x18 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s300;
						end
					else if( x21 && x20 && x18 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s192;
						end
					else if( x21 && x20 && x18 && ~x15 && x16 && x10 && x12 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s259;
						end
					else if( x21 && x20 && x18 && ~x15 && x16 && x10 && ~x12 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( x21 && x20 && x18 && ~x15 && x16 && ~x10 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s259;
						end
					else if( x21 && x20 && x18 && ~x15 && ~x16 )
						begin
							y2 = 1'b1;	y5 = 1'b1;	y6 = 1'b1;	
							y7 = 1'b1;	
							nx_state = s134;
						end
					else if( x21 && x20 && ~x18 )
						begin
							y4 = 1'b1;	y16 = 1'b1;	
							nx_state = s307;
						end
					else if( x21 && ~x20 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s199;
						end
					else if( ~x21 && x18 && x15 && x10 && x11 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x21 && x18 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s301;
						end
					else if( ~x21 && x18 && x15 && x10 && ~x11 && ~x12 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s195;
						end
					else if( ~x21 && x18 && x15 && ~x10 && x12 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s197;
						end
					else if( ~x21 && x18 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y10 = 1'b1;	
							nx_state = s192;
						end
					else if( ~x21 && x18 && ~x15 && x16 && x10 && x12 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s259;
						end
					else if( ~x21 && x18 && ~x15 && x16 && x10 && ~x12 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x21 && x18 && ~x15 && x16 && ~x10 )
						begin
							y1 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s259;
						end
					else if( ~x21 && x18 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s303;
						end
					else if( ~x21 && ~x18 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s57;
						end
					else nx_state = s306;
				s307 : if( x21 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s121;
						end
					else if( ~x21 )
						nx_state = s1;
					else nx_state = s307;
				s308 : if( 1'b1 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	y9 = 1'b1;	
							nx_state = s79;
						end
					else nx_state = s308;
				s309 : if( x22 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x22 )
						begin
							y17 = 1'b1;	
							nx_state = s17;
						end
					else nx_state = s309;
				s310 : if( x21 && x9 && x8 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x21 && x9 && ~x8 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( x21 && x9 && ~x8 && ~x7 )
						nx_state = s1;
					else if( x21 && ~x9 )
						nx_state = s1;
					else if( ~x21 && x22 && x8 && x7 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x21 && x22 && x8 && ~x7 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x8 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x4 && x5 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y9 = 1'b1;	y13 = 1'b1;	
							nx_state = s29;
						end
					else if( ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s310;
				s311 : if( x21 && x16 && x15 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s214;
						end
					else if( x21 && x16 && x15 && ~x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s215;
						end
					else if( x21 && x16 && ~x15 && x10 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else if( x21 && x16 && ~x15 && ~x10 )
						begin
							y14 = 1'b1;	y16 = 1'b1;	
							nx_state = s216;
						end
					else if( x21 && ~x16 && x17 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s215;
						end
					else if( x21 && ~x16 && ~x17 && x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s215;
						end
					else if( x21 && ~x16 && ~x17 && ~x10 )
						begin
							y11 = 1'b1;	y14 = 1'b1;	
							nx_state = s218;
						end
					else if( ~x21 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else nx_state = s311;
				s312 : if( 1'b1 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s118;
						end
					else nx_state = s312;
				s313 : if( 1'b1 )
						begin
							y8 = 1'b1;	y22 = 1'b1;	
							nx_state = s267;
						end
					else nx_state = s313;
				s314 : if( x67 && x22 && x15 && x8 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x67 && x22 && x15 && ~x8 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x67 && x22 && ~x15 && x16 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s302;
						end
					else if( x67 && x22 && ~x15 && ~x16 )
						begin
							y11 = 1'b1;	
							nx_state = s122;
						end
					else if( x67 && ~x22 )
						begin
							y10 = 1'b1;	y26 = 1'b1;	y27 = 1'b1;	
							nx_state = s2;
						end
					else if( ~x67 && x60 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	
							nx_state = s154;
						end
					else if( ~x67 && ~x60 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else nx_state = s314;
				s315 : if( 1'b1 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else nx_state = s315;
				s316 : if( x60 )
						nx_state = s1;
					else if( ~x60 && x61 )
						nx_state = s1;
					else if( ~x60 && ~x61 && x62 )
						begin
							y2 = 1'b1;	y19 = 1'b1;	y24 = 1'b1;	
							nx_state = s321;
						end
					else if( ~x60 && ~x61 && ~x62 )
						nx_state = s40;
					else nx_state = s316;
				s317 : if( x21 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x21 && x16 && x10 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s67;
						end
					else if( ~x21 && x16 && ~x10 )
						begin
							y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s113;
						end
					else if( ~x21 && ~x16 && x17 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x21 && ~x16 && ~x17 )
						begin
							y5 = 1'b1;	y17 = 1'b1;	
							nx_state = s115;
						end
					else nx_state = s317;
				s318 : if( 1'b1 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else nx_state = s318;
				s319 : if( x65 && x61 && x60 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s328;
						end
					else if( x65 && x61 && ~x60 && x62 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else if( x65 && x61 && ~x60 && ~x62 && x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s255;
						end
					else if( x65 && x61 && ~x60 && ~x62 && ~x2 && x19 && x15 )
						nx_state = s73;
					else if( x65 && x61 && ~x60 && ~x62 && ~x2 && x19 && ~x15 && x16 )
						begin
							y12 = 1'b1;	
							nx_state = s291;
						end
					else if( x65 && x61 && ~x60 && ~x62 && ~x2 && x19 && ~x15 && ~x16 )
						nx_state = s73;
					else if( x65 && x61 && ~x60 && ~x62 && ~x2 && ~x19 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y24 = 1'b1;	
							nx_state = s64;
						end
					else if( x65 && ~x61 && x60 && x2 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s255;
						end
					else if( x65 && ~x61 && x60 && ~x2 && x19 && x15 )
						nx_state = s73;
					else if( x65 && ~x61 && x60 && ~x2 && x19 && ~x15 && x16 )
						begin
							y12 = 1'b1;	
							nx_state = s291;
						end
					else if( x65 && ~x61 && x60 && ~x2 && x19 && ~x15 && ~x16 )
						nx_state = s73;
					else if( x65 && ~x61 && x60 && ~x2 && ~x19 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y24 = 1'b1;	
							nx_state = s64;
						end
					else if( x65 && ~x61 && ~x60 && x62 )
						nx_state = s40;
					else if( x65 && ~x61 && ~x60 && ~x62 && x5 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s255;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && x15 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && x15 && ~x7 && x11 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && x15 && ~x7 && ~x11 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s254;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && x4 )
						nx_state = s40;
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && ~x4 && x11 && x9 )
						nx_state = s40;
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && ~x4 && x11 && ~x9 && x7 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s128;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && ~x4 && x11 && ~x9 && ~x7 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s118;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && ~x4 && ~x11 && x9 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && ~x4 && ~x11 && x9 && ~x7 && x10 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && ~x4 && ~x11 && x9 && ~x7 && ~x10 )
						nx_state = s40;
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && x7 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && x7 && ~x8 )
						nx_state = s40;
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && ~x7 && x12 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && x16 && ~x4 && ~x11 && ~x9 && ~x7 && ~x12 )
						nx_state = s40;
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && x18 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( x65 && ~x61 && ~x60 && ~x62 && ~x5 && ~x18 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y24 = 1'b1;	
							nx_state = s64;
						end
					else if( ~x65 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s374;
						end
					else nx_state = s319;
				s320 : if( x65 )
						nx_state = s40;
					else if( ~x65 && x66 && x23 && x18 && x15 && x7 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y9 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s81;
						end
					else if( ~x65 && x66 && x23 && x18 && x15 && ~x7 && x9 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x65 && x66 && x23 && x18 && x15 && ~x7 && ~x9 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x65 && x66 && x23 && x18 && ~x15 && x7 && x9 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s330;
						end
					else if( ~x65 && x66 && x23 && x18 && ~x15 && x7 && ~x9 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x65 && x66 && x23 && x18 && ~x15 && ~x7 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s330;
						end
					else if( ~x65 && x66 && x23 && ~x18 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s84;
						end
					else if( ~x65 && x66 && ~x23 && x9 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && x66 && ~x23 && ~x9 && x7 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x65 && x66 && ~x23 && ~x9 && ~x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x65 && ~x66 )
						begin
							y5 = 1'b1;	
							nx_state = s343;
						end
					else nx_state = s320;
				s321 : if( x61 && x16 && x17 && x11 && x13 )
						begin
							y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s260;
						end
					else if( x61 && x16 && x17 && x11 && ~x13 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s261;
						end
					else if( x61 && x16 && x17 && ~x11 && x12 && x13 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s262;
						end
					else if( x61 && x16 && x17 && ~x11 && x12 && ~x13 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s254;
						end
					else if( x61 && x16 && x17 && ~x11 && ~x12 && x13 && x15 )
						begin
							y15 = 1'b1;	
							nx_state = s355;
						end
					else if( x61 && x16 && x17 && ~x11 && ~x12 && x13 && ~x15 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x61 && x16 && x17 && ~x11 && ~x12 && x13 && ~x15 && x18 && ~x14 )
						nx_state = s1;
					else if( x61 && x16 && x17 && ~x11 && ~x12 && x13 && ~x15 && ~x18 )
						nx_state = s1;
					else if( x61 && x16 && x17 && ~x11 && ~x12 && ~x13 && x14 )
						begin
							y15 = 1'b1;	
							nx_state = s355;
						end
					else if( x61 && x16 && x17 && ~x11 && ~x12 && ~x13 && ~x14 && x18 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x61 && x16 && x17 && ~x11 && ~x12 && ~x13 && ~x14 && x18 && ~x15 )
						nx_state = s1;
					else if( x61 && x16 && x17 && ~x11 && ~x12 && ~x13 && ~x14 && ~x18 )
						nx_state = s1;
					else if( x61 && x16 && ~x17 && x12 && x11 && x13 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( x61 && x16 && ~x17 && x12 && x11 && x13 && ~x3 && x2 )
						nx_state = s40;
					else if( x61 && x16 && ~x17 && x12 && x11 && x13 && ~x3 && ~x2 )
						begin
							y22 = 1'b1;	
							nx_state = s224;
						end
					else if( x61 && x16 && ~x17 && x12 && x11 && ~x13 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s255;
						end
					else if( x61 && x16 && ~x17 && x12 && ~x11 && x13 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else if( x61 && x16 && ~x17 && x12 && ~x11 && ~x13 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s263;
						end
					else if( x61 && x16 && ~x17 && ~x12 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( x61 && x16 && ~x17 && ~x12 && ~x3 && x2 )
						nx_state = s40;
					else if( x61 && x16 && ~x17 && ~x12 && ~x3 && ~x2 && x13 && x11 )
						begin
							y22 = 1'b1;	
							nx_state = s58;
						end
					else if( x61 && x16 && ~x17 && ~x12 && ~x3 && ~x2 && x13 && ~x11 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x61 && x16 && ~x17 && ~x12 && ~x3 && ~x2 && ~x13 && x11 )
						begin
							y4 = 1'b1;	y13 = 1'b1;	y24 = 1'b1;	
							nx_state = s64;
						end
					else if( x61 && x16 && ~x17 && ~x12 && ~x3 && ~x2 && ~x13 && ~x11 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x61 && ~x16 && x3 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( x61 && ~x16 && ~x3 && x17 && x13 && x11 && x9 && x2 )
						nx_state = s40;
					else if( x61 && ~x16 && ~x3 && x17 && x13 && x11 && x9 && ~x2 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s252;
						end
					else if( x61 && ~x16 && ~x3 && x17 && x13 && x11 && ~x9 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x61 && ~x16 && ~x3 && x17 && x13 && x11 && ~x9 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x61 && ~x16 && ~x3 && x17 && x13 && x11 && ~x9 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x61 && ~x16 && ~x3 && x17 && x13 && x11 && ~x9 && ~x18 )
						nx_state = s1;
					else if( x61 && ~x16 && ~x3 && x17 && x13 && ~x11 && x12 && x2 )
						nx_state = s40;
					else if( x61 && ~x16 && ~x3 && x17 && x13 && ~x11 && x12 && ~x2 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s252;
						end
					else if( x61 && ~x16 && ~x3 && x17 && x13 && ~x11 && ~x12 && x8 && x2 )
						nx_state = s40;
					else if( x61 && ~x16 && ~x3 && x17 && x13 && ~x11 && ~x12 && x8 && ~x2 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s252;
						end
					else if( x61 && ~x16 && ~x3 && x17 && x13 && ~x11 && ~x12 && ~x8 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x61 && ~x16 && ~x3 && x17 && x13 && ~x11 && ~x12 && ~x8 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x61 && ~x16 && ~x3 && x17 && x13 && ~x11 && ~x12 && ~x8 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x61 && ~x16 && ~x3 && x17 && x13 && ~x11 && ~x12 && ~x8 && ~x18 )
						nx_state = s1;
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && x11 )
						nx_state = s40;
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && x12 && x10 && x2 )
						nx_state = s40;
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && x12 && x10 && ~x2 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s252;
						end
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && x12 && ~x10 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && x12 && ~x10 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && x12 && ~x10 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && x12 && ~x10 && ~x18 )
						nx_state = s1;
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && x7 && x2 )
						nx_state = s40;
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && x7 && ~x2 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s252;
						end
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && ~x7 && x18 && x14 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && ~x7 && x18 && ~x14 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && ~x7 && x18 && ~x14 && ~x15 )
						nx_state = s1;
					else if( x61 && ~x16 && ~x3 && x17 && ~x13 && ~x11 && ~x12 && ~x7 && ~x18 )
						nx_state = s1;
					else if( x61 && ~x16 && ~x3 && ~x17 && x2 )
						nx_state = s40;
					else if( x61 && ~x16 && ~x3 && ~x17 && ~x2 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s74;
						end
					else if( ~x61 && x62 && x2 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y10 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s261;
						end
					else if( ~x61 && x62 && ~x2 && x19 && x15 && x12 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x61 && x62 && ~x2 && x19 && x15 && x12 && ~x7 )
						begin
							y12 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x61 && x62 && ~x2 && x19 && x15 && ~x12 && x7 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x61 && x62 && ~x2 && x19 && x15 && ~x12 && ~x7 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s263;
						end
					else if( ~x61 && x62 && ~x2 && x19 && ~x15 && x16 && x7 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x61 && x62 && ~x2 && x19 && ~x15 && x16 && x7 && ~x12 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s262;
						end
					else if( ~x61 && x62 && ~x2 && x19 && ~x15 && x16 && ~x7 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s258;
						end
					else if( ~x61 && x62 && ~x2 && x19 && ~x15 && ~x16 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x61 && x62 && ~x2 && x19 && ~x15 && ~x16 && ~x7 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x61 && x62 && ~x2 && ~x19 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y23 = 1'b1;	
							nx_state = s411;
						end
					else if( ~x61 && ~x62 )
						nx_state = s1;
					else nx_state = s321;
				s322 : if( 1'b1 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s262;
						end
					else nx_state = s322;
				s323 : if( x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x3 )
						nx_state = s1;
					else nx_state = s323;
				s324 : if( 1'b1 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s414;
						end
					else nx_state = s324;
				s325 : if( 1'b1 )
						nx_state = s40;
					else nx_state = s325;
				s326 : if( 1'b1 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else nx_state = s326;
				s327 : if( 1'b1 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else nx_state = s327;
				s328 : if( x65 && x60 && x61 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s38;
						end
					else if( x65 && x60 && ~x61 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s68;
						end
					else if( x65 && ~x60 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s68;
						end
					else if( ~x65 && x68 && x19 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s375;
						end
					else if( ~x65 && x68 && ~x19 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x68 && x21 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x65 && ~x68 && ~x21 )
						begin
							y8 = 1'b1;	y14 = 1'b1;	
							nx_state = s378;
						end
					else nx_state = s328;
				s329 : if( x65 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s66;
						end
					else if( ~x65 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else nx_state = s329;
				s330 : if( x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x18 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x21 && x22 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x21 && x22 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x17 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && x18 && x14 )
						nx_state = s40;
					else if( ~x21 && x22 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s40;
					else if( ~x21 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && x7 && x9 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x21 && ~x22 && x23 && x7 && x9 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x21 && ~x22 && x23 && x7 && x9 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && x7 && x9 && ~x19 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && x7 && ~x9 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s333;
						end
					else if( ~x21 && ~x22 && x23 && ~x7 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x21 && ~x22 && x23 && ~x7 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x21 && ~x22 && x23 && ~x7 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x7 && ~x19 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else nx_state = s330;
				s331 : if( x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x18 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && x18 && x14 )
						nx_state = s40;
					else if( ~x21 && x22 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s40;
					else if( ~x21 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x19 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else nx_state = s331;
				s332 : if( x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x18 )
						nx_state = s1;
					else if( ~x21 && x23 && x22 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x21 && x23 && ~x22 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s180;
						end
					else if( ~x21 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else nx_state = s332;
				s333 : if( x21 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s143;
						end
					else if( ~x21 && x22 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x21 && x22 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x21 && x22 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x17 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x19 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 )
						begin
							y3 = 1'b1;	
							nx_state = s320;
						end
					else nx_state = s333;
				s334 : if( 1'b1 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else nx_state = s334;
				s335 : if( 1'b1 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s341;
						end
					else nx_state = s335;
				s336 : if( x68 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( x68 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( x68 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( x68 && ~x7 )
						nx_state = s1;
					else if( ~x68 && x21 )
						begin
							y5 = 1'b1;	
							nx_state = s343;
						end
					else if( ~x68 && ~x21 && x22 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x68 && ~x21 && x22 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x68 && ~x21 && x22 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x68 && ~x21 && x22 && x23 && ~x17 )
						nx_state = s1;
					else if( ~x68 && ~x21 && x22 && ~x23 && x18 && x14 )
						nx_state = s40;
					else if( ~x68 && ~x21 && x22 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s40;
					else if( ~x68 && ~x21 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x68 && ~x21 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x68 && ~x21 && ~x22 && x23 )
						nx_state = s1;
					else if( ~x68 && ~x21 && ~x22 && ~x23 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s180;
						end
					else nx_state = s336;
				s337 : if( x23 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s333;
						end
					else if( ~x23 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else nx_state = s337;
				s338 : if( x65 && x66 )
						nx_state = s316;
					else if( x65 && ~x66 && x67 && x8 && x9 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x65 && ~x66 && x67 && x8 && ~x9 && x10 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	y19 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s136;
						end
					else if( x65 && ~x66 && x67 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( x65 && ~x66 && x67 && ~x8 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x19 && x18 && x14 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	y25 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && ~x66 && ~x67 && x19 && x18 && ~x14 && x17 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	y25 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && ~x66 && ~x67 && x19 && x18 && ~x14 && ~x17 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x19 && x18 && ~x14 && ~x17 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && x19 && x18 && ~x14 && ~x17 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x19 && x18 && ~x14 && ~x17 && ~x5 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && x19 && ~x18 )
						begin
							y6 = 1'b1;	y8 = 1'b1;	y25 = 1'b1;	
							nx_state = s1;
						end
					else if( x65 && ~x66 && ~x67 && ~x19 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && ~x19 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && ~x66 && ~x67 && ~x19 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x66 && ~x67 && ~x19 && ~x5 )
						nx_state = s1;
					else if( ~x65 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else nx_state = s338;
				s339 : if( x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x21 && ~x18 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && x4 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else if( ~x21 && x22 && x23 && ~x4 && x18 && x15 && x10 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x21 && x22 && x23 && ~x4 && x18 && x15 && ~x10 && x12 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && x22 && x23 && ~x4 && x18 && x15 && ~x10 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s285;
						end
					else if( ~x21 && x22 && x23 && ~x4 && x18 && ~x15 && x16 && x10 && x12 )
						begin
							y14 = 1'b1;	
							nx_state = s286;
						end
					else if( ~x21 && x22 && x23 && ~x4 && x18 && ~x15 && x16 && x10 && ~x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x21 && x22 && x23 && ~x4 && x18 && ~x15 && x16 && ~x10 )
						begin
							y14 = 1'b1;	
							nx_state = s286;
						end
					else if( ~x21 && x22 && x23 && ~x4 && x18 && ~x15 && ~x16 )
						nx_state = s40;
					else if( ~x21 && x22 && x23 && ~x4 && ~x18 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x21 && x22 && ~x23 && x18 && x14 )
						nx_state = s40;
					else if( ~x21 && x22 && ~x23 && x18 && ~x14 && x13 )
						nx_state = s40;
					else if( ~x21 && x22 && ~x23 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 && ~x18 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x19 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else nx_state = s339;
				s340 : if( x21 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x21 && x22 && x15 && x10 && x16 && x12 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x21 && x22 && x15 && x10 && x16 && ~x12 )
						begin
							y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s339;
						end
					else if( ~x21 && x22 && x15 && x10 && ~x16 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x21 && x22 && x15 && x10 && ~x16 && ~x3 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x21 && x22 && x15 && x10 && ~x16 && ~x3 && ~x2 && x11 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s126;
						end
					else if( ~x21 && x22 && x15 && x10 && ~x16 && ~x3 && ~x2 && ~x11 && x12 )
						begin
							y3 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							y20 = 1'b1;	
							nx_state = s332;
						end
					else if( ~x21 && x22 && x15 && x10 && ~x16 && ~x3 && ~x2 && ~x11 && ~x12 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	
							nx_state = s330;
						end
					else if( ~x21 && x22 && x15 && ~x10 && x11 && x12 && x16 )
						begin
							y14 = 1'b1;	
							nx_state = s331;
						end
					else if( ~x21 && x22 && x15 && ~x10 && x11 && x12 && ~x16 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x21 && x22 && x15 && ~x10 && x11 && x12 && ~x16 && ~x3 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x21 && x22 && x15 && ~x10 && x11 && x12 && ~x16 && ~x3 && ~x2 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s336;
						end
					else if( ~x21 && x22 && x15 && ~x10 && x11 && ~x12 && x16 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && x15 && ~x10 && x11 && ~x12 && ~x16 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y13 = 1'b1;	
							nx_state = s333;
						end
					else if( ~x21 && x22 && x15 && ~x10 && ~x11 && x16 && x12 && x13 )
						begin
							y11 = 1'b1;	
							nx_state = s122;
						end
					else if( ~x21 && x22 && x15 && ~x10 && ~x11 && x16 && x12 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x22 && x15 && ~x10 && ~x11 && x16 && ~x12 && x14 )
						begin
							y11 = 1'b1;	
							nx_state = s122;
						end
					else if( ~x21 && x22 && x15 && ~x10 && ~x11 && x16 && ~x12 && ~x14 )
						nx_state = s1;
					else if( ~x21 && x22 && x15 && ~x10 && ~x11 && ~x16 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x21 && x22 && x15 && ~x10 && ~x11 && ~x16 && ~x3 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x21 && x22 && x15 && ~x10 && ~x11 && ~x16 && ~x3 && ~x2 && x12 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x21 && x22 && x15 && ~x10 && ~x11 && ~x16 && ~x3 && ~x2 && ~x12 )
						begin
							y14 = 1'b1;	
							nx_state = s48;
						end
					else if( ~x21 && x22 && ~x15 && x16 && x12 && x10 && x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x15 && x16 && x12 && x10 && ~x8 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x21 && x22 && ~x15 && x16 && x12 && x10 && ~x8 && ~x3 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x21 && x22 && ~x15 && x16 && x12 && x10 && ~x8 && ~x3 && ~x2 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x21 && x22 && ~x15 && x16 && x12 && ~x10 && x11 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x21 && x22 && ~x15 && x16 && x12 && ~x10 && x11 && ~x3 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x21 && x22 && ~x15 && x16 && x12 && ~x10 && x11 && ~x3 && ~x2 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x21 && x22 && ~x15 && x16 && x12 && ~x10 && ~x11 && x7 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x21 && x22 && ~x15 && x16 && x12 && ~x10 && ~x11 && x7 && ~x3 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s69;
						end
					else if( ~x21 && x22 && ~x15 && x16 && x12 && ~x10 && ~x11 && x7 && ~x3 && ~x2 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x21 && x22 && ~x15 && x16 && x12 && ~x10 && ~x11 && ~x7 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && x10 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && x10 && ~x3 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s264;
						end
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && x10 && ~x3 && ~x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && ~x10 && x11 && x9 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && ~x10 && x11 && x9 && ~x3 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && ~x10 && x11 && x9 && ~x3 && ~x2 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && ~x10 && x11 && ~x9 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && ~x10 && ~x11 && x8 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && ~x10 && ~x11 && x8 && ~x3 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && ~x10 && ~x11 && x8 && ~x3 && ~x2 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x21 && x22 && ~x15 && x16 && ~x12 && ~x10 && ~x11 && ~x8 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x15 && ~x16 && x3 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x21 && x22 && ~x15 && ~x16 && ~x3 && x2 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x21 && x22 && ~x15 && ~x16 && ~x3 && ~x2 )
						begin
							y7 = 1'b1;	y8 = 1'b1;	
							nx_state = s110;
						end
					else if( ~x21 && ~x22 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x21 && ~x22 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x23 && ~x19 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x23 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else nx_state = s340;
				s341 : if( x68 && x7 && x8 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( x68 && x7 && ~x8 && x9 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( x68 && x7 && ~x8 && ~x9 )
						nx_state = s1;
					else if( x68 && ~x7 )
						nx_state = s1;
					else if( ~x68 && x21 && x18 && x14 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x68 && x21 && x18 && ~x14 && x13 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s144;
						end
					else if( ~x68 && x21 && x18 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x68 && x21 && ~x18 )
						nx_state = s1;
					else if( ~x68 && ~x21 && x22 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x68 && ~x21 && x22 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x68 && ~x21 && x22 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x68 && ~x21 && x22 && x23 && ~x17 )
						nx_state = s1;
					else if( ~x68 && ~x21 && x22 && ~x23 )
						begin
							y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s301;
						end
					else if( ~x68 && ~x21 && ~x22 && x23 && x19 && x14 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x68 && ~x21 && ~x22 && x23 && x19 && ~x14 && x13 )
						begin
							y7 = 1'b1;	y10 = 1'b1;	y21 = 1'b1;	
							y22 = 1'b1;	
							nx_state = s145;
						end
					else if( ~x68 && ~x21 && ~x22 && x23 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x68 && ~x21 && ~x22 && x23 && ~x19 )
						nx_state = s1;
					else if( ~x68 && ~x21 && ~x22 && ~x23 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s180;
						end
					else nx_state = s341;
				s342 : if( x66 && x22 )
						begin
							y11 = 1'b1;	
							nx_state = s122;
						end
					else if( x66 && ~x22 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x66 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	
							nx_state = s142;
						end
					else nx_state = s342;
				s343 : if( x66 && x21 )
						begin
							y1 = 1'b1;	
							nx_state = s22;
						end
					else if( x66 && ~x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s86;
						end
					else if( ~x66 )
						begin
							y10 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else nx_state = s343;
				s344 : if( x21 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x21 && ~x20 )
						nx_state = s1;
					else nx_state = s344;
				s345 : if( x68 && x15 && x10 && x11 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s192;
						end
					else if( x68 && x15 && x10 && ~x11 && x12 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s193;
						end
					else if( x68 && x15 && x10 && ~x11 && ~x12 )
						begin
							y1 = 1'b1;	y8 = 1'b1;	y13 = 1'b1;	
							nx_state = s192;
						end
					else if( x68 && x15 && ~x10 && x12 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s300;
						end
					else if( x68 && x15 && ~x10 && ~x12 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y10 = 1'b1;	
							nx_state = s192;
						end
					else if( x68 && ~x15 && x16 && x10 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x68 && ~x15 && x16 && x10 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x68 && ~x15 && x16 && x10 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x68 && ~x15 && x16 && x10 && ~x19 )
						nx_state = s1;
					else if( x68 && ~x15 && x16 && ~x10 && x12 && x11 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	y7 = 1'b1;	
							y11 = 1'b1;	
							nx_state = s199;
						end
					else if( x68 && ~x15 && x16 && ~x10 && x12 && ~x11 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x68 && ~x15 && x16 && ~x10 && x12 && ~x11 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x68 && ~x15 && x16 && ~x10 && x12 && ~x11 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x68 && ~x15 && x16 && ~x10 && x12 && ~x11 && ~x19 )
						nx_state = s1;
					else if( x68 && ~x15 && x16 && ~x10 && ~x12 && x19 && x14 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x68 && ~x15 && x16 && ~x10 && ~x12 && x19 && ~x14 && x13 )
						begin
							y22 = 1'b1;	
							nx_state = s4;
						end
					else if( x68 && ~x15 && x16 && ~x10 && ~x12 && x19 && ~x14 && ~x13 )
						nx_state = s1;
					else if( x68 && ~x15 && x16 && ~x10 && ~x12 && ~x19 )
						nx_state = s1;
					else if( x68 && ~x15 && ~x16 )
						begin
							y5 = 1'b1;	y7 = 1'b1;	y8 = 1'b1;	
							y9 = 1'b1;	
							nx_state = s201;
						end
					else if( ~x68 )
						begin
							y1 = 1'b1;	y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s72;
						end
					else nx_state = s345;
				s346 : if( x67 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x67 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x67 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x67 && ~x4 )
						nx_state = s1;
					else if( ~x67 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x67 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x67 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x67 && ~x5 )
						nx_state = s1;
					else nx_state = s346;
				s347 : if( x19 && x20 && x11 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x19 && x20 && ~x11 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x19 && x20 && ~x11 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x19 && x20 && ~x11 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x19 && x20 && ~x11 && ~x5 )
						nx_state = s1;
					else if( x19 && ~x20 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x19 && ~x20 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x19 && ~x20 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x19 && ~x20 && ~x5 )
						nx_state = s1;
					else if( ~x19 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x19 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x19 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x19 && ~x5 )
						nx_state = s1;
					else nx_state = s347;
				s348 : if( x19 && x17 && x20 && x14 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( x19 && x17 && x20 && ~x14 )
						begin
							y4 = 1'b1;	y29 = 1'b1;	y32 = 1'b1;	
							nx_state = s351;
						end
					else if( x19 && x17 && ~x20 && x14 )
						begin
							y4 = 1'b1;	y18 = 1'b1;	y29 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s351;
						end
					else if( x19 && x17 && ~x20 && ~x14 && x15 )
						begin
							y16 = 1'b1;	y28 = 1'b1;	
							nx_state = s352;
						end
					else if( x19 && x17 && ~x20 && ~x14 && ~x15 && x16 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	y32 = 1'b1;	
							nx_state = s351;
						end
					else if( x19 && x17 && ~x20 && ~x14 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s351;
						end
					else if( x19 && ~x17 && x18 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	y19 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s349;
						end
					else if( x19 && ~x17 && ~x18 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x19 && x20 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x19 && ~x20 && x17 && x16 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s351;
						end
					else if( ~x19 && ~x20 && x17 && ~x16 && x15 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x19 && ~x20 && x17 && ~x16 && ~x15 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x19 && ~x20 && ~x17 && x18 && x4 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s415;
						end
					else if( ~x19 && ~x20 && ~x17 && x18 && ~x4 )
						begin
							y7 = 1'b1;	
							nx_state = s338;
						end
					else if( ~x19 && ~x20 && ~x17 && ~x18 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else nx_state = s348;
				s349 : if( x19 && x11 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x19 && ~x11 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x19 && ~x11 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x19 && ~x11 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x19 && ~x11 && ~x5 )
						nx_state = s1;
					else if( ~x19 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x19 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x19 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x19 && ~x5 )
						nx_state = s1;
					else nx_state = s349;
				s350 : if( x19 && x14 && x20 )
						begin
							y7 = 1'b1;	
							nx_state = s338;
						end
					else if( x19 && x14 && ~x20 )
						begin
							y2 = 1'b1;	y21 = 1'b1;	
							nx_state = s416;
						end
					else if( x19 && ~x14 )
						begin
							y7 = 1'b1;	
							nx_state = s338;
						end
					else if( ~x19 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x19 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x19 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x19 && ~x5 )
						nx_state = s1;
					else nx_state = s350;
				s351 : if( x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x5 )
						nx_state = s1;
					else nx_state = s351;
				s352 : if( x19 && x20 && x9 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s415;
						end
					else if( x19 && x20 && ~x9 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( x19 && ~x20 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x19 && ~x20 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x19 && ~x20 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x19 && ~x20 && ~x5 )
						nx_state = s1;
					else if( ~x19 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x19 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x19 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( ~x19 && ~x5 )
						nx_state = s1;
					else nx_state = s352;
				s353 : if( x65 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x5 )
						nx_state = s1;
					else if( ~x65 && x21 )
						begin
							y17 = 1'b1;	
							nx_state = s77;
						end
					else if( ~x65 && ~x21 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s344;
						end
					else nx_state = s353;
				s354 : if( 1'b1 )
						begin
							y14 = 1'b1;	
							nx_state = s417;
						end
					else nx_state = s354;
				s355 : if( x65 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x65 )
						begin
							y15 = 1'b1;	y112 = 1'b1;	
							nx_state = s46;
						end
					else nx_state = s355;
				s356 : if( x65 && x60 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s63;
						end
					else if( x65 && ~x60 && x61 && x62 )
						begin
							y1 = 1'b1;	y4 = 1'b1;	y23 = 1'b1;	
							nx_state = s411;
						end
					else if( x65 && ~x60 && x61 && ~x62 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s63;
						end
					else if( x65 && ~x60 && ~x61 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x65 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else nx_state = s356;
				s357 : if( x65 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x65 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else nx_state = s357;
				s358 : if( x21 && x18 && x10 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x21 && x18 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x21 && x18 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x21 && x18 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x21 && x18 && ~x10 && ~x4 )
						nx_state = s1;
					else if( x21 && ~x18 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x21 && ~x18 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x21 && ~x18 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x21 && ~x18 && ~x4 )
						nx_state = s1;
					else if( ~x21 && x22 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && x22 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x4 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x20 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x22 && x20 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x22 && x20 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x20 && ~x4 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x20 && x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x22 && ~x20 && x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x22 && ~x20 && x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x20 && x19 && ~x4 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x20 && ~x19 && x10 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && ~x22 && ~x20 && ~x19 && ~x10 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x22 && ~x20 && ~x19 && ~x10 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x22 && ~x20 && ~x19 && ~x10 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x20 && ~x19 && ~x10 && ~x4 )
						nx_state = s1;
					else nx_state = s358;
				s359 : if( x21 && x16 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x21 && x16 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s360;
						end
					else if( x21 && ~x16 && x17 && x18 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s418;
						end
					else if( x21 && ~x16 && x17 && x18 && ~x3 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s249;
						end
					else if( x21 && ~x16 && x17 && x18 && ~x3 && ~x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( x21 && ~x16 && x17 && ~x18 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( x21 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && x22 && x16 && x19 && x18 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x21 && x22 && x16 && x19 && x18 && ~x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s362;
						end
					else if( ~x21 && x22 && x16 && x19 && ~x18 && x13 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && x16 && x19 && ~x18 && ~x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x21 && x22 && x16 && ~x19 && x13 )
						begin
							y3 = 1'b1;	y16 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && x22 && x16 && ~x19 && ~x13 && x18 && x15 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && x16 && ~x19 && ~x13 && x18 && ~x15 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && x22 && x16 && ~x19 && ~x13 && ~x18 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x21 && x22 && ~x16 && x17 && x18 && x19 && x10 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s418;
						end
					else if( ~x21 && x22 && ~x16 && x17 && x18 && x19 && x10 && ~x3 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else if( ~x21 && x22 && ~x16 && x17 && x18 && x19 && ~x10 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && x22 && ~x16 && x17 && x18 && ~x19 && x13 && x3 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s419;
						end
					else if( ~x21 && x22 && ~x16 && x17 && x18 && ~x19 && x13 && ~x3 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else if( ~x21 && x22 && ~x16 && x17 && x18 && ~x19 && ~x13 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && x22 && ~x16 && x17 && ~x18 && x13 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s418;
						end
					else if( ~x21 && x22 && ~x16 && x17 && ~x18 && x13 && ~x3 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else if( ~x21 && x22 && ~x16 && x17 && ~x18 && ~x13 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && x22 && ~x16 && x17 && ~x18 && ~x13 && ~x19 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( ~x21 && x22 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && ~x22 && x19 && x17 && x13 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && ~x22 && x19 && x17 && ~x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x21 && ~x22 && x19 && ~x17 && x18 && x13 && x3 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else if( ~x21 && ~x22 && x19 && ~x17 && x18 && x13 && ~x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s418;
						end
					else if( ~x21 && ~x22 && x19 && ~x17 && x18 && ~x13 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( ~x21 && ~x22 && x19 && ~x17 && ~x18 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && ~x22 && ~x19 && x16 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x21 && ~x22 && ~x19 && x16 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s360;
						end
					else if( ~x21 && ~x22 && ~x19 && ~x16 && x17 && x20 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( ~x21 && ~x22 && ~x19 && ~x16 && x17 && ~x20 && x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s418;
						end
					else if( ~x21 && ~x22 && ~x19 && ~x16 && x17 && ~x20 && ~x3 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x21 && ~x22 && ~x19 && ~x16 && x17 && ~x20 && ~x3 && ~x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( ~x21 && ~x22 && ~x19 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s146;
						end
					else nx_state = s359;
				s360 : if( x21 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x21 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x21 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x21 && ~x4 )
						nx_state = s1;
					else if( ~x21 && x22 && x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && x22 && x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && x22 && x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && x19 && ~x4 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x18 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && x22 && ~x19 && x18 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && x22 && ~x19 && x18 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && x18 && ~x4 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x19 && ~x18 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	
							nx_state = s300;
						end
					else if( ~x21 && ~x22 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x22 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s360;
				s361 : if( x22 && x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x22 && x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x22 && x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x22 && x19 && ~x4 )
						nx_state = s1;
					else if( x22 && ~x19 && x18 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x22 && ~x19 && x18 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x22 && ~x19 && x18 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x22 && ~x19 && x18 && ~x4 )
						nx_state = s1;
					else if( x22 && ~x19 && ~x18 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x22 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x22 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s361;
				s362 : if( x22 && x19 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x22 && x19 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x22 && x19 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x22 && x19 && ~x4 )
						nx_state = s1;
					else if( x22 && ~x19 && x18 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( x22 && ~x19 && ~x18 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x22 && ~x19 && ~x18 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x22 && ~x19 && ~x18 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x22 && ~x19 && ~x18 && ~x4 )
						nx_state = s1;
					else if( ~x22 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x22 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x22 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s362;
				s363 : if( x65 && x67 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x67 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x65 && x67 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x65 && x67 && ~x4 )
						nx_state = s1;
					else if( x65 && ~x67 && x21 )
						begin
							y4 = 1'b1;	y22 = 1'b1;	y38 = 1'b1;	
							nx_state = s95;
						end
					else if( x65 && ~x67 && ~x21 )
						begin
							y35 = 1'b1;	
							nx_state = s26;
						end
					else if( ~x65 )
						begin
							y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s288;
						end
					else nx_state = s363;
				s364 : if( x19 && x18 && x14 )
						begin
							y7 = 1'b1;	
							nx_state = s338;
						end
					else if( x19 && x18 && ~x14 && x17 )
						begin
							y7 = 1'b1;	
							nx_state = s338;
						end
					else if( x19 && x18 && ~x14 && ~x17 && x20 )
						begin
							y7 = 1'b1;	
							nx_state = s30;
						end
					else if( x19 && x18 && ~x14 && ~x17 && ~x20 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( x19 && ~x18 )
						begin
							y7 = 1'b1;	
							nx_state = s338;
						end
					else if( ~x19 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else nx_state = s364;
				s365 : if( 1'b1 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else nx_state = s365;
				s366 : if( x20 && x15 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s198;
						end
					else if( x20 && ~x15 && x16 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s59;
						end
					else if( x20 && ~x15 && ~x16 )
						begin
							y7 = 1'b1;	y12 = 1'b1;	
							nx_state = s211;
						end
					else if( ~x20 && x21 && x17 && x15 && x8 )
						begin
							y8 = 1'b1;	y10 = 1'b1;	
							nx_state = s254;
						end
					else if( ~x20 && x21 && x17 && x15 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x20 && x21 && x17 && ~x15 && x16 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x20 && x21 && x17 && ~x15 && ~x16 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s209;
						end
					else if( ~x20 && x21 && ~x17 )
						nx_state = s40;
					else if( ~x20 && ~x21 && x3 )
						nx_state = s40;
					else if( ~x20 && ~x21 && ~x3 && x18 && x15 && x8 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( ~x20 && ~x21 && ~x3 && x18 && x15 && ~x8 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	y10 = 1'b1;	
							nx_state = s198;
						end
					else if( ~x20 && ~x21 && ~x3 && x18 && ~x15 && x16 )
						begin
							y10 = 1'b1;	y14 = 1'b1;	
							nx_state = s47;
						end
					else if( ~x20 && ~x21 && ~x3 && x18 && ~x15 && ~x16 )
						begin
							y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s209;
						end
					else if( ~x20 && ~x21 && ~x3 && ~x18 )
						nx_state = s39;
					else nx_state = s366;
				s367 : if( x61 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( ~x61 && x15 && x12 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s292;
						end
					else if( ~x61 && x15 && x12 && ~x7 )
						begin
							y12 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x61 && x15 && ~x12 && x7 )
						begin
							y7 = 1'b1;	y14 = 1'b1;	y23 = 1'b1;	
							nx_state = s63;
						end
					else if( ~x61 && x15 && ~x12 && ~x7 )
						begin
							y2 = 1'b1;	y10 = 1'b1;	y20 = 1'b1;	
							nx_state = s263;
						end
					else if( ~x61 && ~x15 && x16 && x7 && x12 )
						begin
							y12 = 1'b1;	
							nx_state = s290;
						end
					else if( ~x61 && ~x15 && x16 && x7 && ~x12 )
						begin
							y5 = 1'b1;	y10 = 1'b1;	
							nx_state = s262;
						end
					else if( ~x61 && ~x15 && x16 && ~x7 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s258;
						end
					else if( ~x61 && ~x15 && ~x16 && x7 )
						begin
							y12 = 1'b1;	
							nx_state = s100;
						end
					else if( ~x61 && ~x15 && ~x16 && ~x7 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else nx_state = s367;
				s368 : if( x22 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s314;
						end
					else if( ~x22 && x19 && x15 && x8 )
						begin
							y11 = 1'b1;	
							nx_state = s8;
						end
					else if( ~x22 && x19 && x15 && ~x8 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	
							nx_state = s111;
						end
					else if( ~x22 && x19 && ~x15 && x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	
							nx_state = s50;
						end
					else if( ~x22 && x19 && ~x15 && ~x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x22 && ~x19 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	
							nx_state = s314;
						end
					else nx_state = s368;
				s369 : if( x4 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	
							nx_state = s168;
						end
					else if( ~x4 && x42 && x15 && x8 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else if( ~x4 && x42 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x4 && x42 && ~x15 && x16 )
						begin
							y21 = 1'b1;	
							nx_state = s151;
						end
					else if( ~x4 && x42 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y28 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x4 && ~x42 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y14 = 1'b1;	
							y16 = 1'b1;	
							nx_state = s400;
						end
					else nx_state = s369;
				s370 : if( x21 )
						begin
							y14 = 1'b1;	
							nx_state = s155;
						end
					else if( ~x21 && x22 && x23 && x17 && x14 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x21 && x22 && x23 && x17 && ~x14 && x13 )
						begin
							y1 = 1'b1;	y7 = 1'b1;	y16 = 1'b1;	
							nx_state = s87;
						end
					else if( ~x21 && x22 && x23 && x17 && ~x14 && ~x13 )
						nx_state = s1;
					else if( ~x21 && x22 && x23 && ~x17 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x23 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s341;
						end
					else if( ~x21 && ~x22 )
						begin
							y4 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s180;
						end
					else nx_state = s370;
				s371 : if( x22 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x22 && x21 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x22 && ~x21 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x22 && ~x21 && x4 && ~x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x22 && ~x21 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x22 && ~x21 && ~x4 )
						nx_state = s1;
					else nx_state = s371;
				s372 : if( 1'b1 )
						begin
							y2 = 1'b1;	y11 = 1'b1;	y17 = 1'b1;	
							nx_state = s123;
						end
					else nx_state = s372;
				s373 : if( x21 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x21 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x5 && ~x4 && x22 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x5 && ~x4 && x22 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x5 && ~x4 && ~x22 )
						nx_state = s1;
					else if( ~x21 && ~x5 && x22 )
						nx_state = s1;
					else if( ~x21 && ~x5 && ~x22 && x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && ~x5 && ~x22 && x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x5 && ~x22 && ~x4 )
						nx_state = s1;
					else nx_state = s373;
				s374 : if( x66 && x16 && x21 && x7 && x10 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s67;
						end
					else if( x66 && x16 && x21 && x7 && ~x10 )
						begin
							y5 = 1'b1;	y18 = 1'b1;	
							nx_state = s113;
						end
					else if( x66 && x16 && x21 && ~x7 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s67;
						end
					else if( x66 && x16 && ~x21 && x7 && x10 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s75;
						end
					else if( x66 && x16 && ~x21 && x7 && ~x10 )
						begin
							y4 = 1'b1;	y18 = 1'b1;	
							nx_state = s395;
						end
					else if( x66 && x16 && ~x21 && ~x7 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s75;
						end
					else if( x66 && ~x16 && x17 && x9 && x21 && x10 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s67;
						end
					else if( x66 && ~x16 && x17 && x9 && x21 && ~x10 && x13 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s67;
						end
					else if( x66 && ~x16 && x17 && x9 && x21 && ~x10 && ~x13 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && ~x16 && x17 && x9 && x21 && ~x10 && ~x13 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && ~x16 && x17 && x9 && x21 && ~x10 && ~x13 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x66 && ~x16 && x17 && x9 && x21 && ~x10 && ~x13 && ~x19 )
						nx_state = s1;
					else if( x66 && ~x16 && x17 && x9 && ~x21 && x10 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s75;
						end
					else if( x66 && ~x16 && x17 && x9 && ~x21 && ~x10 && x13 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s75;
						end
					else if( x66 && ~x16 && x17 && x9 && ~x21 && ~x10 && ~x13 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x66 && ~x16 && x17 && x9 && ~x21 && ~x10 && ~x13 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x66 && ~x16 && x17 && x9 && ~x21 && ~x10 && ~x13 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x66 && ~x16 && x17 && x9 && ~x21 && ~x10 && ~x13 && ~x20 )
						nx_state = s1;
					else if( x66 && ~x16 && x17 && ~x9 && x21 && x10 && x11 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s67;
						end
					else if( x66 && ~x16 && x17 && ~x9 && x21 && x10 && ~x11 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && ~x16 && x17 && ~x9 && x21 && x10 && ~x11 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && ~x16 && x17 && ~x9 && x21 && x10 && ~x11 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x66 && ~x16 && x17 && ~x9 && x21 && x10 && ~x11 && ~x19 )
						nx_state = s1;
					else if( x66 && ~x16 && x17 && ~x9 && x21 && ~x10 && x12 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s67;
						end
					else if( x66 && ~x16 && x17 && ~x9 && x21 && ~x10 && ~x12 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && ~x16 && x17 && ~x9 && x21 && ~x10 && ~x12 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( x66 && ~x16 && x17 && ~x9 && x21 && ~x10 && ~x12 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x66 && ~x16 && x17 && ~x9 && x21 && ~x10 && ~x12 && ~x19 )
						nx_state = s1;
					else if( x66 && ~x16 && x17 && ~x9 && ~x21 && x10 && x11 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s75;
						end
					else if( x66 && ~x16 && x17 && ~x9 && ~x21 && x10 && ~x11 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x66 && ~x16 && x17 && ~x9 && ~x21 && x10 && ~x11 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x66 && ~x16 && x17 && ~x9 && ~x21 && x10 && ~x11 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x66 && ~x16 && x17 && ~x9 && ~x21 && x10 && ~x11 && ~x20 )
						nx_state = s1;
					else if( x66 && ~x16 && x17 && ~x9 && ~x21 && ~x10 && x12 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s75;
						end
					else if( x66 && ~x16 && x17 && ~x9 && ~x21 && ~x10 && ~x12 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x66 && ~x16 && x17 && ~x9 && ~x21 && ~x10 && ~x12 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( x66 && ~x16 && x17 && ~x9 && ~x21 && ~x10 && ~x12 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( x66 && ~x16 && x17 && ~x9 && ~x21 && ~x10 && ~x12 && ~x20 )
						nx_state = s1;
					else if( x66 && ~x16 && ~x17 && x7 )
						begin
							y4 = 1'b1;	y17 = 1'b1;	
							nx_state = s353;
						end
					else if( x66 && ~x16 && ~x17 && ~x7 && x21 )
						begin
							y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s67;
						end
					else if( x66 && ~x16 && ~x17 && ~x7 && ~x21 )
						begin
							y4 = 1'b1;	y8 = 1'b1;	
							nx_state = s75;
						end
					else if( ~x66 && x21 && x3 && x4 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x66 && x21 && x3 && ~x4 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x66 && x21 && x3 && ~x4 && ~x5 )
						nx_state = s1;
					else if( ~x66 && x21 && ~x3 )
						nx_state = s1;
					else if( ~x66 && ~x21 && x22 && x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x66 && ~x21 && x22 && x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x66 && ~x21 && x22 && x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x66 && ~x21 && x22 && ~x6 )
						nx_state = s1;
					else if( ~x66 && ~x21 && ~x22 && x8 && x9 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x66 && ~x21 && ~x22 && x8 && ~x9 && x10 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	
							nx_state = s88;
						end
					else if( ~x66 && ~x21 && ~x22 && x8 && ~x9 && ~x10 )
						nx_state = s1;
					else if( ~x66 && ~x21 && ~x22 && ~x8 )
						nx_state = s1;
					else nx_state = s374;
				s375 : if( x21 )
						nx_state = s1;
					else if( ~x21 && x22 )
						begin
							y13 = 1'b1;	
							nx_state = s413;
						end
					else if( ~x21 && ~x22 && x5 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else if( ~x21 && ~x22 && ~x5 && x7 && x18 && x15 )
						begin
							y8 = 1'b1;	y18 = 1'b1;	
							nx_state = s82;
						end
					else if( ~x21 && ~x22 && ~x5 && x7 && x18 && ~x15 )
						begin
							y2 = 1'b1;	y4 = 1'b1;	
							nx_state = s374;
						end
					else if( ~x21 && ~x22 && ~x5 && x7 && ~x18 && x19 && x15 )
						begin
							y3 = 1'b1;	
							nx_state = s320;
						end
					else if( ~x21 && ~x22 && ~x5 && x7 && ~x18 && x19 && ~x15 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( ~x21 && ~x22 && ~x5 && x7 && ~x18 && ~x19 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( ~x21 && ~x22 && ~x5 && ~x7 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s385;
						end
					else nx_state = s375;
				s376 : if( x21 )
						begin
							y18 = 1'b1;	
							nx_state = s203;
						end
					else if( ~x21 && x22 )
						begin
							y1 = 1'b1;	y6 = 1'b1;	
							nx_state = s142;
						end
					else if( ~x21 && ~x22 )
						begin
							y18 = 1'b1;	
							nx_state = s114;
						end
					else nx_state = s376;
				s377 : if( x22 && x21 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s123;
						end
					else if( x22 && ~x21 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( x22 && ~x21 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( x22 && ~x21 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( x22 && ~x21 && ~x5 )
						nx_state = s1;
					else if( ~x22 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y17 = 1'b1;	
							y18 = 1'b1;	
							nx_state = s123;
						end
					else nx_state = s377;
				s378 : if( x21 )
						begin
							y18 = 1'b1;	y19 = 1'b1;	
							nx_state = s126;
						end
					else if( ~x21 && x22 && x5 && x4 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && x5 && ~x4 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && x5 && ~x4 && ~x6 )
						nx_state = s1;
					else if( ~x21 && x22 && ~x5 )
						nx_state = s1;
					else if( ~x21 && ~x22 && x19 && x15 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x21 && ~x22 && x19 && ~x15 && x12 )
						begin
							y2 = 1'b1;	y6 = 1'b1;	y18 = 1'b1;	
							nx_state = s123;
						end
					else if( ~x21 && ~x22 && x19 && ~x15 && ~x12 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x21 && ~x22 && ~x19 && x20 && x14 && x15 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x21 && ~x22 && ~x19 && x20 && x14 && ~x15 && x18 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x21 && ~x22 && ~x19 && x20 && x14 && ~x15 && ~x18 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && ~x22 && ~x19 && x20 && x14 && ~x15 && ~x18 && x4 && ~x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && ~x22 && ~x19 && x20 && x14 && ~x15 && ~x18 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x19 && x20 && x14 && ~x15 && ~x18 && ~x4 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x19 && x20 && ~x14 && x15 && x16 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x21 && ~x22 && ~x19 && x20 && ~x14 && x15 && ~x16 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && ~x22 && ~x19 && x20 && ~x14 && x15 && ~x16 && x4 && ~x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && ~x22 && ~x19 && x20 && ~x14 && x15 && ~x16 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x19 && x20 && ~x14 && x15 && ~x16 && ~x4 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x19 && x20 && ~x14 && ~x15 && x17 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s103;
						end
					else if( ~x21 && ~x22 && ~x19 && x20 && ~x14 && ~x15 && ~x17 && x4 && x5 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && ~x22 && ~x19 && x20 && ~x14 && ~x15 && ~x17 && x4 && ~x5 && x6 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && ~x22 && ~x19 && x20 && ~x14 && ~x15 && ~x17 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x19 && x20 && ~x14 && ~x15 && ~x17 && ~x4 )
						nx_state = s1;
					else if( ~x21 && ~x22 && ~x19 && ~x20 && x12 )
						begin
							y6 = 1'b1;	y21 = 1'b1;	
							nx_state = s225;
						end
					else if( ~x21 && ~x22 && ~x19 && ~x20 && ~x12 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	y6 = 1'b1;	
							nx_state = s103;
						end
					else nx_state = s378;
				s379 : if( 1'b1 )
						begin
							y8 = 1'b1;	y12 = 1'b1;	y13 = 1'b1;	
							nx_state = s106;
						end
					else nx_state = s379;
				s380 : if( 1'b1 )
						begin
							y21 = 1'b1;	
							nx_state = s7;
						end
					else nx_state = s380;
				s381 : if( 1'b1 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else nx_state = s381;
				s382 : if( 1'b1 )
						begin
							y11 = 1'b1;	y13 = 1'b1;	
							nx_state = s52;
						end
					else nx_state = s382;
				s383 : if( 1'b1 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else nx_state = s383;
				s384 : if( 1'b1 )
						begin
							y18 = 1'b1;	
							nx_state = s394;
						end
					else nx_state = s384;
				s385 : if( x21 && x8 )
						begin
							y3 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s275;
						end
					else if( x21 && ~x8 && x19 && x18 && x17 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s272;
						end
					else if( x21 && ~x8 && x19 && x18 && x17 && ~x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s272;
						end
					else if( x21 && ~x8 && x19 && x18 && ~x17 && x12 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x21 && ~x8 && x19 && x18 && ~x17 && ~x12 )
						begin
							y4 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s273;
						end
					else if( x21 && ~x8 && x19 && ~x18 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s274;
						end
					else if( x21 && ~x8 && ~x19 && x9 && x20 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s272;
						end
					else if( x21 && ~x8 && ~x19 && x9 && x20 && ~x12 )
						begin
							y2 = 1'b1;	y9 = 1'b1;	y10 = 1'b1;	
							nx_state = s105;
						end
					else if( x21 && ~x8 && ~x19 && x9 && ~x20 && x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s270;
						end
					else if( x21 && ~x8 && ~x19 && x9 && ~x20 && ~x12 )
						begin
							y16 = 1'b1;	y18 = 1'b1;	
							nx_state = s109;
						end
					else if( x21 && ~x8 && ~x19 && ~x9 )
						begin
							y9 = 1'b1;	y17 = 1'b1;	y18 = 1'b1;	
							nx_state = s274;
						end
					else if( ~x21 && x22 )
						nx_state = s1;
					else if( ~x21 && ~x22 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s102;
						end
					else nx_state = s385;
				s386 : if( x6 && x7 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( x6 && ~x7 && x8 )
						begin
							y8 = 1'b1;	y19 = 1'b1;	
							nx_state = s138;
						end
					else if( x6 && ~x7 && ~x8 )
						nx_state = s1;
					else if( ~x6 )
						nx_state = s1;
					else nx_state = s386;
				s387 : if( 1'b1 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s388;
						end
					else nx_state = s387;
				s388 : if( 1'b1 )
						begin
							y13 = 1'b1;	
							nx_state = s265;
						end
					else nx_state = s388;
				s389 : if( 1'b1 )
						begin
							y3 = 1'b1;	y5 = 1'b1;	
							nx_state = s255;
						end
					else nx_state = s389;
				s390 : if( x21 && x20 )
						begin
							y5 = 1'b1;	y6 = 1'b1;	
							nx_state = s133;
						end
					else if( x21 && ~x20 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else nx_state = s390;
				s391 : if( x3 )
						begin
							y3 = 1'b1;	y7 = 1'b1;	y11 = 1'b1;	
							nx_state = s420;
						end
					else if( ~x3 && x8 && x21 && x16 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x3 && x8 && x21 && x16 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s360;
						end
					else if( ~x3 && x8 && x21 && ~x16 && x17 && x18 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x3 && x8 && x21 && ~x16 && x17 && x18 && ~x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( ~x3 && x8 && x21 && ~x16 && x17 && ~x18 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( ~x3 && x8 && x21 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x3 && x8 && ~x21 && x22 && x16 && x19 && x18 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x3 && x8 && ~x21 && x22 && x16 && x19 && x18 && ~x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s362;
						end
					else if( ~x3 && x8 && ~x21 && x22 && x16 && x19 && ~x18 && x13 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x3 && x8 && ~x21 && x22 && x16 && x19 && ~x18 && ~x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x3 && x8 && ~x21 && x22 && x16 && ~x19 && x13 )
						begin
							y3 = 1'b1;	y16 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x3 && x8 && ~x21 && x22 && x16 && ~x19 && ~x13 && x18 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x3 && x8 && ~x21 && x22 && x16 && ~x19 && ~x13 && ~x18 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x3 && x8 && ~x21 && x22 && ~x16 && x17 && x19 && x18 && x10 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else if( ~x3 && x8 && ~x21 && x22 && ~x16 && x17 && x19 && x18 && ~x10 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x3 && x8 && ~x21 && x22 && ~x16 && x17 && x19 && ~x18 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else if( ~x3 && x8 && ~x21 && x22 && ~x16 && x17 && x19 && ~x18 && ~x13 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x3 && x8 && ~x21 && x22 && ~x16 && x17 && ~x19 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else if( ~x3 && x8 && ~x21 && x22 && ~x16 && x17 && ~x19 && ~x13 && x18 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x3 && x8 && ~x21 && x22 && ~x16 && x17 && ~x19 && ~x13 && ~x18 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( ~x3 && x8 && ~x21 && x22 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && x19 && x17 && x13 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && x19 && x17 && ~x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && x19 && ~x17 && x18 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && x19 && ~x17 && x18 && ~x13 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && x19 && ~x17 && ~x18 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && ~x19 && x16 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && ~x19 && x16 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s360;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && ~x19 && ~x16 && x17 && x20 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && ~x19 && ~x16 && x17 && ~x20 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && ~x19 && ~x16 && x17 && ~x20 && ~x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( ~x3 && x8 && ~x21 && ~x22 && ~x19 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x3 && ~x8 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s421;
						end
					else nx_state = s391;
				s392 : if( x68 )
						begin
							y6 = 1'b1;	y7 = 1'b1;	
							nx_state = s76;
						end
					else if( ~x68 )
						begin
							y5 = 1'b1;	y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s282;
						end
					else nx_state = s392;
				s393 : if( x20 && x18 && x13 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x20 && x18 && ~x13 && x12 )
						begin
							y9 = 1'b1;	
							nx_state = s27;
						end
					else if( x20 && x18 && ~x13 && ~x12 )
						nx_state = s1;
					else if( x20 && ~x18 )
						nx_state = s1;
					else if( ~x20 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else nx_state = s393;
				s394 : if( 1'b1 )
						begin
							y4 = 1'b1;	y21 = 1'b1;	
							nx_state = s273;
						end
					else nx_state = s394;
				s395 : if( x65 && x5 && x6 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x5 && ~x6 && x7 )
						begin
							y5 = 1'b1;	
							nx_state = s101;
						end
					else if( x65 && x5 && ~x6 && ~x7 )
						nx_state = s1;
					else if( x65 && ~x5 )
						nx_state = s1;
					else if( ~x65 && x21 && x19 && x15 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && x21 && x19 && ~x15 && x14 )
						begin
							y8 = 1'b1;	
							nx_state = s92;
						end
					else if( ~x65 && x21 && x19 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && x21 && ~x19 )
						nx_state = s1;
					else if( ~x65 && ~x21 && x20 && x15 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x65 && ~x21 && x20 && ~x15 && x14 )
						begin
							y27 = 1'b1;	
							nx_state = s3;
						end
					else if( ~x65 && ~x21 && x20 && ~x15 && ~x14 )
						nx_state = s1;
					else if( ~x65 && ~x21 && ~x20 )
						nx_state = s1;
					else nx_state = s395;
				s396 : if( 1'b1 )
						begin
							y8 = 1'b1;	y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s375;
						end
					else nx_state = s396;
				s397 : if( x63 && x15 && x8 )
						begin
							y2 = 1'b1;	y3 = 1'b1;	
							nx_state = s23;
						end
					else if( x63 && x15 && ~x8 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x63 && ~x15 && x16 )
						begin
							y19 = 1'b1;	
							nx_state = s11;
						end
					else if( x63 && ~x15 && ~x16 )
						begin
							y13 = 1'b1;	y14 = 1'b1;	y29 = 1'b1;	
							nx_state = s135;
						end
					else if( ~x63 )
						nx_state = s1;
					else nx_state = s397;
				s398 : if( x19 && x14 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( x19 && ~x14 && x13 )
						begin
							y11 = 1'b1;	y12 = 1'b1;	
							nx_state = s175;
						end
					else if( x19 && ~x14 && ~x13 )
						nx_state = s398;
					else if( ~x19 )
						nx_state = s1;
					else nx_state = s398;
				s399 : if( x66 )
						begin
							y15 = 1'b1;	y16 = 1'b1;	
							nx_state = s137;
						end
					else if( ~x66 )
						begin
							y11 = 1'b1;	
							nx_state = s53;
						end
					else nx_state = s399;
				s400 : if( 1'b1 )
						begin
							y3 = 1'b1;	y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s130;
						end
					else nx_state = s400;
				s401 : if( x20 )
						begin
							y2 = 1'b1;	y7 = 1'b1;	y13 = 1'b1;	
							nx_state = s366;
						end
					else if( ~x20 )
						nx_state = s1;
					else nx_state = s401;
				s402 : if( x25 && x24 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( x25 && ~x24 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x25 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else nx_state = s402;
				s403 : if( 1'b1 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s59;
						end
					else nx_state = s403;
				s404 : if( x3 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	
							nx_state = s250;
						end
					else if( ~x3 && x19 )
						begin
							y14 = 1'b1;	
							nx_state = s285;
						end
					else if( ~x3 && ~x19 )
						begin
							y14 = 1'b1;	y21 = 1'b1;	y22 = 1'b1;	
							nx_state = s84;
						end
					else nx_state = s404;
				s405 : if( x21 && x20 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( x21 && ~x20 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s302;
						end
					else if( ~x21 )
						begin
							y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s302;
						end
					else nx_state = s405;
				s406 : if( 1'b1 )
						begin
							y8 = 1'b1;	
							nx_state = s246;
						end
					else nx_state = s406;
				s407 : if( 1'b1 )
						begin
							y20 = 1'b1;	
							nx_state = s13;
						end
					else nx_state = s407;
				s408 : if( x21 && x18 && x16 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else if( x21 && x18 && ~x16 && x17 && x13 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else if( x21 && x18 && ~x16 && x17 && ~x13 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x21 && x18 && ~x16 && x17 && ~x13 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x21 && x18 && ~x16 && x17 && ~x13 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x21 && x18 && ~x16 && x17 && ~x13 && ~x4 )
						nx_state = s1;
					else if( x21 && x18 && ~x16 && ~x17 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else if( x21 && ~x18 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x21 && ~x18 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( x21 && ~x18 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( x21 && ~x18 && ~x4 )
						nx_state = s1;
					else if( ~x21 && x19 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x21 && ~x19 && x22 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x21 && ~x19 && ~x22 && x20 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x19 && ~x22 && x20 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x19 && ~x22 && x20 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x19 && ~x22 && x20 && ~x4 )
						nx_state = s1;
					else if( ~x21 && ~x19 && ~x22 && ~x20 && x16 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && x13 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && ~x13 && x17 && x4 && x5 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && ~x13 && x17 && x4 && ~x5 && x6 )
						begin
							y10 = 1'b1;	
							nx_state = s12;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && ~x13 && x17 && x4 && ~x5 && ~x6 )
						nx_state = s1;
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && ~x13 && x17 && ~x4 )
						nx_state = s1;
					else if( ~x21 && ~x19 && ~x22 && ~x20 && ~x16 && ~x13 && ~x17 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s408;
				s409 : if( x21 && x18 && x13 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x21 && x18 && ~x13 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else if( x21 && ~x18 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x21 && x22 && x18 && x19 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && x22 && x18 && ~x19 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( ~x21 && x22 && ~x18 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && ~x22 && x19 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && ~x22 && ~x19 && x13 && x20 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else if( ~x21 && ~x22 && ~x19 && x13 && ~x20 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && ~x22 && ~x19 && ~x13 )
						begin
							y5 = 1'b1;	y16 = 1'b1;	y17 = 1'b1;	
							nx_state = s1;
						end
					else nx_state = s409;
				s410 : if( 1'b1 )
						begin
							y9 = 1'b1;	y14 = 1'b1;	
							nx_state = s336;
						end
					else nx_state = s410;
				s411 : if( x61 )
						nx_state = s1;
					else if( ~x61 )
						begin
							y2 = 1'b1;	y8 = 1'b1;	
							nx_state = s367;
						end
					else nx_state = s411;
				s412 : if( x4 && x19 && x20 && x14 )
						begin
							y16 = 1'b1;	y28 = 1'b1;	
							nx_state = s422;
						end
					else if( x4 && x19 && x20 && ~x14 && x16 )
						begin
							y16 = 1'b1;	y28 = 1'b1;	
							nx_state = s422;
						end
					else if( x4 && x19 && x20 && ~x14 && ~x16 && x17 )
						begin
							y16 = 1'b1;	y28 = 1'b1;	
							nx_state = s352;
						end
					else if( x4 && x19 && x20 && ~x14 && ~x16 && ~x17 )
						begin
							y16 = 1'b1;	y28 = 1'b1;	
							nx_state = s422;
						end
					else if( x4 && x19 && ~x20 )
						begin
							y16 = 1'b1;	y28 = 1'b1;	
							nx_state = s422;
						end
					else if( x4 && ~x19 )
						begin
							y16 = 1'b1;	y28 = 1'b1;	
							nx_state = s422;
						end
					else if( ~x4 && x9 && x17 && x19 && x20 && x14 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( ~x4 && x9 && x17 && x19 && x20 && ~x14 && x16 )
						begin
							y4 = 1'b1;	y29 = 1'b1;	y32 = 1'b1;	
							nx_state = s351;
						end
					else if( ~x4 && x9 && x17 && x19 && x20 && ~x14 && ~x16 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s415;
						end
					else if( ~x4 && x9 && x17 && x19 && ~x20 && x14 )
						begin
							y4 = 1'b1;	y18 = 1'b1;	y29 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s351;
						end
					else if( ~x4 && x9 && x17 && x19 && ~x20 && ~x14 && x16 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	y32 = 1'b1;	
							nx_state = s351;
						end
					else if( ~x4 && x9 && x17 && x19 && ~x20 && ~x14 && ~x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s351;
						end
					else if( ~x4 && x9 && x17 && ~x19 && x16 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s351;
						end
					else if( ~x4 && x9 && x17 && ~x19 && ~x16 && x20 )
						begin
							y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s351;
						end
					else if( ~x4 && x9 && x17 && ~x19 && ~x16 && ~x20 && x15 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x4 && x9 && x17 && ~x19 && ~x16 && ~x20 && ~x15 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x4 && x9 && ~x17 && x18 && x19 && x14 && x16 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	y19 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s349;
						end
					else if( ~x4 && x9 && ~x17 && x18 && x19 && x14 && ~x16 )
						begin
							y2 = 1'b1;	y21 = 1'b1;	
							nx_state = s416;
						end
					else if( ~x4 && x9 && ~x17 && x18 && x19 && ~x14 )
						begin
							y7 = 1'b1;	
							nx_state = s338;
						end
					else if( ~x4 && x9 && ~x17 && x18 && ~x19 )
						begin
							y7 = 1'b1;	
							nx_state = s338;
						end
					else if( ~x4 && x9 && ~x17 && ~x18 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x4 && ~x9 && x19 && x20 && x17 && x16 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s415;
						end
					else if( ~x4 && ~x9 && x19 && x20 && x17 && ~x16 && x14 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s415;
						end
					else if( ~x4 && ~x9 && x19 && x20 && x17 && ~x16 && ~x14 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( ~x4 && ~x9 && x19 && x20 && ~x17 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s415;
						end
					else if( ~x4 && ~x9 && x19 && ~x20 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s415;
						end
					else if( ~x4 && ~x9 && ~x19 && x20 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s415;
						end
					else if( ~x4 && ~x9 && ~x19 && ~x20 && x17 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s415;
						end
					else if( ~x4 && ~x9 && ~x19 && ~x20 && ~x17 && x18 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s241;
						end
					else if( ~x4 && ~x9 && ~x19 && ~x20 && ~x17 && ~x18 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s415;
						end
					else nx_state = s412;
				s413 : if( x22 )
						begin
							y3 = 1'b1;	y14 = 1'b1;	y15 = 1'b1;	
							nx_state = s385;
						end
					else if( ~x22 )
						begin
							y3 = 1'b1;	
							nx_state = s320;
						end
					else nx_state = s413;
				s414 : if( 1'b1 )
						begin
							y7 = 1'b1;	
							nx_state = s140;
						end
					else nx_state = s414;
				s415 : if( x17 && x19 && x20 && x14 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( x17 && x19 && x20 && ~x14 && x16 )
						begin
							y4 = 1'b1;	y29 = 1'b1;	y32 = 1'b1;	
							nx_state = s351;
						end
					else if( x17 && x19 && x20 && ~x14 && ~x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( x17 && x19 && ~x20 && x14 )
						begin
							y4 = 1'b1;	y18 = 1'b1;	y29 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s351;
						end
					else if( x17 && x19 && ~x20 && ~x14 && x16 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	y32 = 1'b1;	
							nx_state = s351;
						end
					else if( x17 && x19 && ~x20 && ~x14 && ~x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s351;
						end
					else if( x17 && ~x19 && x16 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s351;
						end
					else if( x17 && ~x19 && ~x16 && x20 )
						begin
							y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s351;
						end
					else if( x17 && ~x19 && ~x16 && ~x20 && x15 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( x17 && ~x19 && ~x16 && ~x20 && ~x15 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x17 && x18 && x19 && x14 && x16 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	y19 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s349;
						end
					else if( ~x17 && x18 && x19 && x14 && ~x16 )
						begin
							y2 = 1'b1;	y21 = 1'b1;	
							nx_state = s416;
						end
					else if( ~x17 && x18 && x19 && ~x14 )
						begin
							y7 = 1'b1;	
							nx_state = s338;
						end
					else if( ~x17 && x18 && ~x19 )
						begin
							y7 = 1'b1;	
							nx_state = s338;
						end
					else if( ~x17 && ~x18 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else nx_state = s415;
				s416 : if( x20 )
						begin
							y8 = 1'b1;	
							nx_state = s246;
						end
					else if( ~x20 )
						begin
							y6 = 1'b1;	y20 = 1'b1;	
							nx_state = s102;
						end
					else nx_state = s416;
				s417 : if( 1'b1 )
						begin
							y4 = 1'b1;	y5 = 1'b1;	y9 = 1'b1;	
							nx_state = s80;
						end
					else nx_state = s417;
				s418 : if( x21 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s249;
						end
					else if( x21 && ~x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( ~x21 && x19 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else if( ~x21 && ~x19 && x22 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else if( ~x21 && ~x19 && ~x22 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x21 && ~x19 && ~x22 && ~x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else nx_state = s418;
				s419 : if( 1'b1 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else nx_state = s419;
				s420 : if( x8 && x21 && x16 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x8 && x21 && x16 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s360;
						end
					else if( x8 && x21 && ~x16 && x17 && x18 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s249;
						end
					else if( x8 && x21 && ~x16 && x17 && x18 && ~x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( x8 && x21 && ~x16 && x17 && ~x18 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( x8 && x21 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s146;
						end
					else if( x8 && ~x21 && x22 && x16 && x19 && x18 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( x8 && ~x21 && x22 && x16 && x19 && x18 && ~x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s362;
						end
					else if( x8 && ~x21 && x22 && x16 && x19 && ~x18 && x13 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( x8 && ~x21 && x22 && x16 && x19 && ~x18 && ~x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x8 && ~x21 && x22 && x16 && ~x19 && x13 )
						begin
							y3 = 1'b1;	y16 = 1'b1;	
							nx_state = s146;
						end
					else if( x8 && ~x21 && x22 && x16 && ~x19 && ~x13 && x18 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s146;
						end
					else if( x8 && ~x21 && x22 && x16 && ~x19 && ~x13 && ~x18 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( x8 && ~x21 && x22 && ~x16 && x17 && x19 && x18 && x10 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else if( x8 && ~x21 && x22 && ~x16 && x17 && x19 && x18 && ~x10 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s146;
						end
					else if( x8 && ~x21 && x22 && ~x16 && x17 && x19 && ~x18 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else if( x8 && ~x21 && x22 && ~x16 && x17 && x19 && ~x18 && ~x13 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( x8 && ~x21 && x22 && ~x16 && x17 && ~x19 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else if( x8 && ~x21 && x22 && ~x16 && x17 && ~x19 && ~x13 && x18 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( x8 && ~x21 && x22 && ~x16 && x17 && ~x19 && ~x13 && ~x18 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( x8 && ~x21 && x22 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s146;
						end
					else if( x8 && ~x21 && ~x22 && x19 && x17 && x13 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( x8 && ~x21 && ~x22 && x19 && x17 && ~x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( x8 && ~x21 && ~x22 && x19 && ~x17 && x18 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else if( x8 && ~x21 && ~x22 && x19 && ~x17 && x18 && ~x13 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( x8 && ~x21 && ~x22 && x19 && ~x17 && ~x18 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s146;
						end
					else if( x8 && ~x21 && ~x22 && ~x19 && x16 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x8 && ~x21 && ~x22 && ~x19 && x16 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s360;
						end
					else if( x8 && ~x21 && ~x22 && ~x19 && ~x16 && x17 && x20 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( x8 && ~x21 && ~x22 && ~x19 && ~x16 && x17 && ~x20 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s249;
						end
					else if( x8 && ~x21 && ~x22 && ~x19 && ~x16 && x17 && ~x20 && ~x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( x8 && ~x21 && ~x22 && ~x19 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x8 )
						begin
							y3 = 1'b1;	y8 = 1'b1;	y12 = 1'b1;	
							y13 = 1'b1;	
							nx_state = s421;
						end
					else nx_state = s420;
				s421 : if( x21 && x16 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x21 && x16 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s360;
						end
					else if( x21 && ~x16 && x17 && x18 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s249;
						end
					else if( x21 && ~x16 && x17 && x18 && ~x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( x21 && ~x16 && x17 && ~x18 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( x21 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && x22 && x16 && x19 && x18 && x10 )
						begin
							y3 = 1'b1;	
							nx_state = s89;
						end
					else if( ~x21 && x22 && x16 && x19 && x18 && ~x10 )
						begin
							y5 = 1'b1;	y8 = 1'b1;	y11 = 1'b1;	
							y12 = 1'b1;	
							nx_state = s362;
						end
					else if( ~x21 && x22 && x16 && x19 && ~x18 && x13 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && x22 && x16 && x19 && ~x18 && ~x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x21 && x22 && x16 && ~x19 && x13 )
						begin
							y3 = 1'b1;	y16 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && x22 && x16 && ~x19 && ~x13 && x18 )
						begin
							y5 = 1'b1;	y12 = 1'b1;	y26 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && x22 && x16 && ~x19 && ~x13 && ~x18 )
						begin
							y24 = 1'b1;	
							nx_state = s278;
						end
					else if( ~x21 && x22 && ~x16 && x17 && x18 && x19 && x10 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else if( ~x21 && x22 && ~x16 && x17 && x18 && x19 && ~x10 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y18 = 1'b1;	
							y19 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && x22 && ~x16 && x17 && x18 && ~x19 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else if( ~x21 && x22 && ~x16 && x17 && x18 && ~x19 && ~x13 )
						begin
							y16 = 1'b1;	
							nx_state = s16;
						end
					else if( ~x21 && x22 && ~x16 && x17 && ~x18 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else if( ~x21 && x22 && ~x16 && x17 && ~x18 && ~x13 && x19 )
						begin
							y7 = 1'b1;	y15 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && x22 && ~x16 && x17 && ~x18 && ~x13 && ~x19 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( ~x21 && x22 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && ~x22 && x19 && x17 && x13 )
						begin
							y15 = 1'b1;	
							nx_state = s149;
						end
					else if( ~x21 && ~x22 && x19 && x17 && ~x13 )
						begin
							y23 = 1'b1;	
							nx_state = s83;
						end
					else if( ~x21 && ~x22 && x19 && ~x17 && x18 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s248;
						end
					else if( ~x21 && ~x22 && x19 && ~x17 && x18 && ~x13 )
						begin
							y7 = 1'b1;	y11 = 1'b1;	y15 = 1'b1;	
							nx_state = s358;
						end
					else if( ~x21 && ~x22 && x19 && ~x17 && ~x18 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s146;
						end
					else if( ~x21 && ~x22 && ~x19 && x16 && x13 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( ~x21 && ~x22 && ~x19 && x16 && ~x13 )
						begin
							y7 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s360;
						end
					else if( ~x21 && ~x22 && ~x19 && ~x16 && x17 && x20 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( ~x21 && ~x22 && ~x19 && ~x16 && x17 && ~x20 && x13 )
						begin
							y1 = 1'b1;	y25 = 1'b1;	
							nx_state = s249;
						end
					else if( ~x21 && ~x22 && ~x19 && ~x16 && x17 && ~x20 && ~x13 )
						begin
							y2 = 1'b1;	y12 = 1'b1;	y15 = 1'b1;	
							nx_state = s408;
						end
					else if( ~x21 && ~x22 && ~x19 && ~x16 && ~x17 )
						begin
							y8 = 1'b1;	y9 = 1'b1;	y11 = 1'b1;	
							nx_state = s146;
						end
					else nx_state = s421;
				s422 : if( x9 && x17 && x19 && x20 && x14 )
						begin
							y2 = 1'b1;	
							nx_state = s56;
						end
					else if( x9 && x17 && x19 && x20 && ~x14 )
						begin
							y4 = 1'b1;	y29 = 1'b1;	y32 = 1'b1;	
							nx_state = s351;
						end
					else if( x9 && x17 && x19 && ~x20 && x14 )
						begin
							y4 = 1'b1;	y18 = 1'b1;	y29 = 1'b1;	
							y32 = 1'b1;	
							nx_state = s351;
						end
					else if( x9 && x17 && x19 && ~x20 && ~x14 && x16 )
						begin
							y29 = 1'b1;	y31 = 1'b1;	y32 = 1'b1;	
							nx_state = s351;
						end
					else if( x9 && x17 && x19 && ~x20 && ~x14 && ~x16 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	y18 = 1'b1;	
							nx_state = s351;
						end
					else if( x9 && x17 && ~x19 && x16 )
						begin
							y29 = 1'b1;	y30 = 1'b1;	
							nx_state = s351;
						end
					else if( x9 && x17 && ~x19 && ~x16 && x20 )
						begin
							y9 = 1'b1;	y26 = 1'b1;	
							nx_state = s351;
						end
					else if( x9 && x17 && ~x19 && ~x16 && ~x20 && x15 )
						begin
							y4 = 1'b1;	y11 = 1'b1;	
							nx_state = s112;
						end
					else if( x9 && x17 && ~x19 && ~x16 && ~x20 && ~x15 )
						begin
							y25 = 1'b1;	
							nx_state = s78;
						end
					else if( x9 && ~x17 && x18 && x19 && x14 && x16 )
						begin
							y2 = 1'b1;	y14 = 1'b1;	y19 = 1'b1;	
							y29 = 1'b1;	y30 = 1'b1;	y32 = 1'b1;	
							nx_state = s349;
						end
					else if( x9 && ~x17 && x18 && x19 && x14 && ~x16 )
						begin
							y2 = 1'b1;	y21 = 1'b1;	
							nx_state = s416;
						end
					else if( x9 && ~x17 && x18 && x19 && ~x14 )
						begin
							y7 = 1'b1;	
							nx_state = s338;
						end
					else if( x9 && ~x17 && x18 && ~x19 )
						begin
							y7 = 1'b1;	
							nx_state = s338;
						end
					else if( x9 && ~x17 && ~x18 )
						begin
							y4 = 1'b1;	
							nx_state = s43;
						end
					else if( ~x9 && x19 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s415;
						end
					else if( ~x9 && ~x19 && x20 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s415;
						end
					else if( ~x9 && ~x19 && ~x20 && x17 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s415;
						end
					else if( ~x9 && ~x19 && ~x20 && ~x17 && x18 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s241;
						end
					else if( ~x9 && ~x19 && ~x20 && ~x17 && ~x18 )
						begin
							y17 = 1'b1;	y20 = 1'b1;	y28 = 1'b1;	
							nx_state = s415;
						end
					else nx_state = s422;

			default : nx_state = 0;
		endcase
	end
endmodule
